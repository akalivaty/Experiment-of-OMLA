//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n800, new_n802, new_n803, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G141gat), .B(G148gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n204), .B1(KEYINPUT2), .B2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G155gat), .B(G162gat), .Z(new_n207));
  AOI21_X1  g006(.A(KEYINPUT72), .B1(G155gat), .B2(G162gat), .ZN(new_n208));
  OR3_X1    g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n207), .B1(new_n206), .B2(new_n208), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT73), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n213));
  XNOR2_X1  g012(.A(G197gat), .B(G204gat), .ZN(new_n214));
  XOR2_X1   g013(.A(KEYINPUT68), .B(G218gat), .Z(new_n215));
  INV_X1    g014(.A(G211gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n214), .B1(new_n217), .B2(KEYINPUT22), .ZN(new_n218));
  XNOR2_X1  g017(.A(G211gat), .B(G218gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n213), .B1(new_n220), .B2(KEYINPUT29), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n212), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n211), .A2(new_n213), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT29), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n220), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n203), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n211), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n221), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n230), .A2(G228gat), .A3(G233gat), .A4(new_n226), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(new_n232), .B(G22gat), .Z(new_n233));
  XOR2_X1   g032(.A(KEYINPUT31), .B(G50gat), .Z(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n232), .B(G22gat), .ZN(new_n236));
  INV_X1    g035(.A(new_n234), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(G78gat), .B(G106gat), .Z(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(KEYINPUT76), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT77), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n235), .A2(new_n238), .A3(new_n242), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(G15gat), .B(G43gat), .Z(new_n247));
  XNOR2_X1  g046(.A(G71gat), .B(G99gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(G169gat), .A2(G176gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT23), .ZN(new_n251));
  AND2_X1   g050(.A1(G183gat), .A2(G190gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n251), .B1(new_n253), .B2(KEYINPUT24), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(new_n252), .ZN(new_n256));
  NAND2_X1  g055(.A1(G169gat), .A2(G176gat), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n257), .B1(new_n250), .B2(KEYINPUT23), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n254), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT25), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT65), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n261), .B1(KEYINPUT25), .B2(new_n259), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT27), .B(G183gat), .ZN(new_n263));
  INV_X1    g062(.A(G190gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n265), .B(KEYINPUT28), .Z(new_n266));
  INV_X1    g065(.A(KEYINPUT26), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n250), .B1(new_n267), .B2(new_n257), .ZN(new_n268));
  NOR3_X1   g067(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n253), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT66), .ZN(new_n271));
  OR2_X1    g070(.A1(new_n270), .A2(KEYINPUT66), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n266), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n262), .A2(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(G127gat), .B(G134gat), .Z(new_n275));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n276));
  XOR2_X1   g075(.A(G113gat), .B(G120gat), .Z(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n278), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n274), .B(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G227gat), .ZN(new_n284));
  INV_X1    g083(.A(G233gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT64), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n249), .B1(new_n288), .B2(KEYINPUT33), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT32), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OR2_X1    g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT34), .B1(new_n283), .B2(new_n286), .ZN(new_n293));
  OR3_X1    g092(.A1(new_n283), .A2(KEYINPUT34), .A3(new_n287), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(new_n291), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n292), .A2(new_n293), .A3(new_n294), .A4(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n293), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n289), .A2(new_n291), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n289), .A2(new_n291), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n246), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT81), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT81), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(new_n246), .B2(new_n301), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n262), .A2(new_n273), .ZN(new_n307));
  INV_X1    g106(.A(G226gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n308), .A2(new_n285), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n307), .B(KEYINPUT69), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n224), .B1(new_n308), .B2(new_n285), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n220), .B(new_n310), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(G8gat), .B(G36gat), .Z(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(KEYINPUT70), .ZN(new_n315));
  XNOR2_X1  g114(.A(G64gat), .B(G92gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n307), .A2(new_n312), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n319), .B1(new_n311), .B2(new_n309), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n313), .B(new_n318), .C1(new_n320), .C2(new_n220), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT30), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(KEYINPUT71), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n313), .B1(new_n320), .B2(new_n220), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n317), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n322), .B1(new_n321), .B2(KEYINPUT71), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n211), .A2(new_n281), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT4), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT74), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n212), .A2(new_n282), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n331), .B1(new_n332), .B2(KEYINPUT4), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT5), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n229), .A2(KEYINPUT3), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(new_n282), .A3(new_n223), .ZN(new_n336));
  NAND2_X1  g135(.A1(G225gat), .A2(G233gat), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n333), .A2(new_n334), .A3(new_n336), .A4(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G1gat), .B(G29gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT0), .ZN(new_n340));
  XNOR2_X1  g139(.A(G57gat), .B(G85gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  INV_X1    g141(.A(new_n337), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT4), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n343), .B1(new_n329), .B2(new_n344), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n336), .B(new_n345), .C1(new_n332), .C2(new_n344), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n211), .B(new_n281), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n334), .B1(new_n347), .B2(new_n343), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n338), .A2(new_n342), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT6), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(KEYINPUT75), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n342), .B1(new_n338), .B2(new_n349), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n353), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n328), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n202), .B1(new_n306), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n353), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(new_n351), .A3(new_n350), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n353), .A2(KEYINPUT6), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n362), .A2(KEYINPUT80), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(KEYINPUT80), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n361), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AND4_X1   g164(.A1(new_n202), .A2(new_n302), .A3(new_n328), .A4(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n246), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n357), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n324), .A2(KEYINPUT37), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n369), .A2(new_n318), .ZN(new_n370));
  INV_X1    g169(.A(new_n220), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n371), .B(new_n310), .C1(new_n311), .C2(new_n312), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n372), .B(KEYINPUT37), .C1(new_n320), .C2(new_n371), .ZN(new_n373));
  OR2_X1    g172(.A1(new_n373), .A2(KEYINPUT79), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(KEYINPUT79), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT38), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n377), .B1(new_n324), .B2(KEYINPUT37), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n376), .A2(new_n377), .B1(new_n370), .B2(new_n378), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n321), .B(new_n361), .C1(new_n363), .C2(new_n364), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n333), .A2(new_n336), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n343), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n347), .A2(new_n343), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OR2_X1    g183(.A1(new_n384), .A2(KEYINPUT78), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(KEYINPUT78), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n382), .A2(KEYINPUT39), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n387), .B(new_n342), .C1(KEYINPUT39), .C2(new_n382), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT40), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n389), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n360), .A3(new_n391), .ZN(new_n392));
  OAI22_X1  g191(.A1(new_n379), .A2(new_n380), .B1(new_n328), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n368), .B1(new_n393), .B2(new_n367), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n301), .A2(KEYINPUT36), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT36), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n396), .B1(new_n296), .B2(new_n300), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  OAI22_X1  g198(.A1(new_n359), .A2(new_n366), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(G8gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(G15gat), .B(G22gat), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT16), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n402), .B1(new_n403), .B2(G1gat), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n401), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n404), .B1(G1gat), .B2(new_n402), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI221_X1 g207(.A(new_n404), .B1(new_n405), .B2(new_n401), .C1(G1gat), .C2(new_n402), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT88), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT84), .B(KEYINPUT15), .ZN(new_n413));
  INV_X1    g212(.A(G50gat), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT85), .B1(new_n414), .B2(G43gat), .ZN(new_n415));
  INV_X1    g214(.A(G43gat), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n415), .B1(new_n416), .B2(G50gat), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n414), .A2(KEYINPUT85), .A3(G43gat), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n413), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n416), .A2(G50gat), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n414), .A2(G43gat), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT15), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G29gat), .A2(G36gat), .ZN(new_n425));
  OR3_X1    g224(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n419), .A2(new_n424), .A3(new_n425), .A4(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n426), .B1(new_n430), .B2(new_n427), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n427), .A2(new_n430), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n425), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n423), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n412), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n429), .A2(new_n434), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT17), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n435), .A2(KEYINPUT17), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n409), .B(new_n408), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G229gat), .A2(G233gat), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n442), .B(KEYINPUT87), .Z(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n436), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(KEYINPUT89), .A2(KEYINPUT18), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n446), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n436), .A2(new_n441), .A3(new_n444), .A4(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n410), .B(KEYINPUT88), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n437), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n443), .B(KEYINPUT13), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n447), .A2(new_n449), .A3(new_n454), .ZN(new_n455));
  XOR2_X1   g254(.A(G113gat), .B(G141gat), .Z(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(KEYINPUT11), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n457), .B(G169gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(G197gat), .ZN(new_n459));
  INV_X1    g258(.A(G169gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n457), .B(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(G197gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT12), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n464), .A2(KEYINPUT12), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n455), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT82), .B1(new_n466), .B2(new_n467), .ZN(new_n471));
  OR2_X1    g270(.A1(new_n464), .A2(KEYINPUT12), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT82), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n473), .A3(new_n465), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(new_n455), .A3(KEYINPUT90), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT90), .B1(new_n475), .B2(new_n455), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n470), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n400), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT91), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT91), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n400), .A2(new_n482), .A3(new_n479), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G71gat), .B(G78gat), .ZN(new_n485));
  AND2_X1   g284(.A1(G57gat), .A2(G64gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(G57gat), .A2(G64gat), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G71gat), .A2(G78gat), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT92), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT9), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n490), .B1(new_n489), .B2(new_n491), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n485), .B(new_n488), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  OR2_X1    g293(.A1(G57gat), .A2(G64gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(G57gat), .A2(G64gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(KEYINPUT9), .A3(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(G71gat), .A2(G78gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(G71gat), .A2(G78gat), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT21), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(G231gat), .A2(G233gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(KEYINPUT93), .B(KEYINPUT19), .Z(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(G127gat), .B(G155gat), .Z(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT20), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n508), .B(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n450), .B1(new_n503), .B2(new_n502), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT94), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n511), .B(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(G183gat), .B(G211gat), .Z(new_n515));
  AND2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n435), .B(new_n438), .ZN(new_n520));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT8), .ZN(new_n522));
  NAND2_X1  g321(.A1(G85gat), .A2(G92gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G85gat), .ZN(new_n526));
  INV_X1    g325(.A(G92gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n522), .A2(new_n525), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G99gat), .B(G106gat), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(KEYINPUT95), .A3(new_n532), .ZN(new_n533));
  AOI22_X1  g332(.A1(KEYINPUT8), .A2(new_n521), .B1(new_n526), .B2(new_n527), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n534), .A2(new_n531), .A3(new_n525), .A4(new_n529), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT95), .B1(new_n530), .B2(new_n532), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n520), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g338(.A1(G232gat), .A2(G233gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT41), .ZN(new_n541));
  INV_X1    g340(.A(new_n538), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n541), .B1(new_n437), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G190gat), .B(G218gat), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n539), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n539), .B2(new_n543), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n546), .B(new_n547), .C1(KEYINPUT41), .C2(new_n540), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n540), .A2(KEYINPUT41), .ZN(new_n549));
  INV_X1    g348(.A(new_n547), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n549), .B1(new_n550), .B2(new_n545), .ZN(new_n551));
  XOR2_X1   g350(.A(G134gat), .B(G162gat), .Z(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n548), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(new_n548), .B2(new_n551), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G120gat), .B(G148gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(G176gat), .B(G204gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT10), .ZN(new_n561));
  NOR3_X1   g360(.A1(new_n542), .A2(new_n561), .A3(new_n502), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n502), .B1(new_n536), .B2(new_n537), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n495), .A2(new_n496), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(new_n500), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT92), .B1(new_n498), .B2(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n566), .A2(new_n569), .B1(new_n500), .B2(new_n497), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT96), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n530), .A2(new_n532), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .A4(new_n535), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n572), .A2(new_n494), .A3(new_n501), .A4(new_n535), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT96), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n564), .A2(new_n573), .A3(new_n575), .A4(new_n561), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n576), .A2(KEYINPUT97), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(KEYINPUT97), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n563), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT99), .ZN(new_n580));
  NAND2_X1  g379(.A1(G230gat), .A2(G233gat), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n574), .B(new_n571), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT97), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n583), .A2(new_n584), .A3(new_n561), .A4(new_n564), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n576), .A2(KEYINPUT97), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n562), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n581), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT99), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n582), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n583), .A2(new_n564), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n588), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n560), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT98), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n595), .A3(new_n581), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT98), .B1(new_n587), .B2(new_n588), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n593), .A2(new_n560), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  NOR3_X1   g400(.A1(new_n519), .A2(new_n557), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT100), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n354), .A2(new_n603), .A3(new_n355), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n603), .B1(new_n354), .B2(new_n355), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n484), .A2(new_n602), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(G1gat), .ZN(G1324gat));
  INV_X1    g408(.A(new_n328), .ZN(new_n610));
  INV_X1    g409(.A(new_n483), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n482), .B1(new_n400), .B2(new_n479), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n610), .B(new_n602), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT16), .B(G8gat), .Z(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n613), .A2(KEYINPUT42), .A3(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n613), .A2(new_n615), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT42), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n618), .B1(new_n613), .B2(G8gat), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n616), .B1(new_n617), .B2(new_n619), .ZN(G1325gat));
  NAND3_X1  g419(.A1(new_n484), .A2(new_n399), .A3(new_n602), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(G15gat), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n301), .A2(G15gat), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n484), .A2(new_n602), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(G1326gat));
  NAND3_X1  g424(.A1(new_n484), .A2(new_n246), .A3(new_n602), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT43), .B(G22gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(G1327gat));
  INV_X1    g427(.A(new_n601), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n519), .A2(new_n557), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT101), .Z(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n632), .B1(new_n481), .B2(new_n483), .ZN(new_n633));
  INV_X1    g432(.A(G29gat), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n633), .A2(new_n634), .A3(new_n607), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT45), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n633), .A2(KEYINPUT45), .A3(new_n634), .A4(new_n607), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n393), .A2(new_n367), .ZN(new_n639));
  INV_X1    g438(.A(new_n368), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n399), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n305), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n246), .A2(new_n301), .A3(new_n304), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n358), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n366), .B1(new_n644), .B2(KEYINPUT35), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n557), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n400), .A2(KEYINPUT44), .A3(new_n557), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n518), .B(KEYINPUT102), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(new_n479), .A3(new_n629), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT103), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n650), .A2(new_n607), .A3(new_n654), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n637), .B(new_n638), .C1(new_n634), .C2(new_n655), .ZN(G1328gat));
  NOR2_X1   g455(.A1(new_n328), .A2(G36gat), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n633), .A2(KEYINPUT46), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT46), .B1(new_n633), .B2(new_n657), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n650), .A2(new_n610), .A3(new_n654), .ZN(new_n660));
  INV_X1    g459(.A(G36gat), .ZN(new_n661));
  OAI22_X1  g460(.A1(new_n658), .A2(new_n659), .B1(new_n660), .B2(new_n661), .ZN(G1329gat));
  INV_X1    g461(.A(new_n301), .ZN(new_n663));
  AOI21_X1  g462(.A(G43gat), .B1(new_n633), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n398), .A2(new_n416), .ZN(new_n665));
  AND4_X1   g464(.A1(new_n648), .A2(new_n649), .A3(new_n654), .A4(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT47), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n663), .B(new_n631), .C1(new_n611), .C2(new_n612), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n416), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT47), .ZN(new_n670));
  INV_X1    g469(.A(new_n666), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n667), .A2(new_n672), .ZN(G1330gat));
  AOI21_X1  g472(.A(G50gat), .B1(new_n633), .B2(new_n246), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n367), .A2(new_n414), .ZN(new_n675));
  AND4_X1   g474(.A1(new_n648), .A2(new_n649), .A3(new_n654), .A4(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT48), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n246), .B(new_n631), .C1(new_n611), .C2(new_n612), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n414), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT48), .ZN(new_n680));
  INV_X1    g479(.A(new_n676), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n677), .A2(new_n682), .ZN(G1331gat));
  NAND2_X1  g482(.A1(new_n475), .A2(new_n455), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT90), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n469), .B1(new_n686), .B2(new_n476), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n518), .A2(new_n687), .A3(new_n556), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(new_n629), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n400), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n607), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g491(.A(new_n328), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT104), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n694), .B(new_n696), .ZN(G1333gat));
  NAND3_X1  g496(.A1(new_n690), .A2(KEYINPUT105), .A3(new_n663), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n400), .A2(new_n663), .A3(new_n689), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700));
  AOI21_X1  g499(.A(G71gat), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n690), .A2(G71gat), .A3(new_n399), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n246), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g506(.A1(new_n518), .A2(new_n479), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n557), .B(new_n708), .C1(new_n641), .C2(new_n645), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT51), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n400), .A2(KEYINPUT51), .A3(new_n557), .A4(new_n708), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n606), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n604), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(G85gat), .A3(new_n629), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT106), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n518), .A2(new_n479), .A3(new_n629), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n650), .A2(new_n607), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(new_n720), .B2(new_n526), .ZN(G1336gat));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n711), .A2(new_n712), .A3(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n328), .A2(G92gat), .A3(new_n629), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n709), .A2(KEYINPUT107), .A3(new_n710), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n648), .A2(new_n649), .A3(new_n610), .A4(new_n719), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G92gat), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT52), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT52), .B1(new_n713), .B2(new_n724), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n728), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(G1337gat));
  NAND3_X1  g532(.A1(new_n650), .A2(new_n399), .A3(new_n719), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G99gat), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n301), .A2(G99gat), .A3(new_n629), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT108), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n713), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n738), .ZN(G1338gat));
  NOR3_X1   g538(.A1(new_n367), .A2(G106gat), .A3(new_n629), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n723), .A2(new_n725), .A3(new_n740), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n648), .A2(new_n649), .A3(new_n246), .A4(new_n719), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G106gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT53), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT53), .B1(new_n713), .B2(new_n740), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1339gat));
  NOR2_X1   g547(.A1(new_n688), .A2(new_n601), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n452), .A2(new_n453), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n444), .B1(new_n436), .B2(new_n441), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n464), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n470), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n556), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT54), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n758), .B1(new_n587), .B2(new_n588), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n597), .A2(new_n596), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n582), .A2(new_n589), .A3(new_n758), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n560), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT109), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n762), .A2(new_n765), .A3(new_n560), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n761), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n760), .A2(KEYINPUT55), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n768), .B1(new_n764), .B2(new_n766), .ZN(new_n769));
  INV_X1    g568(.A(new_n600), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n769), .A2(KEYINPUT110), .A3(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n772));
  INV_X1    g571(.A(new_n768), .ZN(new_n773));
  INV_X1    g572(.A(new_n766), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n765), .B1(new_n762), .B2(new_n560), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n772), .B1(new_n776), .B2(new_n600), .ZN(new_n777));
  OAI221_X1 g576(.A(new_n757), .B1(KEYINPUT55), .B2(new_n767), .C1(new_n771), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n629), .A2(new_n756), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT110), .B1(new_n769), .B2(new_n770), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n776), .A2(new_n772), .A3(new_n600), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n760), .B1(new_n774), .B2(new_n775), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n687), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n779), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n778), .B1(new_n786), .B2(new_n557), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n749), .B1(new_n787), .B2(new_n652), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n788), .A2(new_n610), .A3(new_n715), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n789), .A2(new_n306), .ZN(new_n790));
  AOI21_X1  g589(.A(G113gat), .B1(new_n790), .B2(new_n479), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n302), .ZN(new_n792));
  INV_X1    g591(.A(G113gat), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n792), .A2(new_n793), .A3(new_n687), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT112), .ZN(G1340gat));
  NOR2_X1   g595(.A1(new_n629), .A2(G120gat), .ZN(new_n797));
  XOR2_X1   g596(.A(new_n797), .B(KEYINPUT113), .Z(new_n798));
  NAND2_X1  g597(.A1(new_n790), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(G120gat), .B1(new_n792), .B2(new_n629), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(G1341gat));
  INV_X1    g600(.A(G127gat), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n790), .A2(new_n802), .A3(new_n518), .ZN(new_n803));
  OAI21_X1  g602(.A(G127gat), .B1(new_n792), .B2(new_n652), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(G1342gat));
  NOR2_X1   g604(.A1(new_n788), .A2(new_n715), .ZN(new_n806));
  INV_X1    g605(.A(G134gat), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n610), .A2(new_n556), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n806), .A2(new_n807), .A3(new_n306), .A4(new_n808), .ZN(new_n809));
  XOR2_X1   g608(.A(new_n809), .B(KEYINPUT56), .Z(new_n810));
  NAND3_X1  g609(.A1(new_n789), .A2(new_n302), .A3(new_n557), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n811), .A2(KEYINPUT114), .A3(G134gat), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT114), .B1(new_n811), .B2(G134gat), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT115), .ZN(G1343gat));
  NOR3_X1   g614(.A1(new_n399), .A2(new_n610), .A3(new_n715), .ZN(new_n816));
  INV_X1    g615(.A(G141gat), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n687), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n246), .A2(KEYINPUT57), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n769), .A2(new_n770), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n779), .B1(new_n785), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(new_n557), .ZN(new_n822));
  XOR2_X1   g621(.A(new_n822), .B(KEYINPUT116), .Z(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n778), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n519), .ZN(new_n825));
  INV_X1    g624(.A(new_n749), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n819), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n785), .B1(new_n771), .B2(new_n777), .ZN(new_n828));
  INV_X1    g627(.A(new_n779), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n557), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n757), .B1(KEYINPUT55), .B2(new_n767), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n831), .B1(new_n780), .B2(new_n781), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n652), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n367), .B1(new_n833), .B2(new_n826), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(KEYINPUT57), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n816), .B(new_n818), .C1(new_n827), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n398), .A2(new_n246), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n789), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n817), .B1(new_n839), .B2(new_n687), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n836), .A2(KEYINPUT58), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT58), .B1(new_n836), .B2(new_n840), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI211_X1 g643(.A(KEYINPUT117), .B(KEYINPUT58), .C1(new_n836), .C2(new_n840), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n841), .B1(new_n844), .B2(new_n845), .ZN(G1344gat));
  INV_X1    g645(.A(new_n839), .ZN(new_n847));
  INV_X1    g646(.A(G148gat), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n847), .A2(new_n848), .A3(new_n601), .ZN(new_n849));
  INV_X1    g648(.A(new_n816), .ZN(new_n850));
  INV_X1    g649(.A(new_n827), .ZN(new_n851));
  INV_X1    g650(.A(new_n835), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI211_X1 g652(.A(KEYINPUT59), .B(new_n848), .C1(new_n853), .C2(new_n601), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n778), .B1(new_n821), .B2(new_n557), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n749), .B1(new_n857), .B2(new_n519), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n856), .B1(new_n858), .B2(new_n367), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n860), .B1(new_n834), .B2(KEYINPUT57), .ZN(new_n861));
  NOR4_X1   g660(.A1(new_n788), .A2(KEYINPUT118), .A3(new_n856), .A4(new_n367), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n601), .A3(new_n816), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n855), .B1(new_n864), .B2(G148gat), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n849), .B1(new_n854), .B2(new_n865), .ZN(G1345gat));
  INV_X1    g665(.A(G155gat), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n847), .A2(new_n867), .A3(new_n518), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n853), .A2(new_n651), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n868), .B1(new_n869), .B2(new_n867), .ZN(G1346gat));
  INV_X1    g669(.A(G162gat), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n806), .A2(new_n871), .A3(new_n808), .A4(new_n838), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT119), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n853), .A2(new_n557), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n871), .ZN(G1347gat));
  OAI21_X1  g674(.A(KEYINPUT120), .B1(new_n607), .B2(new_n328), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n715), .A2(new_n877), .A3(new_n610), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n876), .A2(new_n302), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n833), .A2(new_n826), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n881), .A2(new_n460), .A3(new_n687), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n788), .A2(new_n607), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n328), .B1(new_n303), .B2(new_n305), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n479), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n882), .B1(new_n887), .B2(new_n460), .ZN(G1348gat));
  AOI21_X1  g687(.A(G176gat), .B1(new_n886), .B2(new_n601), .ZN(new_n889));
  INV_X1    g688(.A(G176gat), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n881), .A2(new_n890), .A3(new_n629), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n891), .A2(KEYINPUT121), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(KEYINPUT121), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(G1349gat));
  OAI21_X1  g693(.A(G183gat), .B1(new_n881), .B2(new_n652), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n518), .A2(new_n263), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n885), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g697(.A1(new_n886), .A2(new_n264), .A3(new_n557), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n879), .A2(new_n880), .A3(new_n557), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n900), .A2(new_n901), .A3(G190gat), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n900), .B2(G190gat), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(G1351gat));
  NOR2_X1   g703(.A1(new_n837), .A2(new_n328), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n883), .A2(new_n905), .ZN(new_n906));
  XOR2_X1   g705(.A(KEYINPUT122), .B(G197gat), .Z(new_n907));
  NOR3_X1   g706(.A1(new_n906), .A2(new_n687), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT123), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n876), .A2(new_n398), .A3(new_n878), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n910), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n479), .B1(new_n767), .B2(KEYINPUT55), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n913), .B1(new_n780), .B2(new_n781), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n556), .B1(new_n914), .B2(new_n779), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n651), .B1(new_n915), .B2(new_n778), .ZN(new_n916));
  OAI211_X1 g715(.A(KEYINPUT57), .B(new_n246), .C1(new_n916), .C2(new_n749), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT118), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n880), .A2(new_n860), .A3(KEYINPUT57), .A4(new_n246), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n912), .B1(new_n920), .B2(new_n859), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(KEYINPUT125), .A3(new_n479), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n907), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT125), .B1(new_n921), .B2(new_n479), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n909), .B1(new_n923), .B2(new_n924), .ZN(G1352gat));
  NOR3_X1   g724(.A1(new_n906), .A2(G204gat), .A3(new_n629), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT62), .ZN(new_n927));
  INV_X1    g726(.A(G204gat), .ZN(new_n928));
  AOI211_X1 g727(.A(new_n629), .B(new_n912), .C1(new_n920), .C2(new_n859), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(G1353gat));
  INV_X1    g729(.A(new_n906), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n216), .A3(new_n518), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n933));
  AOI211_X1 g732(.A(new_n933), .B(new_n216), .C1(new_n921), .C2(new_n518), .ZN(new_n934));
  INV_X1    g733(.A(new_n912), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n863), .A2(new_n518), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n932), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT126), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n940), .B(new_n932), .C1(new_n934), .C2(new_n937), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1354gat));
  AOI21_X1  g741(.A(G218gat), .B1(new_n931), .B2(new_n557), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n921), .B(KEYINPUT127), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n556), .A2(new_n215), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(G1355gat));
endmodule


