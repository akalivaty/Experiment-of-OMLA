

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595;

  NAND2_X1 U322 ( .A1(n390), .A2(n389), .ZN(n392) );
  NOR2_X1 U323 ( .A1(n552), .A2(n478), .ZN(n592) );
  XNOR2_X1 U324 ( .A(n454), .B(n453), .ZN(n507) );
  NOR2_X1 U325 ( .A1(n580), .A2(n579), .ZN(n290) );
  XOR2_X1 U326 ( .A(G43GAT), .B(G99GAT), .Z(n291) );
  XOR2_X1 U327 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n292) );
  NOR2_X1 U328 ( .A1(n579), .A2(n525), .ZN(n365) );
  XNOR2_X1 U329 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n473) );
  XNOR2_X1 U330 ( .A(KEYINPUT54), .B(KEYINPUT122), .ZN(n475) );
  XNOR2_X1 U331 ( .A(n474), .B(n473), .ZN(n532) );
  INV_X1 U332 ( .A(KEYINPUT97), .ZN(n391) );
  XNOR2_X1 U333 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U334 ( .A(n392), .B(n391), .ZN(n486) );
  XNOR2_X1 U335 ( .A(n346), .B(n291), .ZN(n347) );
  XNOR2_X1 U336 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U337 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U338 ( .A(n410), .B(n409), .ZN(n417) );
  INV_X1 U339 ( .A(G204GAT), .ZN(n480) );
  INV_X1 U340 ( .A(G29GAT), .ZN(n455) );
  XNOR2_X1 U341 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U342 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U343 ( .A(n483), .B(n482), .ZN(G1353GAT) );
  XNOR2_X1 U344 ( .A(n458), .B(n457), .ZN(G1328GAT) );
  XOR2_X1 U345 ( .A(G113GAT), .B(G1GAT), .Z(n432) );
  XOR2_X1 U346 ( .A(G148GAT), .B(G134GAT), .Z(n294) );
  XNOR2_X1 U347 ( .A(G29GAT), .B(G85GAT), .ZN(n293) );
  XNOR2_X1 U348 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U349 ( .A(n432), .B(n295), .Z(n297) );
  NAND2_X1 U350 ( .A1(G225GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U351 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U352 ( .A(n298), .B(KEYINPUT90), .Z(n301) );
  XNOR2_X1 U353 ( .A(G120GAT), .B(KEYINPUT0), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n299), .B(KEYINPUT81), .ZN(n336) );
  XNOR2_X1 U355 ( .A(n336), .B(KEYINPUT5), .ZN(n300) );
  XNOR2_X1 U356 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U357 ( .A(KEYINPUT6), .B(G57GAT), .Z(n303) );
  XNOR2_X1 U358 ( .A(G141GAT), .B(G127GAT), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U360 ( .A(n305), .B(n304), .Z(n314) );
  XNOR2_X1 U361 ( .A(KEYINPUT3), .B(KEYINPUT87), .ZN(n306) );
  XNOR2_X1 U362 ( .A(n306), .B(KEYINPUT2), .ZN(n307) );
  XOR2_X1 U363 ( .A(n307), .B(KEYINPUT88), .Z(n309) );
  XNOR2_X1 U364 ( .A(G155GAT), .B(G162GAT), .ZN(n308) );
  XNOR2_X1 U365 ( .A(n309), .B(n308), .ZN(n367) );
  XOR2_X1 U366 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n311) );
  XNOR2_X1 U367 ( .A(KEYINPUT4), .B(KEYINPUT1), .ZN(n310) );
  XNOR2_X1 U368 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n367), .B(n312), .ZN(n313) );
  XOR2_X1 U370 ( .A(n314), .B(n313), .Z(n490) );
  INV_X1 U371 ( .A(n490), .ZN(n535) );
  XOR2_X1 U372 ( .A(KEYINPUT105), .B(KEYINPUT38), .Z(n454) );
  XOR2_X1 U373 ( .A(G211GAT), .B(G22GAT), .Z(n316) );
  XNOR2_X1 U374 ( .A(G155GAT), .B(G78GAT), .ZN(n315) );
  XNOR2_X1 U375 ( .A(n316), .B(n315), .ZN(n329) );
  XOR2_X1 U376 ( .A(G8GAT), .B(G64GAT), .Z(n318) );
  XNOR2_X1 U377 ( .A(G1GAT), .B(G183GAT), .ZN(n317) );
  XNOR2_X1 U378 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U379 ( .A(KEYINPUT80), .B(KEYINPUT12), .Z(n320) );
  XNOR2_X1 U380 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n319) );
  XNOR2_X1 U381 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U382 ( .A(n322), .B(n321), .ZN(n327) );
  XOR2_X1 U383 ( .A(G127GAT), .B(G15GAT), .Z(n343) );
  XNOR2_X1 U384 ( .A(G57GAT), .B(G71GAT), .ZN(n323) );
  XNOR2_X1 U385 ( .A(n323), .B(KEYINPUT13), .ZN(n447) );
  XOR2_X1 U386 ( .A(n343), .B(n447), .Z(n325) );
  NAND2_X1 U387 ( .A1(G231GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U388 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U390 ( .A(n329), .B(n328), .Z(n577) );
  INV_X1 U391 ( .A(n577), .ZN(n590) );
  XOR2_X1 U392 ( .A(G169GAT), .B(G176GAT), .Z(n331) );
  XNOR2_X1 U393 ( .A(G113GAT), .B(KEYINPUT85), .ZN(n330) );
  XNOR2_X1 U394 ( .A(n331), .B(n330), .ZN(n350) );
  XOR2_X1 U395 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n333) );
  NAND2_X1 U396 ( .A1(G227GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U397 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U398 ( .A(n334), .B(KEYINPUT83), .Z(n338) );
  XNOR2_X1 U399 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n292), .B(n335), .ZN(n354) );
  XNOR2_X1 U401 ( .A(n336), .B(n354), .ZN(n337) );
  XNOR2_X1 U402 ( .A(n338), .B(n337), .ZN(n348) );
  XOR2_X1 U403 ( .A(KEYINPUT84), .B(G71GAT), .Z(n345) );
  INV_X1 U404 ( .A(G190GAT), .ZN(n339) );
  NAND2_X1 U405 ( .A1(G134GAT), .A2(n339), .ZN(n342) );
  INV_X1 U406 ( .A(G134GAT), .ZN(n340) );
  NAND2_X1 U407 ( .A1(n340), .A2(G190GAT), .ZN(n341) );
  NAND2_X1 U408 ( .A1(n342), .A2(n341), .ZN(n396) );
  XNOR2_X1 U409 ( .A(n396), .B(n343), .ZN(n344) );
  XNOR2_X1 U410 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n567) );
  INV_X1 U412 ( .A(n567), .ZN(n579) );
  XOR2_X1 U413 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n356) );
  XOR2_X1 U414 ( .A(G190GAT), .B(G36GAT), .Z(n352) );
  NAND2_X1 U415 ( .A1(G226GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n358) );
  XNOR2_X1 U419 ( .A(G92GAT), .B(G64GAT), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n357), .B(G176GAT), .ZN(n446) );
  XOR2_X1 U421 ( .A(n358), .B(n446), .Z(n364) );
  XOR2_X1 U422 ( .A(KEYINPUT86), .B(G204GAT), .Z(n360) );
  XNOR2_X1 U423 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U425 ( .A(G211GAT), .B(n361), .Z(n366) );
  XNOR2_X1 U426 ( .A(G8GAT), .B(G169GAT), .ZN(n362) );
  XNOR2_X1 U427 ( .A(n362), .B(G197GAT), .ZN(n426) );
  XNOR2_X1 U428 ( .A(n366), .B(n426), .ZN(n363) );
  XOR2_X1 U429 ( .A(n364), .B(n363), .Z(n495) );
  INV_X1 U430 ( .A(n495), .ZN(n525) );
  XNOR2_X1 U431 ( .A(KEYINPUT95), .B(n365), .ZN(n379) );
  XNOR2_X1 U432 ( .A(n367), .B(n366), .ZN(n378) );
  XOR2_X1 U433 ( .A(G141GAT), .B(G22GAT), .Z(n431) );
  XOR2_X1 U434 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n369) );
  XNOR2_X1 U435 ( .A(G50GAT), .B(KEYINPUT89), .ZN(n368) );
  XNOR2_X1 U436 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U437 ( .A(n431), .B(n370), .Z(n372) );
  NAND2_X1 U438 ( .A1(G228GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U439 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U440 ( .A(n373), .B(KEYINPUT22), .Z(n376) );
  XNOR2_X1 U441 ( .A(G148GAT), .B(G106GAT), .ZN(n374) );
  XNOR2_X1 U442 ( .A(n374), .B(G78GAT), .ZN(n439) );
  XNOR2_X1 U443 ( .A(G197GAT), .B(n439), .ZN(n375) );
  XNOR2_X1 U444 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n378), .B(n377), .ZN(n565) );
  NAND2_X1 U446 ( .A1(n379), .A2(n565), .ZN(n380) );
  XNOR2_X1 U447 ( .A(n380), .B(KEYINPUT25), .ZN(n383) );
  XOR2_X1 U448 ( .A(n495), .B(KEYINPUT27), .Z(n386) );
  OR2_X1 U449 ( .A1(n565), .A2(n567), .ZN(n381) );
  XNOR2_X1 U450 ( .A(n381), .B(KEYINPUT26), .ZN(n552) );
  NOR2_X1 U451 ( .A1(n386), .A2(n552), .ZN(n382) );
  NOR2_X1 U452 ( .A1(n383), .A2(n382), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n384), .B(KEYINPUT96), .ZN(n385) );
  NAND2_X1 U454 ( .A1(n385), .A2(n535), .ZN(n390) );
  INV_X1 U455 ( .A(n386), .ZN(n533) );
  XOR2_X1 U456 ( .A(KEYINPUT28), .B(n565), .Z(n537) );
  NOR2_X1 U457 ( .A1(n537), .A2(n567), .ZN(n387) );
  NAND2_X1 U458 ( .A1(n533), .A2(n387), .ZN(n388) );
  NAND2_X1 U459 ( .A1(n490), .A2(n388), .ZN(n389) );
  NOR2_X1 U460 ( .A1(n590), .A2(n486), .ZN(n393) );
  XNOR2_X1 U461 ( .A(n393), .B(KEYINPUT104), .ZN(n418) );
  XOR2_X1 U462 ( .A(KEYINPUT10), .B(G92GAT), .Z(n400) );
  XNOR2_X1 U463 ( .A(G85GAT), .B(G99GAT), .ZN(n395) );
  INV_X1 U464 ( .A(n396), .ZN(n394) );
  NAND2_X1 U465 ( .A1(n395), .A2(n394), .ZN(n398) );
  INV_X1 U466 ( .A(n395), .ZN(n437) );
  NAND2_X1 U467 ( .A1(n437), .A2(n396), .ZN(n397) );
  NAND2_X1 U468 ( .A1(n398), .A2(n397), .ZN(n399) );
  XNOR2_X1 U469 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U470 ( .A(n401), .B(G106GAT), .Z(n410) );
  XOR2_X1 U471 ( .A(KEYINPUT9), .B(KEYINPUT65), .Z(n403) );
  XNOR2_X1 U472 ( .A(KEYINPUT11), .B(KEYINPUT78), .ZN(n402) );
  XNOR2_X1 U473 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U474 ( .A(n404), .B(G218GAT), .ZN(n408) );
  XOR2_X1 U475 ( .A(KEYINPUT79), .B(KEYINPUT77), .Z(n406) );
  NAND2_X1 U476 ( .A1(G232GAT), .A2(G233GAT), .ZN(n405) );
  XOR2_X1 U477 ( .A(n406), .B(n405), .Z(n407) );
  XOR2_X1 U478 ( .A(G50GAT), .B(KEYINPUT8), .Z(n412) );
  XNOR2_X1 U479 ( .A(KEYINPUT7), .B(KEYINPUT70), .ZN(n411) );
  XNOR2_X1 U480 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U481 ( .A(n413), .B(G43GAT), .Z(n415) );
  XNOR2_X1 U482 ( .A(G29GAT), .B(G36GAT), .ZN(n414) );
  XNOR2_X1 U483 ( .A(n415), .B(n414), .ZN(n423) );
  XNOR2_X1 U484 ( .A(G162GAT), .B(n423), .ZN(n416) );
  XOR2_X1 U485 ( .A(n417), .B(n416), .Z(n580) );
  XOR2_X1 U486 ( .A(KEYINPUT36), .B(n580), .Z(n593) );
  NAND2_X1 U487 ( .A1(n418), .A2(n593), .ZN(n419) );
  XNOR2_X1 U488 ( .A(n419), .B(KEYINPUT37), .ZN(n522) );
  XOR2_X1 U489 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n421) );
  XNOR2_X1 U490 ( .A(KEYINPUT69), .B(KEYINPUT30), .ZN(n420) );
  XNOR2_X1 U491 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U492 ( .A(n423), .B(n422), .ZN(n436) );
  XOR2_X1 U493 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n425) );
  XNOR2_X1 U494 ( .A(G15GAT), .B(KEYINPUT72), .ZN(n424) );
  XNOR2_X1 U495 ( .A(n425), .B(n424), .ZN(n430) );
  XOR2_X1 U496 ( .A(n426), .B(KEYINPUT71), .Z(n428) );
  NAND2_X1 U497 ( .A1(G229GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U498 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U499 ( .A(n430), .B(n429), .Z(n434) );
  XNOR2_X1 U500 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U501 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U502 ( .A(n436), .B(n435), .ZN(n585) );
  XNOR2_X1 U503 ( .A(KEYINPUT73), .B(n585), .ZN(n568) );
  XNOR2_X1 U504 ( .A(G120GAT), .B(G204GAT), .ZN(n438) );
  XOR2_X1 U505 ( .A(n438), .B(n437), .Z(n451) );
  XOR2_X1 U506 ( .A(KEYINPUT33), .B(n439), .Z(n441) );
  NAND2_X1 U507 ( .A1(G230GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U508 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U509 ( .A(KEYINPUT32), .B(KEYINPUT75), .Z(n443) );
  XNOR2_X1 U510 ( .A(KEYINPUT74), .B(KEYINPUT31), .ZN(n442) );
  XNOR2_X1 U511 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U512 ( .A(n445), .B(n444), .Z(n449) );
  XNOR2_X1 U513 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U514 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U515 ( .A(n451), .B(n450), .ZN(n479) );
  NOR2_X1 U516 ( .A1(n568), .A2(n479), .ZN(n452) );
  XNOR2_X1 U517 ( .A(n452), .B(KEYINPUT76), .ZN(n488) );
  NAND2_X1 U518 ( .A1(n522), .A2(n488), .ZN(n453) );
  NOR2_X1 U519 ( .A1(n535), .A2(n507), .ZN(n458) );
  XNOR2_X1 U520 ( .A(KEYINPUT103), .B(KEYINPUT39), .ZN(n456) );
  NAND2_X1 U521 ( .A1(n593), .A2(n590), .ZN(n459) );
  XOR2_X1 U522 ( .A(KEYINPUT45), .B(n459), .Z(n460) );
  NAND2_X1 U523 ( .A1(n460), .A2(n568), .ZN(n461) );
  NOR2_X1 U524 ( .A1(n479), .A2(n461), .ZN(n462) );
  XNOR2_X1 U525 ( .A(KEYINPUT113), .B(n462), .ZN(n472) );
  INV_X1 U526 ( .A(n580), .ZN(n561) );
  XNOR2_X1 U527 ( .A(n479), .B(KEYINPUT64), .ZN(n464) );
  INV_X1 U528 ( .A(KEYINPUT41), .ZN(n463) );
  XNOR2_X1 U529 ( .A(n464), .B(n463), .ZN(n510) );
  NAND2_X1 U530 ( .A1(n585), .A2(n510), .ZN(n466) );
  INV_X1 U531 ( .A(KEYINPUT46), .ZN(n465) );
  XOR2_X1 U532 ( .A(n466), .B(n465), .Z(n467) );
  NAND2_X1 U533 ( .A1(n467), .A2(n577), .ZN(n468) );
  NOR2_X1 U534 ( .A1(n561), .A2(n468), .ZN(n470) );
  XNOR2_X1 U535 ( .A(KEYINPUT47), .B(KEYINPUT112), .ZN(n469) );
  XNOR2_X1 U536 ( .A(n470), .B(n469), .ZN(n471) );
  NAND2_X1 U537 ( .A1(n472), .A2(n471), .ZN(n474) );
  NAND2_X1 U538 ( .A1(n532), .A2(n495), .ZN(n476) );
  NOR2_X1 U539 ( .A1(n490), .A2(n477), .ZN(n564) );
  INV_X1 U540 ( .A(n564), .ZN(n478) );
  NAND2_X1 U541 ( .A1(n592), .A2(n479), .ZN(n483) );
  XOR2_X1 U542 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n481) );
  XNOR2_X1 U543 ( .A(KEYINPUT101), .B(KEYINPUT100), .ZN(n494) );
  XOR2_X1 U544 ( .A(G1GAT), .B(KEYINPUT34), .Z(n492) );
  NOR2_X1 U545 ( .A1(n561), .A2(n577), .ZN(n484) );
  XOR2_X1 U546 ( .A(KEYINPUT16), .B(n484), .Z(n485) );
  NOR2_X1 U547 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U548 ( .A(KEYINPUT98), .B(n487), .ZN(n512) );
  NAND2_X1 U549 ( .A1(n488), .A2(n512), .ZN(n489) );
  XNOR2_X1 U550 ( .A(KEYINPUT99), .B(n489), .ZN(n500) );
  NAND2_X1 U551 ( .A1(n500), .A2(n490), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(G1324GAT) );
  NAND2_X1 U554 ( .A1(n500), .A2(n495), .ZN(n496) );
  XNOR2_X1 U555 ( .A(G8GAT), .B(n496), .ZN(G1325GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT35), .B(KEYINPUT102), .Z(n498) );
  NAND2_X1 U557 ( .A1(n500), .A2(n567), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U559 ( .A(G15GAT), .B(n499), .ZN(G1326GAT) );
  NAND2_X1 U560 ( .A1(n500), .A2(n537), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n501), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U562 ( .A1(n525), .A2(n507), .ZN(n502) );
  XOR2_X1 U563 ( .A(KEYINPUT106), .B(n502), .Z(n503) );
  XNOR2_X1 U564 ( .A(G36GAT), .B(n503), .ZN(G1329GAT) );
  XNOR2_X1 U565 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n505) );
  NOR2_X1 U566 ( .A1(n579), .A2(n507), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U568 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  INV_X1 U569 ( .A(n537), .ZN(n529) );
  NOR2_X1 U570 ( .A1(n507), .A2(n529), .ZN(n508) );
  XOR2_X1 U571 ( .A(G50GAT), .B(n508), .Z(n509) );
  XNOR2_X1 U572 ( .A(KEYINPUT108), .B(n509), .ZN(G1331GAT) );
  INV_X1 U573 ( .A(n510), .ZN(n573) );
  NOR2_X1 U574 ( .A1(n585), .A2(n573), .ZN(n511) );
  XOR2_X1 U575 ( .A(KEYINPUT109), .B(n511), .Z(n521) );
  NAND2_X1 U576 ( .A1(n521), .A2(n512), .ZN(n518) );
  NOR2_X1 U577 ( .A1(n535), .A2(n518), .ZN(n513) );
  XOR2_X1 U578 ( .A(G57GAT), .B(n513), .Z(n514) );
  XNOR2_X1 U579 ( .A(KEYINPUT42), .B(n514), .ZN(G1332GAT) );
  NOR2_X1 U580 ( .A1(n525), .A2(n518), .ZN(n515) );
  XOR2_X1 U581 ( .A(KEYINPUT110), .B(n515), .Z(n516) );
  XNOR2_X1 U582 ( .A(G64GAT), .B(n516), .ZN(G1333GAT) );
  NOR2_X1 U583 ( .A1(n579), .A2(n518), .ZN(n517) );
  XOR2_X1 U584 ( .A(G71GAT), .B(n517), .Z(G1334GAT) );
  NOR2_X1 U585 ( .A1(n529), .A2(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NAND2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n528) );
  NOR2_X1 U589 ( .A1(n535), .A2(n528), .ZN(n524) );
  XNOR2_X1 U590 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n524), .B(n523), .ZN(G1336GAT) );
  NOR2_X1 U592 ( .A1(n525), .A2(n528), .ZN(n526) );
  XOR2_X1 U593 ( .A(G92GAT), .B(n526), .Z(G1337GAT) );
  NOR2_X1 U594 ( .A1(n579), .A2(n528), .ZN(n527) );
  XOR2_X1 U595 ( .A(G99GAT), .B(n527), .Z(G1338GAT) );
  NOR2_X1 U596 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U597 ( .A(KEYINPUT44), .B(n530), .Z(n531) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NAND2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U601 ( .A(KEYINPUT115), .B(n536), .ZN(n551) );
  INV_X1 U602 ( .A(n551), .ZN(n539) );
  NOR2_X1 U603 ( .A1(n579), .A2(n537), .ZN(n538) );
  NAND2_X1 U604 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U605 ( .A(KEYINPUT116), .B(n540), .ZN(n548) );
  NOR2_X1 U606 ( .A1(n548), .A2(n568), .ZN(n542) );
  XNOR2_X1 U607 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G113GAT), .B(n543), .ZN(G1340GAT) );
  XNOR2_X1 U610 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n545) );
  NOR2_X1 U611 ( .A1(n573), .A2(n548), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  NOR2_X1 U613 ( .A1(n577), .A2(n548), .ZN(n546) );
  XOR2_X1 U614 ( .A(KEYINPUT50), .B(n546), .Z(n547) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  NOR2_X1 U616 ( .A1(n548), .A2(n580), .ZN(n550) );
  XNOR2_X1 U617 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  XOR2_X1 U619 ( .A(G141GAT), .B(KEYINPUT119), .Z(n554) );
  NOR2_X1 U620 ( .A1(n552), .A2(n551), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n562), .A2(n585), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n556) );
  NAND2_X1 U624 ( .A1(n562), .A2(n510), .ZN(n555) );
  XNOR2_X1 U625 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(n557), .ZN(G1345GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n559) );
  NAND2_X1 U628 ( .A1(n562), .A2(n590), .ZN(n558) );
  XNOR2_X1 U629 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U630 ( .A(G155GAT), .B(n560), .ZN(G1346GAT) );
  NAND2_X1 U631 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n563), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U633 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n566), .B(KEYINPUT55), .ZN(n581) );
  NAND2_X1 U635 ( .A1(n581), .A2(n567), .ZN(n576) );
  NOR2_X1 U636 ( .A1(n568), .A2(n576), .ZN(n570) );
  XNOR2_X1 U637 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n569) );
  XNOR2_X1 U638 ( .A(n570), .B(n569), .ZN(G1348GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT124), .B(KEYINPUT57), .Z(n572) );
  XNOR2_X1 U640 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n571) );
  XNOR2_X1 U641 ( .A(n572), .B(n571), .ZN(n575) );
  NOR2_X1 U642 ( .A1(n573), .A2(n576), .ZN(n574) );
  XOR2_X1 U643 ( .A(n575), .B(n574), .Z(G1349GAT) );
  NOR2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U645 ( .A(G183GAT), .B(n578), .Z(G1350GAT) );
  AND2_X1 U646 ( .A1(n581), .A2(n290), .ZN(n583) );
  XNOR2_X1 U647 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(G190GAT), .B(n584), .ZN(G1351GAT) );
  NAND2_X1 U650 ( .A1(n592), .A2(n585), .ZN(n589) );
  XOR2_X1 U651 ( .A(KEYINPUT126), .B(KEYINPUT59), .Z(n587) );
  XNOR2_X1 U652 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1352GAT) );
  NAND2_X1 U655 ( .A1(n590), .A2(n592), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n591), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(n594), .B(KEYINPUT62), .ZN(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

