//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352, new_n1353;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n202), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0003(.A(KEYINPUT65), .ZN(new_n204));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  OAI21_X1  g0005(.A(new_n204), .B1(new_n205), .B2(G13), .ZN(new_n206));
  INV_X1    g0006(.A(G13), .ZN(new_n207));
  NAND4_X1  g0007(.A1(new_n207), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  OAI21_X1  g0010(.A(G250), .B1(G257), .B2(G264), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(new_n212), .A2(KEYINPUT0), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n221), .B1(KEYINPUT0), .B2(new_n212), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT66), .Z(new_n223));
  NAND2_X1  g0023(.A1(G116), .A2(G270), .ZN(new_n224));
  INV_X1    g0024(.A(G50), .ZN(new_n225));
  INV_X1    g0025(.A(G226), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(G77), .B2(G244), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n229), .A2(new_n230), .A3(KEYINPUT68), .ZN(new_n231));
  INV_X1    g0031(.A(G238), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT67), .B(G68), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n228), .B(new_n231), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(KEYINPUT68), .B1(new_n229), .B2(new_n230), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n205), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT1), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n223), .A2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT2), .B(G226), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G264), .B(G270), .Z(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT69), .ZN(new_n249));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  OR2_X1    g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n259), .A2(G223), .B1(new_n262), .B2(G77), .ZN(new_n263));
  INV_X1    g0063(.A(G222), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT3), .B(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n256), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(G1), .A2(G13), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G274), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n268), .B2(new_n269), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G41), .A2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n274), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  OR2_X1    g0078(.A1(KEYINPUT70), .A2(G1), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT70), .A2(G1), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n270), .B1(new_n281), .B2(new_n276), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n278), .B1(new_n283), .B2(G226), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n272), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT71), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n272), .A2(KEYINPUT71), .A3(new_n284), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G190), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(G200), .A3(new_n288), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n225), .A2(new_n216), .A3(new_n217), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n292), .A2(G20), .B1(G150), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT72), .ZN(new_n295));
  INV_X1    g0095(.A(G33), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n295), .B1(new_n296), .B2(G20), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n214), .A2(KEYINPUT72), .A3(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT8), .B(G58), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n294), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n213), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n279), .A2(G13), .A3(G20), .A4(new_n280), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n301), .A2(new_n303), .B1(new_n225), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n303), .ZN(new_n307));
  AND2_X1   g0107(.A1(KEYINPUT70), .A2(G1), .ZN(new_n308));
  NOR2_X1   g0108(.A1(KEYINPUT70), .A2(G1), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G20), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n307), .A2(G50), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT9), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n290), .A2(new_n291), .A3(new_n314), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n315), .A2(KEYINPUT10), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(KEYINPUT10), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G179), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n289), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n287), .A2(new_n321), .A3(new_n288), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n313), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n259), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n265), .A2(G223), .A3(new_n256), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n271), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n278), .B1(new_n283), .B2(G232), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G169), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n319), .B2(new_n330), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT16), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n218), .B1(new_n233), .B2(new_n216), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G20), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n293), .A2(G159), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT7), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n265), .B2(G20), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n262), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n233), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n333), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  NOR3_X1   g0142(.A1(new_n265), .A2(new_n338), .A3(G20), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT7), .B1(new_n262), .B2(new_n214), .ZN(new_n344));
  OAI21_X1  g0144(.A(G68), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n345), .A2(KEYINPUT16), .A3(new_n335), .A4(new_n336), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n342), .A2(new_n346), .A3(new_n303), .ZN(new_n347));
  NOR3_X1   g0147(.A1(new_n308), .A2(new_n309), .A3(new_n214), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(new_n300), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n307), .A2(new_n349), .B1(new_n305), .B2(new_n300), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n332), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT18), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n330), .A2(G200), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n328), .A2(new_n329), .A3(G190), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n356), .A2(KEYINPUT17), .A3(new_n347), .A4(new_n350), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT18), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n332), .A2(new_n351), .A3(new_n358), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n347), .A2(new_n354), .A3(new_n350), .A4(new_n355), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT17), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n353), .A2(new_n357), .A3(new_n359), .A4(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NOR4_X1   g0164(.A1(new_n305), .A2(new_n348), .A3(new_n217), .A4(new_n303), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT12), .B1(new_n305), .B2(new_n217), .ZN(new_n366));
  INV_X1    g0166(.A(new_n233), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT12), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n367), .A2(new_n304), .A3(new_n368), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n365), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n233), .A2(G20), .B1(G50), .B2(new_n293), .ZN(new_n371));
  INV_X1    g0171(.A(G77), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n372), .B2(new_n299), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n303), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT11), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n373), .A2(KEYINPUT11), .A3(new_n303), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n370), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n274), .A2(new_n275), .A3(new_n277), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n282), .B2(new_n232), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n240), .A2(G1698), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n265), .B(new_n383), .C1(G226), .C2(G1698), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G33), .A2(G97), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n271), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT13), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n382), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n270), .B1(new_n384), .B2(new_n385), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT13), .B1(new_n390), .B2(new_n381), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n321), .B1(new_n389), .B2(new_n391), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT14), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n393), .A2(G179), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n394), .A2(new_n395), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n379), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G200), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G190), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n392), .A2(new_n401), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n400), .A2(new_n378), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n300), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n405), .A2(new_n293), .B1(G20), .B2(G77), .ZN(new_n406));
  XNOR2_X1  g0206(.A(KEYINPUT15), .B(G87), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n406), .B1(new_n299), .B2(new_n407), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(new_n303), .B1(new_n372), .B2(new_n305), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n307), .A2(G77), .A3(new_n311), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G244), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n380), .B1(new_n282), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n259), .A2(G238), .ZN(new_n414));
  INV_X1    g0214(.A(G107), .ZN(new_n415));
  OAI221_X1 g0215(.A(new_n414), .B1(new_n415), .B2(new_n265), .C1(new_n240), .C2(new_n266), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n413), .B1(new_n416), .B2(new_n271), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n411), .B1(G190), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n417), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G200), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n321), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n417), .A2(new_n319), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n411), .A3(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n364), .A2(new_n404), .A3(new_n421), .A4(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n324), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n348), .A2(G13), .A3(new_n415), .A4(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n427), .B1(new_n304), .B2(G107), .ZN(new_n430));
  NAND2_X1  g0230(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n279), .A2(G33), .A3(new_n280), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n302), .A2(new_n213), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n304), .A2(new_n433), .A3(new_n434), .A4(G107), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n432), .A2(KEYINPUT81), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT81), .B1(new_n432), .B2(new_n435), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n214), .B(G87), .C1(new_n260), .C2(new_n261), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT22), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT22), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n265), .A2(new_n441), .A3(new_n214), .A4(G87), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT23), .B1(new_n214), .B2(G107), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT23), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n445), .A2(new_n415), .A3(G20), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  OR2_X1    g0247(.A1(KEYINPUT77), .A2(G116), .ZN(new_n448));
  NAND2_X1  g0248(.A1(KEYINPUT77), .A2(G116), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n296), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n447), .B1(new_n450), .B2(new_n214), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n443), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT24), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n443), .A2(KEYINPUT24), .A3(new_n451), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n454), .A2(new_n303), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT82), .B1(new_n438), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n432), .A2(new_n435), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT81), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n432), .A2(KEYINPUT81), .A3(new_n435), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT82), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n434), .B1(new_n452), .B2(new_n453), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n455), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G294), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n467), .A2(KEYINPUT83), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(KEYINPUT83), .ZN(new_n469));
  OAI21_X1  g0269(.A(G33), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(G257), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n471));
  OAI211_X1 g0271(.A(G250), .B(new_n256), .C1(new_n260), .C2(new_n261), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n271), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT5), .B(G41), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n274), .A2(new_n310), .A3(new_n475), .A4(G45), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n310), .A2(new_n475), .A3(G45), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(G264), .A3(new_n270), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G169), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n319), .B2(new_n479), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n457), .A2(new_n466), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n399), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n474), .A2(new_n401), .A3(new_n476), .A4(new_n478), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n483), .A2(KEYINPUT84), .A3(new_n484), .ZN(new_n485));
  OR2_X1    g0285(.A1(new_n484), .A2(KEYINPUT84), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n485), .A2(new_n462), .A3(new_n486), .A4(new_n465), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(G20), .B1(G33), .B2(G283), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n296), .A2(G97), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n448), .A2(new_n449), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n303), .B(new_n491), .C1(new_n492), .C2(new_n214), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT20), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n449), .ZN(new_n496));
  NOR2_X1   g0296(.A1(KEYINPUT77), .A2(G116), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G20), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n489), .A2(new_n490), .B1(new_n302), .B2(new_n213), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(KEYINPUT20), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n304), .A2(new_n433), .A3(new_n434), .A4(G116), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n305), .A2(new_n498), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n477), .A2(G270), .A3(new_n270), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n476), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n265), .A2(G264), .A3(G1698), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n265), .A2(G257), .A3(new_n256), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n262), .A2(G303), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT79), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT79), .A4(new_n510), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n507), .B1(new_n515), .B2(new_n271), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n505), .B1(new_n517), .B2(G200), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n401), .B2(new_n517), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n515), .A2(new_n271), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n507), .A2(new_n319), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n520), .A2(new_n505), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n505), .A2(G169), .ZN(new_n523));
  OAI21_X1  g0323(.A(KEYINPUT21), .B1(new_n516), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n495), .A2(new_n501), .B1(new_n305), .B2(new_n498), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n321), .B1(new_n525), .B2(new_n503), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT21), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n270), .B1(new_n513), .B2(new_n514), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n526), .B(new_n527), .C1(new_n507), .C2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n522), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n519), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n293), .A2(G77), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT6), .ZN(new_n533));
  INV_X1    g0333(.A(G97), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n533), .A2(new_n534), .A3(G107), .ZN(new_n535));
  XNOR2_X1  g0335(.A(G97), .B(G107), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n535), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n532), .B1(new_n537), .B2(new_n214), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n415), .B1(new_n339), .B2(new_n340), .ZN(new_n539));
  OR2_X1    g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT73), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n348), .A2(new_n541), .A3(G13), .A4(new_n534), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT73), .B1(new_n304), .B2(G97), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n304), .A2(new_n433), .A3(new_n434), .A4(G97), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT74), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT74), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n542), .A2(new_n543), .A3(new_n544), .A4(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n540), .A2(new_n303), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n259), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n550));
  OAI211_X1 g0350(.A(G244), .B(new_n256), .C1(new_n260), .C2(new_n261), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT4), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g0353(.A1(KEYINPUT4), .A2(G244), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n256), .B(new_n554), .C1(new_n260), .C2(new_n261), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT75), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n265), .A2(KEYINPUT75), .A3(new_n256), .A4(new_n554), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n550), .A2(new_n553), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT76), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n279), .A2(G45), .A3(new_n280), .ZN(new_n561));
  AND2_X1   g0361(.A1(KEYINPUT5), .A2(G41), .ZN(new_n562));
  NOR2_X1   g0362(.A1(KEYINPUT5), .A2(G41), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(G257), .B(new_n270), .C1(new_n561), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n476), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n559), .A2(new_n271), .B1(new_n560), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(KEYINPUT76), .A3(new_n476), .ZN(new_n568));
  AOI21_X1  g0368(.A(G200), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G283), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n265), .A2(G250), .A3(G1698), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n553), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n557), .A2(new_n558), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n271), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n566), .A2(new_n560), .ZN(new_n575));
  AND4_X1   g0375(.A1(new_n401), .A2(new_n574), .A3(new_n568), .A4(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n549), .B1(new_n569), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n568), .A3(new_n575), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n321), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n546), .A2(new_n548), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n303), .B1(new_n538), .B2(new_n539), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n574), .A2(new_n575), .A3(new_n319), .A4(new_n568), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n232), .A2(new_n256), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n412), .A2(G1698), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n586), .B(new_n587), .C1(new_n260), .C2(new_n261), .ZN(new_n588));
  OAI21_X1  g0388(.A(G33), .B1(new_n496), .B2(new_n497), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT78), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n588), .A2(new_n589), .A3(KEYINPUT78), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n271), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n561), .A2(G250), .A3(new_n270), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n274), .A2(G45), .A3(new_n310), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G200), .ZN(new_n600));
  INV_X1    g0400(.A(new_n407), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(new_n304), .ZN(new_n602));
  AND4_X1   g0402(.A1(G87), .A2(new_n304), .A3(new_n434), .A4(new_n433), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT19), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n299), .B2(new_n534), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n265), .A2(new_n214), .A3(G68), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n214), .B1(new_n385), .B2(new_n604), .ZN(new_n607));
  NOR2_X1   g0407(.A1(G97), .A2(G107), .ZN(new_n608));
  INV_X1    g0408(.A(G87), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n605), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  AOI211_X1 g0412(.A(new_n602), .B(new_n603), .C1(new_n612), .C2(new_n303), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n270), .B1(new_n590), .B2(new_n591), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n597), .B1(new_n614), .B2(new_n593), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G190), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n600), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n612), .A2(new_n303), .ZN(new_n618));
  INV_X1    g0418(.A(new_n602), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n307), .A2(new_n601), .A3(new_n433), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n594), .A2(new_n319), .A3(new_n598), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n621), .B(new_n622), .C1(G169), .C2(new_n615), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n585), .A2(new_n624), .ZN(new_n625));
  AND4_X1   g0425(.A1(new_n426), .A2(new_n488), .A3(new_n531), .A4(new_n625), .ZN(G372));
  INV_X1    g0426(.A(new_n323), .ZN(new_n627));
  INV_X1    g0427(.A(new_n403), .ZN(new_n628));
  INV_X1    g0428(.A(new_n424), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n398), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n357), .A2(new_n362), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n353), .B(new_n359), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n627), .B1(new_n632), .B2(new_n318), .ZN(new_n633));
  INV_X1    g0433(.A(new_n426), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n602), .B1(new_n612), .B2(new_n303), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n615), .A2(new_n319), .B1(new_n635), .B2(new_n620), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT85), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n637), .B1(new_n599), .B2(new_n321), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n615), .A2(KEYINPUT85), .A3(G169), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n574), .A2(new_n568), .A3(new_n575), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n642), .A2(new_n319), .B1(new_n581), .B2(new_n580), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n643), .A2(new_n623), .A3(new_n617), .A4(new_n579), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n641), .B1(new_n644), .B2(KEYINPUT26), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n599), .A2(new_n637), .A3(new_n321), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT85), .B1(new_n615), .B2(G169), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n399), .B1(new_n594), .B2(new_n598), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(G190), .B2(new_n615), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n636), .A2(new_n648), .B1(new_n650), .B2(new_n613), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n645), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n651), .A2(new_n487), .A3(new_n584), .A4(new_n577), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT87), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT86), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n481), .B(new_n658), .C1(new_n438), .C2(new_n456), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n479), .A2(new_n319), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(G169), .B2(new_n479), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n460), .A2(new_n461), .B1(new_n464), .B2(new_n455), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT86), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n530), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n656), .B1(new_n657), .B2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n530), .A2(new_n659), .A3(new_n663), .A4(KEYINPUT87), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n655), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n633), .B1(new_n634), .B2(new_n667), .ZN(G369));
  NOR2_X1   g0468(.A1(new_n207), .A2(G20), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n310), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n505), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n531), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n530), .B2(new_n676), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G330), .ZN(new_n679));
  INV_X1    g0479(.A(new_n675), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n482), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n457), .A2(new_n466), .A3(new_n675), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n482), .A2(new_n682), .A3(new_n487), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n683), .A2(KEYINPUT88), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(KEYINPUT88), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n681), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n679), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n530), .A2(new_n675), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n684), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n663), .A2(new_n659), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n680), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n687), .A2(new_n692), .ZN(G399));
  NOR2_X1   g0493(.A1(new_n210), .A2(G41), .ZN(new_n694));
  NOR4_X1   g0494(.A1(new_n694), .A2(new_n275), .A3(G116), .A4(new_n610), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n695), .B1(new_n220), .B2(new_n694), .ZN(new_n696));
  XOR2_X1   g0496(.A(new_n696), .B(KEYINPUT28), .Z(new_n697));
  INV_X1    g0497(.A(KEYINPUT91), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n487), .A2(new_n640), .A3(new_n617), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n585), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n482), .A2(new_n530), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n641), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n652), .B1(new_n624), .B2(new_n584), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT90), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n653), .A2(KEYINPUT26), .A3(new_n640), .A4(new_n617), .ZN(new_n706));
  OAI211_X1 g0506(.A(KEYINPUT90), .B(new_n652), .C1(new_n624), .C2(new_n584), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n702), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n698), .B1(new_n709), .B2(new_n680), .ZN(new_n710));
  AOI211_X1 g0510(.A(KEYINPUT91), .B(new_n675), .C1(new_n702), .C2(new_n708), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT29), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n664), .A2(new_n657), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n666), .A3(new_n700), .ZN(new_n714));
  INV_X1    g0514(.A(new_n655), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n680), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT29), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT89), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n474), .A2(new_n478), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n520), .A2(new_n723), .A3(new_n521), .A4(new_n615), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n724), .B2(new_n578), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n521), .A2(new_n723), .A3(new_n615), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n726), .A2(KEYINPUT30), .A3(new_n520), .A4(new_n642), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n615), .A2(G179), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n517), .A2(new_n728), .A3(new_n479), .A4(new_n578), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n725), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT31), .B1(new_n730), .B2(new_n675), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n721), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n730), .A2(new_n675), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(KEYINPUT89), .A3(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n531), .A2(new_n488), .A3(new_n625), .A4(new_n680), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n733), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n720), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n697), .B1(new_n743), .B2(G1), .ZN(G364));
  NOR2_X1   g0544(.A1(new_n678), .A2(G330), .ZN(new_n745));
  INV_X1    g0545(.A(new_n679), .ZN(new_n746));
  INV_X1    g0546(.A(new_n694), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n275), .B1(new_n669), .B2(G45), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n745), .B(new_n746), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n213), .B1(G20), .B2(new_n321), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n214), .A2(new_n319), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(G190), .A3(G200), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT93), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n468), .A2(new_n469), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n319), .A2(new_n399), .A3(G190), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n754), .A2(G326), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT94), .ZN(new_n760));
  NOR4_X1   g0560(.A1(new_n214), .A2(new_n319), .A3(new_n401), .A4(G200), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n265), .B1(new_n761), .B2(G322), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G190), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n752), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n214), .A2(G179), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n763), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G311), .A2(new_n765), .B1(new_n768), .B2(G329), .ZN(new_n769));
  INV_X1    g0569(.A(G283), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n766), .A2(new_n401), .A3(G200), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n766), .A2(G190), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(G303), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n770), .A2(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR4_X1   g0574(.A1(new_n214), .A2(new_n319), .A3(new_n399), .A4(G190), .ZN(new_n775));
  INV_X1    g0575(.A(G317), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n776), .A2(KEYINPUT33), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(KEYINPUT33), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n774), .B1(new_n775), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n760), .A2(new_n762), .A3(new_n769), .A4(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n761), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n265), .B1(new_n782), .B2(new_n216), .ZN(new_n783));
  INV_X1    g0583(.A(new_n775), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n784), .A2(new_n217), .B1(new_n771), .B2(new_n415), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n783), .B(new_n785), .C1(G97), .C2(new_n758), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n772), .A2(new_n609), .ZN(new_n787));
  INV_X1    g0587(.A(G159), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n767), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT32), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n790), .B1(new_n225), .B2(new_n753), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n787), .B(new_n791), .C1(new_n790), .C2(new_n789), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n764), .A2(KEYINPUT92), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n764), .A2(KEYINPUT92), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n786), .B(new_n792), .C1(new_n372), .C2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n751), .B1(new_n781), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n748), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n694), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(G355), .A2(new_n209), .A3(new_n265), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(G116), .B2(new_n209), .ZN(new_n801));
  INV_X1    g0601(.A(G45), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n251), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n209), .A2(new_n262), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(new_n802), .B2(new_n220), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n801), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(G13), .A2(G33), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(G20), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n750), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n799), .B1(new_n806), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n797), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n809), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n678), .B2(new_n814), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT95), .Z(new_n816));
  NOR2_X1   g0616(.A1(new_n749), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G396));
  INV_X1    g0618(.A(new_n799), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n750), .A2(new_n807), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT96), .Z(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n819), .B1(new_n822), .B2(new_n372), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n753), .A2(new_n773), .B1(new_n772), .B2(new_n415), .ZN(new_n824));
  INV_X1    g0624(.A(G311), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n262), .B1(new_n767), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G294), .B2(new_n761), .ZN(new_n827));
  INV_X1    g0627(.A(new_n771), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n828), .A2(G87), .B1(new_n758), .B2(G97), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n827), .B(new_n829), .C1(new_n795), .C2(new_n498), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n824), .B(new_n830), .C1(G283), .C2(new_n775), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n265), .B1(new_n767), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT98), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n771), .A2(new_n217), .ZN(new_n835));
  INV_X1    g0635(.A(new_n758), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n836), .A2(new_n216), .B1(new_n772), .B2(new_n225), .ZN(new_n837));
  OR3_X1    g0637(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n753), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n839), .A2(G137), .B1(new_n761), .B2(G143), .ZN(new_n840));
  INV_X1    g0640(.A(G150), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n840), .B1(new_n841), .B2(new_n784), .C1(new_n795), .C2(new_n788), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  XOR2_X1   g0643(.A(KEYINPUT97), .B(KEYINPUT34), .Z(new_n844));
  AOI21_X1  g0644(.A(new_n838), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n831), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n424), .A2(new_n675), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n411), .A2(new_n675), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT99), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n411), .A2(KEYINPUT99), .A3(new_n675), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n421), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n848), .B1(new_n853), .B2(new_n424), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n823), .B1(new_n847), .B2(new_n751), .C1(new_n854), .C2(new_n808), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n853), .A2(new_n424), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n717), .B1(new_n848), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n854), .A2(new_n680), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n858), .B1(new_n667), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n741), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n819), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n860), .A2(new_n741), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n855), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT100), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(G384));
  NOR2_X1   g0666(.A1(new_n310), .A2(new_n669), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT39), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n217), .B1(new_n339), .B2(new_n340), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n333), .B1(new_n337), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(new_n346), .A3(new_n303), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n350), .ZN(new_n872));
  INV_X1    g0672(.A(new_n673), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n363), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n351), .A2(new_n873), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n352), .A2(new_n877), .A3(new_n878), .A4(new_n360), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n332), .A2(new_n872), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n880), .A2(new_n874), .A3(new_n360), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n879), .B1(new_n881), .B2(new_n878), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n876), .A2(new_n882), .A3(KEYINPUT38), .ZN(new_n883));
  INV_X1    g0683(.A(new_n877), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n363), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n352), .A2(new_n877), .A3(new_n360), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT37), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n879), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT38), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n868), .B1(new_n883), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n876), .A2(new_n882), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n876), .A2(new_n882), .A3(KEYINPUT38), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(KEYINPUT39), .A3(new_n894), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n398), .A2(new_n680), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n848), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n667), .B2(new_n859), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n893), .A2(new_n894), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n396), .A2(new_n397), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n378), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n379), .A2(KEYINPUT101), .A3(new_n680), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT101), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n378), .B2(new_n675), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n904), .A2(new_n628), .A3(new_n908), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n398), .A2(new_n403), .B1(new_n907), .B2(new_n905), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n901), .A2(new_n902), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n353), .A2(new_n359), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n673), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n899), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n712), .A2(new_n426), .A3(new_n719), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n633), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n916), .B(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(G330), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n909), .A2(new_n854), .A3(new_n910), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n731), .A2(new_n732), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n921), .B1(new_n922), .B2(new_n739), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n363), .A2(new_n884), .B1(new_n887), .B2(new_n879), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n894), .B1(KEYINPUT38), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT40), .B1(new_n893), .B2(new_n894), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n926), .A2(KEYINPUT40), .B1(new_n927), .B2(new_n923), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n634), .B1(new_n922), .B2(new_n739), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n920), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n930), .B2(new_n929), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n867), .B1(new_n919), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n919), .B2(new_n932), .ZN(new_n934));
  INV_X1    g0734(.A(new_n537), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(KEYINPUT35), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(KEYINPUT35), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n936), .A2(G116), .A3(new_n215), .A4(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT36), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n220), .B(G77), .C1(new_n216), .C2(new_n233), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(G50), .B2(new_n217), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(new_n207), .A3(new_n281), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n934), .A2(new_n939), .A3(new_n942), .ZN(G367));
  NOR2_X1   g0743(.A1(new_n246), .A2(new_n804), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n810), .B1(new_n209), .B2(new_n407), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n799), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(KEYINPUT46), .A2(G116), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n534), .A2(new_n771), .B1(new_n772), .B2(new_n947), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n784), .A2(new_n755), .B1(new_n415), .B2(new_n836), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n948), .B(new_n949), .C1(new_n754), .C2(G311), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n262), .B1(new_n767), .B2(new_n776), .C1(new_n782), .C2(new_n773), .ZN(new_n951));
  INV_X1    g0751(.A(new_n795), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n951), .B1(new_n952), .B2(G283), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n772), .A2(new_n498), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n950), .B(new_n953), .C1(KEYINPUT46), .C2(new_n954), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n836), .A2(new_n217), .B1(new_n772), .B2(new_n216), .ZN(new_n956));
  INV_X1    g0756(.A(G137), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n265), .B1(new_n767), .B2(new_n957), .C1(new_n782), .C2(new_n841), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n956), .B(new_n958), .C1(G77), .C2(new_n828), .ZN(new_n959));
  INV_X1    g0759(.A(G143), .ZN(new_n960));
  INV_X1    g0760(.A(new_n754), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n795), .A2(new_n225), .B1(new_n788), .B2(new_n784), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT103), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n955), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT47), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n946), .B1(new_n966), .B2(new_n750), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n640), .A2(new_n613), .A3(new_n680), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n680), .A2(new_n613), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n968), .B1(new_n651), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n809), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n686), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n689), .B1(new_n973), .B2(new_n688), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(new_n746), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT45), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n577), .B(new_n584), .C1(new_n549), .C2(new_n680), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n653), .A2(new_n675), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n976), .B1(new_n692), .B2(new_n980), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n689), .A2(KEYINPUT45), .A3(new_n691), .A4(new_n979), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT102), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n981), .A2(new_n982), .B1(new_n687), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n979), .B1(new_n689), .B2(new_n691), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT44), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n687), .A2(new_n983), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n984), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n988), .B1(new_n984), .B2(new_n986), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n743), .B(new_n975), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n743), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n694), .B(KEYINPUT41), .Z(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n798), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT43), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n970), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n689), .A2(new_n980), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n999), .A2(KEYINPUT42), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n584), .B1(new_n977), .B2(new_n482), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n999), .A2(KEYINPUT42), .B1(new_n680), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n998), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n970), .A2(new_n997), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1000), .A2(new_n1002), .A3(new_n997), .A4(new_n970), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n687), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(new_n980), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1006), .A2(new_n1010), .A3(new_n1007), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n972), .B1(new_n996), .B2(new_n1014), .ZN(G387));
  OR3_X1    g0815(.A1(new_n243), .A2(new_n802), .A3(new_n265), .ZN(new_n1016));
  OAI21_X1  g0816(.A(KEYINPUT50), .B1(new_n300), .B2(G50), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1017), .B(new_n802), .C1(new_n217), .C2(new_n372), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n300), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n262), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(G116), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1020), .A2(new_n609), .A3(new_n1021), .A4(new_n608), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n210), .B1(new_n1016), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n810), .B1(new_n415), .B2(new_n209), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G311), .A2(new_n775), .B1(new_n761), .B2(G317), .ZN(new_n1025));
  XOR2_X1   g0825(.A(KEYINPUT105), .B(G322), .Z(new_n1026));
  OAI221_X1 g0826(.A(new_n1025), .B1(new_n795), .B2(new_n773), .C1(new_n961), .C2(new_n1026), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1027), .A2(KEYINPUT106), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(KEYINPUT106), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(KEYINPUT48), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT48), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1028), .A2(new_n1032), .A3(new_n1029), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n772), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n756), .A2(new_n1034), .B1(G283), .B2(new_n758), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT49), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n265), .B1(new_n768), .B2(G326), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n498), .B2(new_n771), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n836), .A2(new_n407), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G50), .B2(new_n761), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT104), .Z(new_n1045));
  OAI22_X1  g0845(.A1(new_n784), .A2(new_n300), .B1(new_n771), .B2(new_n534), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n265), .B1(new_n767), .B2(new_n841), .C1(new_n217), .C2(new_n764), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n772), .A2(new_n372), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n753), .A2(new_n788), .ZN(new_n1049));
  NOR4_X1   g0849(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1041), .A2(new_n1042), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n799), .B1(new_n1023), .B2(new_n1024), .C1(new_n1051), .C2(new_n751), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT107), .Z(new_n1053));
  NAND2_X1  g0853(.A1(new_n686), .A2(new_n809), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1053), .A2(new_n1054), .B1(new_n798), .B2(new_n975), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n743), .A2(new_n975), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n743), .A2(new_n975), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n694), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1055), .B1(new_n1056), .B2(new_n1058), .ZN(G393));
  INV_X1    g0859(.A(new_n991), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1060), .A2(new_n1057), .A3(new_n989), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n992), .A2(new_n1061), .A3(new_n694), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n989), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n980), .A2(new_n809), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n254), .A2(new_n804), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n810), .B1(new_n534), .B2(new_n209), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n799), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n265), .B1(new_n767), .B2(new_n960), .C1(new_n609), .C2(new_n771), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n952), .B2(new_n405), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n836), .A2(new_n372), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G50), .B2(new_n775), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1069), .B(new_n1071), .C1(new_n233), .C2(new_n772), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n839), .A2(G150), .B1(new_n761), .B2(G159), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT51), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1076), .A2(KEYINPUT108), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n262), .B1(new_n764), .B2(new_n467), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n784), .A2(new_n773), .B1(new_n498), .B2(new_n836), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(G107), .C2(new_n828), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n782), .A2(new_n825), .B1(new_n776), .B2(new_n753), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT52), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n767), .A2(new_n1026), .B1(new_n772), .B2(new_n770), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1084), .A2(KEYINPUT109), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(KEYINPUT109), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1080), .A2(new_n1082), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1076), .A2(KEYINPUT108), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1077), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1067), .B1(new_n1089), .B2(new_n750), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1063), .A2(new_n798), .B1(new_n1064), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1062), .A2(new_n1091), .ZN(G390));
  AOI21_X1  g0892(.A(new_n920), .B1(new_n922), .B2(new_n739), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n912), .B1(new_n1093), .B2(new_n854), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n482), .A2(new_n530), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n640), .B1(new_n1095), .B2(new_n656), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n707), .A2(new_n706), .ZN(new_n1097));
  AOI21_X1  g0897(.A(KEYINPUT90), .B1(new_n644), .B2(new_n652), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n680), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(KEYINPUT91), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n709), .A2(new_n698), .A3(new_n680), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1101), .A2(new_n1102), .A3(new_n900), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1094), .B1(new_n856), .B2(new_n1103), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n740), .A2(G330), .A3(new_n854), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n912), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n740), .A2(G330), .A3(new_n854), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT111), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(new_n1109), .A3(new_n911), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1109), .B1(new_n1108), .B2(new_n911), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1093), .A2(new_n854), .A3(new_n912), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1111), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n859), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n848), .B1(new_n716), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1107), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n426), .A2(new_n1093), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n917), .A2(new_n633), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1103), .A2(new_n856), .A3(new_n912), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n897), .B(KEYINPUT110), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n925), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n890), .A2(new_n895), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n897), .B1(new_n1117), .B2(new_n911), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1123), .A2(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n710), .A2(new_n711), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n857), .B1(new_n1130), .B2(new_n900), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1125), .B1(new_n1131), .B2(new_n912), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n898), .B1(new_n901), .B2(new_n912), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1106), .B1(new_n1133), .B2(new_n896), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n1129), .A2(new_n1113), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1122), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1108), .A2(new_n911), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(KEYINPUT111), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n1113), .A3(new_n1110), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1139), .A2(new_n901), .B1(new_n1106), .B2(new_n1104), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1140), .A2(new_n1120), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1135), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1136), .A2(new_n1143), .A3(new_n694), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT112), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n798), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1128), .A2(new_n1127), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1113), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1145), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1128), .A2(new_n1127), .B1(new_n1105), .B2(new_n912), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n748), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1152), .B(KEYINPUT112), .C1(new_n1129), .C2(new_n1113), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n799), .B1(new_n821), .B2(new_n405), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n262), .B1(new_n767), .B2(new_n467), .C1(new_n782), .C2(new_n1021), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1156), .A2(new_n787), .A3(new_n835), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n753), .A2(new_n770), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1158), .B(new_n1070), .C1(G107), .C2(new_n775), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1157), .B(new_n1159), .C1(new_n534), .C2(new_n795), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT113), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n782), .A2(new_n832), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n262), .B(new_n1163), .C1(G125), .C2(new_n768), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n784), .A2(new_n957), .B1(new_n788), .B2(new_n836), .ZN(new_n1165));
  INV_X1    g0965(.A(G128), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n753), .A2(new_n1166), .B1(new_n771), .B2(new_n225), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT54), .B(G143), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n952), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n772), .A2(new_n841), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT53), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1164), .A2(new_n1168), .A3(new_n1171), .A4(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1162), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1155), .B1(new_n1176), .B2(new_n750), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n896), .B2(new_n808), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT114), .B1(new_n1154), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT114), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1178), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(new_n1150), .C2(new_n1153), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1144), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT115), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT115), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1185), .B(new_n1144), .C1(new_n1179), .C2(new_n1182), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1184), .A2(new_n1186), .ZN(G378));
  AOI21_X1  g0987(.A(new_n819), .B1(new_n225), .B2(new_n820), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT118), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n265), .A2(G41), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G283), .B2(new_n768), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n415), .B2(new_n782), .C1(new_n407), .C2(new_n764), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1048), .B(new_n1192), .C1(G68), .C2(new_n758), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n771), .A2(new_n216), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G116), .B2(new_n839), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1193), .B(new_n1195), .C1(new_n534), .C2(new_n784), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT58), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(G33), .A2(G41), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1198), .A2(G50), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1196), .A2(new_n1197), .B1(new_n1190), .B2(new_n1199), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT116), .Z(new_n1201));
  INV_X1    g1001(.A(G124), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1198), .B1(new_n767), .B2(new_n1202), .C1(new_n788), .C2(new_n771), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n782), .A2(new_n1166), .B1(new_n764), .B2(new_n957), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G125), .B2(new_n839), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1034), .A2(new_n1170), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT117), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n775), .A2(G132), .B1(new_n758), .B2(G150), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1205), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1203), .B1(new_n1209), .B2(KEYINPUT59), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(KEYINPUT59), .B2(new_n1209), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1201), .B(new_n1211), .C1(new_n1197), .C2(new_n1196), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1189), .B1(new_n1212), .B2(new_n750), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n313), .A2(new_n873), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n318), .A2(new_n323), .A3(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1216), .B1(new_n318), .B2(new_n323), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1215), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1219), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1221), .A2(new_n1217), .A3(new_n1214), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1213), .B1(new_n1223), .B2(new_n808), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT119), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n916), .B2(KEYINPUT120), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1223), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n928), .B2(new_n920), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n927), .A2(new_n923), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT40), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n923), .B2(new_n925), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G330), .B(new_n1223), .C1(new_n1230), .C2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1228), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1226), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1228), .A2(new_n1225), .A3(new_n1233), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT120), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n916), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1235), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1224), .B1(new_n1240), .B2(new_n748), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT57), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1120), .B(KEYINPUT121), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1242), .B1(new_n1240), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1243), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1122), .B2(new_n1135), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1234), .A2(new_n916), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1239), .A2(new_n1228), .A3(new_n1233), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1242), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n747), .B1(new_n1247), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1241), .B1(new_n1245), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(G375));
  OAI211_X1 g1053(.A(new_n1107), .B(new_n1120), .C1(new_n1115), .C2(new_n1117), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1122), .A2(new_n995), .A3(new_n1254), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(G150), .A2(new_n765), .B1(new_n761), .B2(G137), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1256), .B(new_n265), .C1(new_n1166), .C2(new_n767), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1194), .B(new_n1257), .C1(new_n775), .C2(new_n1170), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n836), .A2(new_n225), .B1(new_n772), .B2(new_n788), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(G132), .B2(new_n839), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n262), .B1(new_n767), .B2(new_n773), .C1(new_n372), .C2(new_n771), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n839), .A2(G294), .B1(new_n775), .B2(new_n492), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n534), .B2(new_n772), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1261), .B(new_n1263), .C1(G107), .C2(new_n952), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1043), .B1(G283), .B2(new_n761), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(KEYINPUT122), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1258), .A2(new_n1260), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n799), .B1(G68), .B2(new_n821), .C1(new_n1267), .C2(new_n751), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(new_n911), .B2(new_n807), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n1118), .B2(new_n798), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1255), .A2(new_n1270), .ZN(G381));
  INV_X1    g1071(.A(new_n1183), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1252), .A2(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1055), .B(new_n817), .C1(new_n1056), .C2(new_n1058), .ZN(new_n1274));
  OR4_X1    g1074(.A1(G384), .A2(G381), .A3(new_n1274), .A4(G390), .ZN(new_n1275));
  OR3_X1    g1075(.A1(new_n1273), .A2(new_n1275), .A3(G387), .ZN(G407));
  OAI211_X1 g1076(.A(G407), .B(G213), .C1(G343), .C2(new_n1273), .ZN(G409));
  NAND3_X1  g1077(.A1(new_n1184), .A2(new_n1186), .A3(new_n1252), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1240), .A2(new_n1244), .A3(new_n994), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1224), .B1(new_n1280), .B2(new_n748), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1272), .B1(new_n1279), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n674), .A2(G213), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1140), .A2(KEYINPUT124), .A3(KEYINPUT60), .A4(new_n1120), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1286), .A2(new_n694), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT60), .B1(new_n1140), .B2(new_n1120), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT123), .B1(new_n1288), .B2(new_n1141), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT124), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT60), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1290), .B1(new_n1254), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1254), .A2(new_n1291), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT123), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n1294), .A3(new_n1122), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1287), .A2(new_n1289), .A3(new_n1292), .A4(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1296), .A2(G384), .A3(new_n1270), .ZN(new_n1297));
  AOI21_X1  g1097(.A(G384), .B1(new_n1296), .B2(new_n1270), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1284), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(G2897), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1297), .A2(new_n1298), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1289), .A2(new_n1295), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1292), .A2(new_n694), .A3(new_n1286), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1270), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n865), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1296), .A2(G384), .A3(new_n1270), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1300), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1302), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT61), .B1(new_n1285), .B2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1299), .B1(new_n1278), .B2(new_n1282), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1311), .A2(KEYINPUT62), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT62), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1310), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n972), .B(G390), .C1(new_n996), .C2(new_n1014), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT125), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(G393), .A2(G396), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1274), .ZN(new_n1320));
  INV_X1    g1120(.A(G390), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1057), .B1(new_n1060), .B2(new_n989), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n995), .B1(new_n1322), .B2(new_n742), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1014), .B1(new_n1323), .B2(new_n748), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n972), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1321), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  AOI22_X1  g1126(.A1(new_n1318), .A2(new_n1320), .B1(new_n1316), .B2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1326), .A2(new_n1316), .A3(KEYINPUT125), .A4(new_n1320), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  XNOR2_X1  g1130(.A(new_n1330), .B(KEYINPUT127), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1315), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT126), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT63), .ZN(new_n1334));
  NOR3_X1   g1134(.A1(new_n1297), .A2(new_n1298), .A3(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1283), .A2(new_n1284), .A3(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1330), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT61), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1301), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1306), .A2(new_n1307), .A3(new_n1300), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1338), .B1(new_n1311), .B2(new_n1341), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1337), .A2(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1283), .A2(new_n1284), .A3(new_n1312), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(new_n1334), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1333), .B1(new_n1343), .B2(new_n1345), .ZN(new_n1346));
  AOI22_X1  g1146(.A1(new_n1311), .A2(new_n1335), .B1(new_n1329), .B2(new_n1328), .ZN(new_n1347));
  AND4_X1   g1147(.A1(new_n1333), .A2(new_n1310), .A3(new_n1347), .A4(new_n1345), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1332), .B1(new_n1346), .B2(new_n1348), .ZN(G405));
  NAND2_X1  g1149(.A1(G375), .A2(new_n1272), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(new_n1278), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1312), .ZN(new_n1352));
  XNOR2_X1  g1152(.A(new_n1351), .B(new_n1352), .ZN(new_n1353));
  XNOR2_X1  g1153(.A(new_n1353), .B(new_n1330), .ZN(G402));
endmodule


