

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743;

  NOR2_X1 U369 ( .A1(n538), .A2(n537), .ZN(n599) );
  INV_X1 U370 ( .A(G953), .ZN(n406) );
  AND2_X2 U371 ( .A1(n741), .A2(KEYINPUT44), .ZN(n530) );
  XNOR2_X2 U372 ( .A(n425), .B(KEYINPUT35), .ZN(n741) );
  NOR2_X2 U373 ( .A1(n553), .A2(n552), .ZN(n681) );
  NOR2_X1 U374 ( .A1(n630), .A2(n631), .ZN(n362) );
  XNOR2_X1 U375 ( .A(n503), .B(n502), .ZN(n653) );
  INV_X2 U376 ( .A(n482), .ZN(n483) );
  NOR2_X1 U377 ( .A1(n374), .A2(n715), .ZN(n708) );
  NAND2_X1 U378 ( .A1(n411), .A2(n352), .ZN(n619) );
  XNOR2_X1 U379 ( .A(n412), .B(n606), .ZN(n411) );
  NOR2_X1 U380 ( .A1(n609), .A2(n612), .ZN(n386) );
  XNOR2_X1 U381 ( .A(n423), .B(KEYINPUT19), .ZN(n592) );
  NOR2_X1 U382 ( .A1(n688), .A2(n602), .ZN(n603) );
  NOR2_X1 U383 ( .A1(n643), .A2(n644), .ZN(n542) );
  XNOR2_X1 U384 ( .A(n375), .B(KEYINPUT108), .ZN(n602) );
  OR2_X1 U385 ( .A1(n601), .A2(n600), .ZN(n375) );
  XNOR2_X1 U386 ( .A(n653), .B(KEYINPUT6), .ZN(n601) );
  XNOR2_X1 U387 ( .A(n481), .B(n424), .ZN(n716) );
  NAND2_X1 U388 ( .A1(n399), .A2(n485), .ZN(n504) );
  INV_X1 U389 ( .A(KEYINPUT36), .ZN(n385) );
  XNOR2_X1 U390 ( .A(G110), .B(KEYINPUT70), .ZN(n441) );
  NOR2_X2 U391 ( .A1(n681), .A2(n742), .ZN(n559) );
  XNOR2_X1 U392 ( .A(n453), .B(n452), .ZN(n717) );
  INV_X1 U393 ( .A(n618), .ZN(n721) );
  NOR2_X1 U394 ( .A1(n633), .A2(n634), .ZN(n638) );
  INV_X1 U395 ( .A(KEYINPUT0), .ZN(n378) );
  NAND2_X1 U396 ( .A1(n592), .A2(n463), .ZN(n379) );
  BUF_X1 U397 ( .A(n653), .Z(n416) );
  NAND2_X2 U398 ( .A1(n415), .A2(n617), .ZN(n356) );
  NAND2_X1 U399 ( .A1(n721), .A2(n395), .ZN(n394) );
  NOR2_X1 U400 ( .A1(n619), .A2(n396), .ZN(n395) );
  INV_X1 U401 ( .A(KEYINPUT2), .ZN(n396) );
  INV_X1 U402 ( .A(KEYINPUT44), .ZN(n381) );
  NOR2_X1 U403 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U404 ( .A1(n401), .A2(n371), .ZN(n412) );
  AND2_X1 U405 ( .A1(n597), .A2(n402), .ZN(n371) );
  XNOR2_X1 U406 ( .A(G902), .B(KEYINPUT15), .ZN(n464) );
  INV_X1 U407 ( .A(G134), .ZN(n484) );
  XNOR2_X1 U408 ( .A(n716), .B(n446), .ZN(n447) );
  XOR2_X1 U409 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n445) );
  XNOR2_X1 U410 ( .A(G146), .B(G125), .ZN(n469) );
  XNOR2_X1 U411 ( .A(n480), .B(n479), .ZN(n647) );
  XNOR2_X1 U412 ( .A(n478), .B(n429), .ZN(n479) );
  NOR2_X1 U413 ( .A1(n713), .A2(G902), .ZN(n480) );
  XOR2_X1 U414 ( .A(G122), .B(G104), .Z(n517) );
  XNOR2_X1 U415 ( .A(G143), .B(G140), .ZN(n516) );
  XNOR2_X1 U416 ( .A(n524), .B(n373), .ZN(n372) );
  INV_X1 U417 ( .A(KEYINPUT98), .ZN(n373) );
  XNOR2_X1 U418 ( .A(G113), .B(G131), .ZN(n524) );
  XNOR2_X1 U419 ( .A(n382), .B(n491), .ZN(n620) );
  XNOR2_X1 U420 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U421 ( .A(n495), .B(n481), .ZN(n382) );
  NOR2_X1 U422 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U423 ( .A1(n534), .A2(n542), .ZN(n398) );
  XNOR2_X1 U424 ( .A(n376), .B(KEYINPUT41), .ZN(n665) );
  XNOR2_X1 U425 ( .A(n579), .B(KEYINPUT39), .ZN(n608) );
  INV_X1 U426 ( .A(n633), .ZN(n585) );
  BUF_X1 U427 ( .A(n644), .Z(n370) );
  INV_X1 U428 ( .A(KEYINPUT34), .ZN(n428) );
  XNOR2_X1 U429 ( .A(n533), .B(KEYINPUT22), .ZN(n556) );
  INV_X1 U430 ( .A(n370), .ZN(n610) );
  AND2_X1 U431 ( .A1(n417), .A2(n416), .ZN(n582) );
  INV_X1 U432 ( .A(n600), .ZN(n417) );
  NAND2_X2 U433 ( .A1(n390), .A2(n387), .ZN(n584) );
  OR2_X1 U434 ( .A1(n620), .A2(n388), .ZN(n387) );
  AND2_X1 U435 ( .A1(n392), .A2(n391), .ZN(n390) );
  NAND2_X1 U436 ( .A1(G469), .A2(n389), .ZN(n388) );
  INV_X1 U437 ( .A(n416), .ZN(n418) );
  AND2_X1 U438 ( .A1(n394), .A2(G472), .ZN(n363) );
  AND2_X1 U439 ( .A1(n394), .A2(G469), .ZN(n364) );
  AND2_X1 U440 ( .A1(n365), .A2(n356), .ZN(n704) );
  AND2_X1 U441 ( .A1(n394), .A2(G210), .ZN(n365) );
  XNOR2_X1 U442 ( .A(n404), .B(n403), .ZN(n402) );
  INV_X1 U443 ( .A(KEYINPUT81), .ZN(n403) );
  INV_X1 U444 ( .A(KEYINPUT47), .ZN(n367) );
  INV_X1 U445 ( .A(KEYINPUT48), .ZN(n606) );
  INV_X1 U446 ( .A(KEYINPUT45), .ZN(n563) );
  OR2_X1 U447 ( .A1(G237), .A2(G902), .ZN(n457) );
  XOR2_X1 U448 ( .A(KEYINPUT92), .B(KEYINPUT20), .Z(n466) );
  NOR2_X1 U449 ( .A1(G953), .A2(G237), .ZN(n520) );
  XOR2_X1 U450 ( .A(KEYINPUT85), .B(KEYINPUT74), .Z(n434) );
  NAND2_X1 U451 ( .A1(G234), .A2(G237), .ZN(n461) );
  XNOR2_X1 U452 ( .A(n598), .B(n578), .ZN(n633) );
  XNOR2_X1 U453 ( .A(n584), .B(KEYINPUT1), .ZN(n644) );
  NOR2_X1 U454 ( .A1(n408), .A2(n580), .ZN(n407) );
  AND2_X1 U455 ( .A1(n653), .A2(n604), .ZN(n565) );
  INV_X1 U456 ( .A(G902), .ZN(n389) );
  NAND2_X1 U457 ( .A1(n393), .A2(G902), .ZN(n391) );
  XOR2_X1 U458 ( .A(KEYINPUT5), .B(G137), .Z(n497) );
  INV_X1 U459 ( .A(G146), .ZN(n357) );
  XNOR2_X1 U460 ( .A(KEYINPUT69), .B(KEYINPUT96), .ZN(n492) );
  XOR2_X1 U461 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n493) );
  XNOR2_X1 U462 ( .A(n717), .B(n489), .ZN(n499) );
  XNOR2_X1 U463 ( .A(G113), .B(KEYINPUT3), .ZN(n449) );
  XNOR2_X1 U464 ( .A(KEYINPUT16), .B(G122), .ZN(n424) );
  XNOR2_X1 U465 ( .A(KEYINPUT65), .B(KEYINPUT8), .ZN(n472) );
  XNOR2_X1 U466 ( .A(G116), .B(G107), .ZN(n505) );
  XOR2_X1 U467 ( .A(KEYINPUT7), .B(G122), .Z(n506) );
  NAND2_X1 U468 ( .A1(n598), .A2(n604), .ZN(n423) );
  XNOR2_X1 U469 ( .A(n523), .B(n372), .ZN(n525) );
  INV_X1 U470 ( .A(KEYINPUT78), .ZN(n361) );
  INV_X1 U471 ( .A(n394), .ZN(n631) );
  AND2_X1 U472 ( .A1(n669), .A2(n406), .ZN(n405) );
  XNOR2_X1 U473 ( .A(n586), .B(n587), .ZN(n740) );
  XNOR2_X1 U474 ( .A(n414), .B(n413), .ZN(n743) );
  NAND2_X1 U475 ( .A1(n427), .A2(n426), .ZN(n425) );
  INV_X1 U476 ( .A(n591), .ZN(n426) );
  XNOR2_X1 U477 ( .A(n397), .B(n428), .ZN(n427) );
  XNOR2_X1 U478 ( .A(n558), .B(n368), .ZN(n742) );
  INV_X1 U479 ( .A(KEYINPUT32), .ZN(n368) );
  NOR2_X1 U480 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U481 ( .A1(n418), .A2(n554), .ZN(n553) );
  NAND2_X1 U482 ( .A1(n421), .A2(n420), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n422), .B(n354), .ZN(n421) );
  XNOR2_X1 U484 ( .A(n624), .B(n623), .ZN(n625) );
  INV_X1 U485 ( .A(KEYINPUT56), .ZN(n383) );
  XNOR2_X1 U486 ( .A(n704), .B(n353), .ZN(n377) );
  XOR2_X1 U487 ( .A(KEYINPUT86), .B(n432), .Z(n346) );
  XNOR2_X1 U488 ( .A(KEYINPUT23), .B(KEYINPUT90), .ZN(n347) );
  XOR2_X1 U489 ( .A(KEYINPUT24), .B(G110), .Z(n348) );
  XNOR2_X1 U490 ( .A(G131), .B(KEYINPUT66), .ZN(n349) );
  AND2_X1 U491 ( .A1(n356), .A2(n394), .ZN(n350) );
  INV_X1 U492 ( .A(G469), .ZN(n393) );
  AND2_X1 U493 ( .A1(n647), .A2(n407), .ZN(n351) );
  AND2_X1 U494 ( .A1(n614), .A2(n701), .ZN(n352) );
  XOR2_X1 U495 ( .A(n703), .B(n702), .Z(n353) );
  XNOR2_X1 U496 ( .A(n672), .B(n671), .ZN(n354) );
  XOR2_X1 U497 ( .A(n670), .B(KEYINPUT121), .Z(n355) );
  INV_X1 U498 ( .A(n715), .ZN(n420) );
  NAND2_X1 U499 ( .A1(n364), .A2(n356), .ZN(n624) );
  NAND2_X1 U500 ( .A1(n363), .A2(n356), .ZN(n422) );
  NAND2_X1 U501 ( .A1(n366), .A2(n356), .ZN(n706) );
  XNOR2_X2 U502 ( .A(n358), .B(n357), .ZN(n495) );
  XNOR2_X1 U503 ( .A(n358), .B(KEYINPUT126), .ZN(n730) );
  XNOR2_X2 U504 ( .A(n504), .B(n349), .ZN(n358) );
  XNOR2_X1 U505 ( .A(n359), .B(n355), .ZN(G75) );
  NAND2_X1 U506 ( .A1(n360), .A2(n405), .ZN(n359) );
  XNOR2_X1 U507 ( .A(n362), .B(n361), .ZN(n360) );
  AND2_X1 U508 ( .A1(n394), .A2(G475), .ZN(n366) );
  NAND2_X1 U509 ( .A1(n350), .A2(G217), .ZN(n712) );
  NAND2_X1 U510 ( .A1(n350), .A2(G478), .ZN(n709) );
  XNOR2_X1 U511 ( .A(n706), .B(n707), .ZN(n374) );
  XNOR2_X1 U512 ( .A(n530), .B(n529), .ZN(n549) );
  NAND2_X1 U513 ( .A1(n540), .A2(n532), .ZN(n533) );
  XNOR2_X2 U514 ( .A(n379), .B(n378), .ZN(n540) );
  XNOR2_X1 U515 ( .A(n595), .B(n367), .ZN(n596) );
  NOR2_X2 U516 ( .A1(n556), .A2(n610), .ZN(n551) );
  XNOR2_X2 U517 ( .A(n369), .B(n563), .ZN(n618) );
  NAND2_X1 U518 ( .A1(n562), .A2(n561), .ZN(n369) );
  NOR2_X1 U519 ( .A1(n743), .A2(n740), .ZN(n588) );
  NAND2_X1 U520 ( .A1(n603), .A2(n604), .ZN(n609) );
  INV_X1 U521 ( .A(n646), .ZN(n408) );
  XNOR2_X1 U522 ( .A(n386), .B(n385), .ZN(n605) );
  NAND2_X1 U523 ( .A1(n638), .A2(n635), .ZN(n376) );
  NAND2_X1 U524 ( .A1(n377), .A2(n420), .ZN(n384) );
  NAND2_X1 U525 ( .A1(n380), .A2(n560), .ZN(n561) );
  XNOR2_X1 U526 ( .A(n559), .B(n381), .ZN(n380) );
  XNOR2_X1 U527 ( .A(n384), .B(n383), .ZN(G51) );
  XNOR2_X1 U528 ( .A(n410), .B(KEYINPUT72), .ZN(n574) );
  NOR2_X1 U529 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U530 ( .A1(n409), .A2(n351), .ZN(n410) );
  XNOR2_X1 U531 ( .A(n588), .B(KEYINPUT46), .ZN(n401) );
  XNOR2_X1 U532 ( .A(n476), .B(n731), .ZN(n713) );
  NAND2_X1 U533 ( .A1(n444), .A2(n443), .ZN(n481) );
  XNOR2_X2 U534 ( .A(G128), .B(G143), .ZN(n482) );
  NAND2_X1 U535 ( .A1(n483), .A2(n484), .ZN(n399) );
  NAND2_X1 U536 ( .A1(n620), .A2(n393), .ZN(n392) );
  NAND2_X1 U537 ( .A1(n540), .A2(n664), .ZN(n397) );
  XNOR2_X2 U538 ( .A(n398), .B(KEYINPUT33), .ZN(n664) );
  NOR2_X2 U539 ( .A1(n400), .A2(n618), .ZN(n628) );
  XNOR2_X1 U540 ( .A(n400), .B(n735), .ZN(n734) );
  XNOR2_X2 U541 ( .A(n619), .B(KEYINPUT80), .ZN(n400) );
  INV_X1 U542 ( .A(n404), .ZN(n696) );
  OR2_X2 U543 ( .A1(n605), .A2(n370), .ZN(n404) );
  INV_X1 U544 ( .A(n584), .ZN(n409) );
  NOR2_X1 U545 ( .A1(n584), .A2(n643), .ZN(n573) );
  NAND2_X1 U546 ( .A1(n647), .A2(n646), .ZN(n643) );
  XNOR2_X1 U547 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U548 ( .A(n499), .B(n469), .ZN(n454) );
  NOR2_X1 U549 ( .A1(n703), .A2(n615), .ZN(n456) );
  INV_X1 U550 ( .A(KEYINPUT40), .ZN(n413) );
  NAND2_X1 U551 ( .A1(n608), .A2(n599), .ZN(n414) );
  NAND2_X1 U552 ( .A1(n628), .A2(n615), .ZN(n415) );
  NAND2_X1 U553 ( .A1(n573), .A2(n418), .ZN(n541) );
  XNOR2_X1 U554 ( .A(n419), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X2 U555 ( .A(n456), .B(n346), .ZN(n598) );
  NAND2_X1 U556 ( .A1(n625), .A2(n420), .ZN(n626) );
  XOR2_X1 U557 ( .A(KEYINPUT25), .B(KEYINPUT93), .Z(n429) );
  AND2_X1 U558 ( .A1(n462), .A2(n632), .ZN(n463) );
  INV_X1 U559 ( .A(G472), .ZN(n502) );
  INV_X1 U560 ( .A(KEYINPUT71), .ZN(n576) );
  NOR2_X1 U561 ( .A1(G952), .A2(n406), .ZN(n715) );
  XNOR2_X1 U562 ( .A(n626), .B(KEYINPUT123), .ZN(G54) );
  INV_X1 U563 ( .A(n464), .ZN(n615) );
  XOR2_X1 U564 ( .A(KEYINPUT75), .B(KEYINPUT87), .Z(n431) );
  NAND2_X1 U565 ( .A1(G210), .A2(n457), .ZN(n430) );
  XNOR2_X1 U566 ( .A(n431), .B(n430), .ZN(n432) );
  NAND2_X1 U567 ( .A1(G224), .A2(n406), .ZN(n433) );
  XNOR2_X1 U568 ( .A(n434), .B(n433), .ZN(n448) );
  INV_X1 U569 ( .A(G107), .ZN(n435) );
  NAND2_X1 U570 ( .A1(G104), .A2(n435), .ZN(n438) );
  INV_X1 U571 ( .A(G104), .ZN(n436) );
  NAND2_X1 U572 ( .A1(n436), .A2(G107), .ZN(n437) );
  NAND2_X1 U573 ( .A1(n438), .A2(n437), .ZN(n442) );
  INV_X1 U574 ( .A(n442), .ZN(n440) );
  INV_X1 U575 ( .A(n441), .ZN(n439) );
  NAND2_X1 U576 ( .A1(n440), .A2(n439), .ZN(n444) );
  NAND2_X1 U577 ( .A1(n442), .A2(n441), .ZN(n443) );
  XNOR2_X1 U578 ( .A(n483), .B(n445), .ZN(n446) );
  XNOR2_X1 U579 ( .A(n448), .B(n447), .ZN(n455) );
  XNOR2_X1 U580 ( .A(KEYINPUT4), .B(KEYINPUT64), .ZN(n733) );
  XNOR2_X1 U581 ( .A(G101), .B(n733), .ZN(n489) );
  INV_X1 U582 ( .A(n449), .ZN(n451) );
  XNOR2_X1 U583 ( .A(G119), .B(G116), .ZN(n450) );
  XNOR2_X1 U584 ( .A(n451), .B(n450), .ZN(n453) );
  XOR2_X1 U585 ( .A(KEYINPUT67), .B(KEYINPUT84), .Z(n452) );
  XNOR2_X1 U586 ( .A(n454), .B(n455), .ZN(n703) );
  NAND2_X1 U587 ( .A1(n457), .A2(G214), .ZN(n458) );
  XNOR2_X1 U588 ( .A(KEYINPUT88), .B(n458), .ZN(n604) );
  NOR2_X1 U589 ( .A1(G898), .A2(n406), .ZN(n459) );
  XOR2_X1 U590 ( .A(KEYINPUT89), .B(n459), .Z(n719) );
  NAND2_X1 U591 ( .A1(n719), .A2(G902), .ZN(n460) );
  NAND2_X1 U592 ( .A1(G952), .A2(n406), .ZN(n569) );
  NAND2_X1 U593 ( .A1(n460), .A2(n569), .ZN(n462) );
  XNOR2_X1 U594 ( .A(KEYINPUT14), .B(n461), .ZN(n632) );
  INV_X1 U595 ( .A(n632), .ZN(n570) );
  NAND2_X1 U596 ( .A1(G234), .A2(n464), .ZN(n465) );
  XNOR2_X1 U597 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U598 ( .A(KEYINPUT91), .B(n467), .ZN(n477) );
  NAND2_X1 U599 ( .A1(G221), .A2(n477), .ZN(n468) );
  XOR2_X1 U600 ( .A(KEYINPUT21), .B(n468), .Z(n646) );
  XOR2_X1 U601 ( .A(G137), .B(G140), .Z(n486) );
  XNOR2_X1 U602 ( .A(KEYINPUT10), .B(n469), .ZN(n519) );
  XNOR2_X1 U603 ( .A(n486), .B(n519), .ZN(n731) );
  XNOR2_X1 U604 ( .A(G119), .B(G128), .ZN(n470) );
  XNOR2_X1 U605 ( .A(n348), .B(n470), .ZN(n471) );
  XNOR2_X1 U606 ( .A(n471), .B(n347), .ZN(n475) );
  NAND2_X1 U607 ( .A1(n406), .A2(G234), .ZN(n473) );
  XNOR2_X1 U608 ( .A(n473), .B(n472), .ZN(n509) );
  NAND2_X1 U609 ( .A1(G221), .A2(n509), .ZN(n474) );
  NAND2_X1 U610 ( .A1(G217), .A2(n477), .ZN(n478) );
  NAND2_X1 U611 ( .A1(G134), .A2(n482), .ZN(n485) );
  XOR2_X1 U612 ( .A(n486), .B(KEYINPUT73), .Z(n488) );
  NAND2_X1 U613 ( .A1(G227), .A2(n406), .ZN(n487) );
  XNOR2_X1 U614 ( .A(n488), .B(n487), .ZN(n490) );
  XNOR2_X1 U615 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U616 ( .A(n495), .B(n494), .ZN(n501) );
  NAND2_X1 U617 ( .A1(n520), .A2(G210), .ZN(n496) );
  XNOR2_X1 U618 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U619 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U620 ( .A(n501), .B(n500), .ZN(n671) );
  NOR2_X1 U621 ( .A1(n671), .A2(G902), .ZN(n503) );
  INV_X1 U622 ( .A(n601), .ZN(n534) );
  XNOR2_X1 U623 ( .A(KEYINPUT101), .B(G478), .ZN(n515) );
  INV_X1 U624 ( .A(n504), .ZN(n508) );
  XNOR2_X1 U625 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U626 ( .A(n508), .B(n507), .Z(n513) );
  XOR2_X1 U627 ( .A(KEYINPUT9), .B(KEYINPUT100), .Z(n511) );
  NAND2_X1 U628 ( .A1(G217), .A2(n509), .ZN(n510) );
  XNOR2_X1 U629 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U630 ( .A(n513), .B(n512), .ZN(n710) );
  NOR2_X1 U631 ( .A1(G902), .A2(n710), .ZN(n514) );
  XNOR2_X1 U632 ( .A(n515), .B(n514), .ZN(n538) );
  XNOR2_X1 U633 ( .A(KEYINPUT13), .B(G475), .ZN(n528) );
  XNOR2_X1 U634 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U635 ( .A(n519), .B(n518), .ZN(n526) );
  XOR2_X1 U636 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n522) );
  NAND2_X1 U637 ( .A1(G214), .A2(n520), .ZN(n521) );
  XNOR2_X1 U638 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U639 ( .A(n526), .B(n525), .ZN(n705) );
  NOR2_X1 U640 ( .A1(G902), .A2(n705), .ZN(n527) );
  XNOR2_X1 U641 ( .A(n528), .B(n527), .ZN(n536) );
  NAND2_X1 U642 ( .A1(n538), .A2(n536), .ZN(n591) );
  INV_X1 U643 ( .A(KEYINPUT83), .ZN(n529) );
  NOR2_X1 U644 ( .A1(n538), .A2(n536), .ZN(n635) );
  AND2_X1 U645 ( .A1(n646), .A2(n635), .ZN(n531) );
  XNOR2_X1 U646 ( .A(KEYINPUT104), .B(n531), .ZN(n532) );
  INV_X1 U647 ( .A(n647), .ZN(n554) );
  NOR2_X1 U648 ( .A1(n534), .A2(n554), .ZN(n535) );
  NAND2_X1 U649 ( .A1(n551), .A2(n535), .ZN(n673) );
  XNOR2_X1 U650 ( .A(KEYINPUT99), .B(n536), .ZN(n537) );
  NAND2_X1 U651 ( .A1(n538), .A2(n537), .ZN(n682) );
  XOR2_X1 U652 ( .A(KEYINPUT102), .B(n682), .Z(n607) );
  NOR2_X1 U653 ( .A1(n599), .A2(n607), .ZN(n539) );
  XNOR2_X1 U654 ( .A(KEYINPUT103), .B(n539), .ZN(n637) );
  INV_X1 U655 ( .A(n637), .ZN(n594) );
  INV_X1 U656 ( .A(n540), .ZN(n543) );
  NOR2_X1 U657 ( .A1(n543), .A2(n541), .ZN(n677) );
  NAND2_X1 U658 ( .A1(n416), .A2(n542), .ZN(n642) );
  NOR2_X1 U659 ( .A1(n543), .A2(n642), .ZN(n545) );
  XNOR2_X1 U660 ( .A(KEYINPUT97), .B(KEYINPUT31), .ZN(n544) );
  XNOR2_X1 U661 ( .A(n545), .B(n544), .ZN(n694) );
  NOR2_X1 U662 ( .A1(n677), .A2(n694), .ZN(n546) );
  OR2_X1 U663 ( .A1(n594), .A2(n546), .ZN(n547) );
  NAND2_X1 U664 ( .A1(n673), .A2(n547), .ZN(n548) );
  XNOR2_X1 U665 ( .A(n550), .B(KEYINPUT82), .ZN(n562) );
  XNOR2_X1 U666 ( .A(n551), .B(KEYINPUT105), .ZN(n552) );
  NAND2_X1 U667 ( .A1(n554), .A2(n601), .ZN(n555) );
  NAND2_X1 U668 ( .A1(n610), .A2(n557), .ZN(n558) );
  NAND2_X1 U669 ( .A1(n559), .A2(n741), .ZN(n560) );
  INV_X1 U670 ( .A(n604), .ZN(n634) );
  XNOR2_X1 U671 ( .A(KEYINPUT109), .B(KEYINPUT30), .ZN(n564) );
  XNOR2_X1 U672 ( .A(n565), .B(n564), .ZN(n575) );
  NAND2_X1 U673 ( .A1(G953), .A2(G902), .ZN(n566) );
  NOR2_X1 U674 ( .A1(n570), .A2(n566), .ZN(n567) );
  XNOR2_X1 U675 ( .A(n567), .B(KEYINPUT107), .ZN(n568) );
  NOR2_X1 U676 ( .A1(G900), .A2(n568), .ZN(n572) );
  NOR2_X1 U677 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U678 ( .A1(n572), .A2(n571), .ZN(n580) );
  XNOR2_X1 U679 ( .A(n577), .B(n576), .ZN(n589) );
  XNOR2_X1 U680 ( .A(KEYINPUT68), .B(KEYINPUT38), .ZN(n578) );
  NAND2_X1 U681 ( .A1(n589), .A2(n585), .ZN(n579) );
  XOR2_X1 U682 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n587) );
  NOR2_X1 U683 ( .A1(n580), .A2(n647), .ZN(n581) );
  NAND2_X1 U684 ( .A1(n581), .A2(n646), .ZN(n600) );
  XOR2_X1 U685 ( .A(KEYINPUT28), .B(n582), .Z(n583) );
  NOR2_X1 U686 ( .A1(n584), .A2(n583), .ZN(n593) );
  NAND2_X1 U687 ( .A1(n593), .A2(n665), .ZN(n586) );
  NAND2_X1 U688 ( .A1(n589), .A2(n598), .ZN(n590) );
  NOR2_X1 U689 ( .A1(n591), .A2(n590), .ZN(n686) );
  NAND2_X1 U690 ( .A1(n593), .A2(n592), .ZN(n687) );
  NOR2_X1 U691 ( .A1(n687), .A2(n594), .ZN(n595) );
  NOR2_X1 U692 ( .A1(n686), .A2(n596), .ZN(n597) );
  INV_X1 U693 ( .A(n598), .ZN(n612) );
  XNOR2_X1 U694 ( .A(n599), .B(KEYINPUT106), .ZN(n690) );
  INV_X1 U695 ( .A(n690), .ZN(n688) );
  AND2_X1 U696 ( .A1(n608), .A2(n607), .ZN(n699) );
  INV_X1 U697 ( .A(n699), .ZN(n614) );
  OR2_X1 U698 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U699 ( .A(KEYINPUT43), .B(n611), .ZN(n613) );
  NAND2_X1 U700 ( .A1(n613), .A2(n612), .ZN(n701) );
  XOR2_X1 U701 ( .A(KEYINPUT79), .B(n615), .Z(n616) );
  NAND2_X1 U702 ( .A1(n616), .A2(KEYINPUT2), .ZN(n617) );
  XNOR2_X1 U703 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n622) );
  XNOR2_X1 U704 ( .A(n620), .B(KEYINPUT57), .ZN(n621) );
  XNOR2_X1 U705 ( .A(n622), .B(n621), .ZN(n623) );
  XOR2_X1 U706 ( .A(KEYINPUT2), .B(KEYINPUT77), .Z(n627) );
  XNOR2_X1 U707 ( .A(n629), .B(KEYINPUT76), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n632), .A2(G952), .ZN(n663) );
  NAND2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U711 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U712 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n664), .A2(n641), .ZN(n659) );
  INV_X1 U714 ( .A(n642), .ZN(n655) );
  NAND2_X1 U715 ( .A1(n370), .A2(n643), .ZN(n645) );
  XNOR2_X1 U716 ( .A(KEYINPUT50), .B(n645), .ZN(n651) );
  XOR2_X1 U717 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n649) );
  OR2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U719 ( .A(n649), .B(n648), .ZN(n650) );
  NAND2_X1 U720 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U721 ( .A1(n416), .A2(n652), .ZN(n654) );
  NOR2_X1 U722 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U723 ( .A(KEYINPUT51), .B(n656), .ZN(n657) );
  NAND2_X1 U724 ( .A1(n657), .A2(n665), .ZN(n658) );
  NAND2_X1 U725 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U726 ( .A(n660), .B(KEYINPUT119), .ZN(n661) );
  XNOR2_X1 U727 ( .A(n661), .B(KEYINPUT52), .ZN(n662) );
  NOR2_X1 U728 ( .A1(n663), .A2(n662), .ZN(n667) );
  AND2_X1 U729 ( .A1(n664), .A2(n665), .ZN(n666) );
  NOR2_X1 U730 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U731 ( .A(KEYINPUT120), .B(n668), .ZN(n669) );
  INV_X1 U732 ( .A(KEYINPUT53), .ZN(n670) );
  XNOR2_X1 U733 ( .A(KEYINPUT111), .B(KEYINPUT62), .ZN(n672) );
  XNOR2_X1 U734 ( .A(G101), .B(n673), .ZN(G3) );
  XOR2_X1 U735 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n675) );
  NAND2_X1 U736 ( .A1(n677), .A2(n690), .ZN(n674) );
  XNOR2_X1 U737 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U738 ( .A(G104), .B(n676), .ZN(G6) );
  XOR2_X1 U739 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n679) );
  INV_X1 U740 ( .A(n682), .ZN(n693) );
  NAND2_X1 U741 ( .A1(n677), .A2(n693), .ZN(n678) );
  XNOR2_X1 U742 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U743 ( .A(G107), .B(n680), .ZN(G9) );
  XOR2_X1 U744 ( .A(n681), .B(G110), .Z(G12) );
  NOR2_X1 U745 ( .A1(n682), .A2(n687), .ZN(n684) );
  XNOR2_X1 U746 ( .A(KEYINPUT114), .B(KEYINPUT29), .ZN(n683) );
  XNOR2_X1 U747 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U748 ( .A(G128), .B(n685), .ZN(G30) );
  XOR2_X1 U749 ( .A(G143), .B(n686), .Z(G45) );
  NOR2_X1 U750 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U751 ( .A(G146), .B(n689), .Z(G48) );
  XOR2_X1 U752 ( .A(G113), .B(KEYINPUT115), .Z(n692) );
  NAND2_X1 U753 ( .A1(n694), .A2(n690), .ZN(n691) );
  XNOR2_X1 U754 ( .A(n692), .B(n691), .ZN(G15) );
  NAND2_X1 U755 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U756 ( .A(n695), .B(G116), .ZN(G18) );
  XNOR2_X1 U757 ( .A(n696), .B(KEYINPUT116), .ZN(n697) );
  XNOR2_X1 U758 ( .A(n697), .B(KEYINPUT37), .ZN(n698) );
  XNOR2_X1 U759 ( .A(G125), .B(n698), .ZN(G27) );
  XNOR2_X1 U760 ( .A(G134), .B(n699), .ZN(n700) );
  XNOR2_X1 U761 ( .A(n700), .B(KEYINPUT117), .ZN(G36) );
  XNOR2_X1 U762 ( .A(G140), .B(n701), .ZN(G42) );
  XNOR2_X1 U763 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n702) );
  XOR2_X1 U764 ( .A(n705), .B(KEYINPUT59), .Z(n707) );
  XNOR2_X1 U765 ( .A(n708), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U766 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U767 ( .A1(n715), .A2(n711), .ZN(G63) );
  XNOR2_X1 U768 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U769 ( .A1(n715), .A2(n714), .ZN(G66) );
  XNOR2_X1 U770 ( .A(n716), .B(G101), .ZN(n718) );
  XNOR2_X1 U771 ( .A(n717), .B(n718), .ZN(n720) );
  NOR2_X1 U772 ( .A1(n720), .A2(n719), .ZN(n729) );
  NAND2_X1 U773 ( .A1(n721), .A2(n406), .ZN(n722) );
  XNOR2_X1 U774 ( .A(n722), .B(KEYINPUT124), .ZN(n726) );
  NAND2_X1 U775 ( .A1(G953), .A2(G224), .ZN(n723) );
  XNOR2_X1 U776 ( .A(KEYINPUT61), .B(n723), .ZN(n724) );
  NAND2_X1 U777 ( .A1(n724), .A2(G898), .ZN(n725) );
  NAND2_X1 U778 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U779 ( .A(n727), .B(KEYINPUT125), .Z(n728) );
  XNOR2_X1 U780 ( .A(n729), .B(n728), .ZN(G69) );
  XNOR2_X1 U781 ( .A(n731), .B(n730), .ZN(n732) );
  XNOR2_X1 U782 ( .A(n733), .B(n732), .ZN(n735) );
  NAND2_X1 U783 ( .A1(n734), .A2(n406), .ZN(n739) );
  XNOR2_X1 U784 ( .A(G227), .B(n735), .ZN(n736) );
  NAND2_X1 U785 ( .A1(n736), .A2(G900), .ZN(n737) );
  NAND2_X1 U786 ( .A1(n737), .A2(G953), .ZN(n738) );
  NAND2_X1 U787 ( .A1(n739), .A2(n738), .ZN(G72) );
  XOR2_X1 U788 ( .A(G137), .B(n740), .Z(G39) );
  XOR2_X1 U789 ( .A(n741), .B(G122), .Z(G24) );
  XOR2_X1 U790 ( .A(G119), .B(n742), .Z(G21) );
  XOR2_X1 U791 ( .A(n743), .B(G131), .Z(G33) );
endmodule

