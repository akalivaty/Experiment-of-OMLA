//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1299, new_n1300, new_n1301, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n212));
  XNOR2_X1  g0012(.A(new_n211), .B(new_n212), .ZN(new_n213));
  AND2_X1   g0013(.A1(KEYINPUT65), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(KEYINPUT65), .A2(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI22_X1  g0024(.A1(new_n222), .A2(new_n223), .B1(new_n206), .B2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT68), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT67), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n228));
  AOI22_X1  g0028(.A1(new_n225), .A2(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT66), .B(G77), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G244), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n229), .B(new_n232), .C1(new_n227), .C2(new_n228), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G116), .A2(G270), .ZN(new_n234));
  AOI22_X1  g0034(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n234), .B(new_n235), .C1(new_n225), .C2(new_n226), .ZN(new_n236));
  OAI21_X1  g0036(.A(new_n209), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  OAI211_X1 g0037(.A(new_n213), .B(new_n221), .C1(new_n237), .C2(KEYINPUT1), .ZN(new_n238));
  AOI21_X1  g0038(.A(new_n238), .B1(KEYINPUT1), .B2(new_n237), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G264), .B(G270), .Z(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT69), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G68), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G68), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n256), .A2(G50), .B1(G20), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n216), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G77), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n217), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT11), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT72), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n267), .A2(KEYINPUT72), .A3(G13), .A4(G20), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OR3_X1    g0072(.A1(new_n272), .A2(KEYINPUT12), .A3(G68), .ZN(new_n273));
  OAI21_X1  g0073(.A(KEYINPUT12), .B1(new_n272), .B2(G68), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n263), .B1(new_n270), .B2(new_n271), .ZN(new_n276));
  INV_X1    g0076(.A(G20), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n276), .B(G68), .C1(G1), .C2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n261), .A2(KEYINPUT11), .A3(new_n263), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n266), .A2(new_n275), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT14), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT13), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G226), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n223), .A2(G1698), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n284), .A2(new_n287), .A3(new_n289), .A4(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G97), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G41), .ZN(new_n296));
  INV_X1    g0096(.A(G45), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(G1), .A2(G13), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G41), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n267), .A2(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OR2_X1    g0101(.A1(KEYINPUT70), .A2(G45), .ZN(new_n302));
  NAND2_X1  g0102(.A1(KEYINPUT70), .A2(G45), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(new_n296), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n267), .A2(G274), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n301), .A2(G238), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n282), .B1(new_n295), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n300), .A2(G1), .A3(G13), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n291), .B2(new_n292), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(G238), .A3(new_n311), .ZN(new_n312));
  AND2_X1   g0112(.A1(KEYINPUT70), .A2(G45), .ZN(new_n313));
  NOR2_X1   g0113(.A1(KEYINPUT70), .A2(G45), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n313), .A2(new_n314), .A3(G41), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n312), .B1(new_n315), .B2(new_n305), .ZN(new_n316));
  NOR3_X1   g0116(.A1(new_n310), .A2(new_n316), .A3(KEYINPUT13), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n281), .B(G169), .C1(new_n308), .C2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n295), .A2(new_n282), .A3(new_n307), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT13), .B1(new_n310), .B2(new_n316), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n320), .A3(G179), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n320), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n281), .B1(new_n323), .B2(G169), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n280), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT3), .B(G33), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(G238), .A3(G1698), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(G232), .A3(new_n286), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n284), .A2(new_n289), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G107), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n327), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n294), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n304), .A2(new_n306), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n309), .A2(G244), .A3(new_n311), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT73), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n333), .A2(KEYINPUT73), .A3(new_n334), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n332), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G200), .ZN(new_n340));
  INV_X1    g0140(.A(G190), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT15), .B(G87), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n259), .A2(new_n342), .B1(new_n230), .B2(new_n216), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n277), .A2(new_n288), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT74), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n222), .A2(KEYINPUT8), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT8), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G58), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n344), .A2(KEYINPUT74), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n346), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n263), .B1(new_n343), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT75), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n270), .A2(new_n271), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n260), .B1(new_n267), .B2(G20), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n230), .A2(new_n355), .B1(new_n276), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n353), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n354), .B1(new_n353), .B2(new_n357), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n340), .B1(new_n341), .B2(new_n339), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n323), .A2(new_n341), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(new_n280), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n323), .A2(G200), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G169), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n339), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n332), .A2(new_n337), .A3(new_n368), .A4(new_n338), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n353), .A2(new_n357), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n325), .A2(new_n361), .A3(new_n365), .A4(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(G222), .A2(G1698), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n286), .A2(G223), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n326), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n375), .B(new_n294), .C1(new_n231), .C2(new_n326), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n301), .A2(G226), .B1(new_n304), .B2(new_n306), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(G179), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n366), .B2(new_n378), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n355), .A2(new_n202), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n202), .B1(new_n267), .B2(G20), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n276), .A2(new_n382), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n263), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT71), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n347), .A2(new_n349), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n222), .A2(KEYINPUT71), .A3(KEYINPUT8), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n387), .A2(G33), .A3(new_n216), .A4(new_n388), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n256), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n385), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n384), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n380), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT9), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n384), .A2(new_n395), .A3(new_n392), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n381), .A2(new_n383), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT9), .B1(new_n397), .B2(new_n391), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n378), .A2(new_n341), .ZN(new_n400));
  INV_X1    g0200(.A(G200), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(new_n376), .B2(new_n377), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT10), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n399), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n404), .B1(new_n399), .B2(new_n403), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n394), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n372), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n387), .A2(new_n388), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n267), .B2(G20), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n276), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n355), .A2(new_n409), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g0213(.A(G58), .B(G68), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(G20), .B1(G159), .B2(new_n256), .ZN(new_n415));
  AOI21_X1  g0215(.A(G20), .B1(new_n284), .B2(new_n289), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT7), .ZN(new_n417));
  OAI21_X1  g0217(.A(G68), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OR2_X1    g0218(.A1(KEYINPUT65), .A2(G20), .ZN(new_n419));
  NAND2_X1  g0219(.A1(KEYINPUT65), .A2(G20), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n421), .A2(new_n326), .ZN(new_n422));
  OAI211_X1 g0222(.A(KEYINPUT16), .B(new_n415), .C1(new_n418), .C2(new_n422), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n423), .A2(new_n263), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT16), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT76), .B1(new_n288), .B2(KEYINPUT3), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT76), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(new_n283), .A3(G33), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n428), .A3(new_n289), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n214), .A2(new_n215), .A3(new_n417), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n417), .B1(new_n326), .B2(G20), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n257), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n415), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n425), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n413), .B1(new_n424), .B2(new_n435), .ZN(new_n436));
  OR2_X1    g0236(.A1(G223), .A2(G1698), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n285), .A2(G1698), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n284), .A2(new_n437), .A3(new_n289), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(G33), .A2(G87), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n309), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n309), .A2(G232), .A3(new_n311), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(new_n315), .B2(new_n305), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G179), .ZN(new_n445));
  OAI21_X1  g0245(.A(G169), .B1(new_n441), .B2(new_n443), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT18), .B1(new_n436), .B2(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n410), .A2(new_n276), .B1(new_n355), .B2(new_n409), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n431), .A2(new_n432), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(G68), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT16), .B1(new_n452), .B2(new_n415), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n423), .A2(new_n263), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT18), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n456), .A3(new_n447), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n449), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT17), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n439), .A2(new_n440), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n294), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n301), .A2(G232), .B1(new_n304), .B2(new_n306), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT77), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .A4(new_n341), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n401), .B1(new_n441), .B2(new_n443), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n463), .B1(new_n444), .B2(new_n341), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n459), .B1(new_n455), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n461), .A2(new_n341), .A3(new_n462), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT77), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(new_n465), .A3(new_n464), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n435), .A2(new_n263), .A3(new_n423), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n472), .A2(new_n473), .A3(KEYINPUT17), .A4(new_n450), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n458), .A2(new_n475), .A3(KEYINPUT78), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n449), .A2(new_n469), .A3(new_n457), .A4(new_n474), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT78), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n408), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  OR2_X1    g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  NAND2_X1  g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  AOI211_X1 g0282(.A(G1), .B(new_n297), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G274), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n481), .A2(new_n482), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n297), .A2(G1), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(G270), .A3(new_n309), .ZN(new_n488));
  INV_X1    g0288(.A(G303), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n329), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n286), .A2(G264), .ZN(new_n491));
  NOR2_X1   g0291(.A1(G257), .A2(G1698), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n284), .B(new_n289), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n490), .A2(new_n493), .A3(new_n294), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n484), .A2(new_n488), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G169), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n288), .A2(G97), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G283), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n419), .A2(new_n498), .A3(new_n420), .A4(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G116), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n262), .A2(new_n217), .B1(G20), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT20), .ZN(new_n504));
  OR2_X1    g0304(.A1(new_n504), .A2(KEYINPUT85), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(KEYINPUT85), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n267), .A2(G33), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n272), .A2(G116), .A3(new_n385), .A4(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n270), .A2(new_n501), .A3(new_n271), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n500), .A2(KEYINPUT85), .A3(new_n502), .A4(new_n504), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n507), .A2(new_n509), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT86), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n512), .A2(new_n513), .ZN(new_n515));
  OAI211_X1 g0315(.A(KEYINPUT21), .B(new_n497), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  AND4_X1   g0316(.A1(G179), .A2(new_n484), .A3(new_n488), .A4(new_n494), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n514), .B2(new_n515), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n509), .A2(new_n510), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n520), .A2(KEYINPUT86), .A3(new_n511), .A4(new_n507), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n512), .A2(new_n513), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT21), .B1(new_n523), .B2(new_n497), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n495), .A2(G200), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n341), .B2(new_n495), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n519), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n419), .A2(new_n420), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT87), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT23), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .A4(new_n206), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n206), .ZN(new_n533));
  OAI21_X1  g0333(.A(KEYINPUT87), .B1(new_n216), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n531), .B1(G20), .B2(new_n206), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G116), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(G20), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n532), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n216), .A2(new_n326), .A3(G87), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT22), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT22), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n216), .A2(new_n326), .A3(new_n542), .A4(G87), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT24), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n539), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n545), .B1(new_n539), .B2(new_n544), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n263), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n272), .A2(new_n385), .A3(new_n508), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT80), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n276), .A2(KEYINPUT80), .A3(new_n508), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(KEYINPUT25), .B1(new_n355), .B2(new_n206), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n355), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n553), .A2(new_n206), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n487), .A2(new_n309), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n484), .B1(new_n558), .B2(new_n224), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n284), .A2(new_n289), .A3(G257), .A4(G1698), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT88), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT88), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n326), .A2(new_n562), .A3(G257), .A4(G1698), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n284), .A2(new_n289), .A3(G250), .A4(new_n286), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G33), .A2(G294), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n561), .A2(new_n563), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n309), .B1(new_n566), .B2(KEYINPUT89), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n564), .A2(new_n565), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT89), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n568), .A2(new_n569), .A3(new_n561), .A4(new_n563), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n559), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n548), .A2(new_n557), .B1(new_n368), .B2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n564), .B(new_n565), .C1(new_n560), .C2(KEYINPUT88), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n560), .A2(KEYINPUT88), .ZN(new_n574));
  OAI21_X1  g0374(.A(KEYINPUT89), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(new_n294), .A3(new_n570), .ZN(new_n576));
  INV_X1    g0376(.A(new_n559), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n366), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n539), .A2(new_n544), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT24), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n539), .A2(new_n544), .A3(new_n545), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n556), .B1(new_n583), .B2(new_n263), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n576), .A2(new_n341), .A3(new_n577), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n571), .B2(G200), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n572), .A2(new_n579), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n342), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n272), .A2(new_n588), .ZN(new_n589));
  OR2_X1    g0389(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n590));
  NAND2_X1  g0390(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n292), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI22_X1  g0392(.A1(new_n592), .A2(new_n529), .B1(G87), .B2(new_n207), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n216), .A2(new_n326), .A3(G68), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n419), .A2(G33), .A3(G97), .A4(new_n420), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(new_n590), .A3(new_n591), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n589), .B1(new_n597), .B2(new_n263), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n551), .A2(new_n552), .A3(G87), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n284), .A2(new_n289), .A3(G238), .A4(new_n286), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n284), .A2(new_n289), .A3(G244), .A4(G1698), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n602), .A3(new_n536), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n294), .ZN(new_n604));
  OAI21_X1  g0404(.A(G250), .B1(new_n297), .B2(G1), .ZN(new_n605));
  OAI22_X1  g0405(.A1(new_n294), .A2(new_n605), .B1(new_n297), .B2(new_n305), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT82), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n604), .A2(KEYINPUT82), .A3(new_n607), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(G190), .A3(new_n611), .ZN(new_n612));
  AOI211_X1 g0412(.A(new_n609), .B(new_n606), .C1(new_n603), .C2(new_n294), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT82), .B1(new_n604), .B2(new_n607), .ZN(new_n614));
  OAI21_X1  g0414(.A(G200), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n600), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n610), .A2(new_n368), .A3(new_n611), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n366), .B1(new_n613), .B2(new_n614), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n597), .A2(new_n263), .ZN(new_n620));
  INV_X1    g0420(.A(new_n589), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n551), .A2(new_n552), .A3(new_n588), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT84), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT84), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n551), .A2(new_n552), .A3(new_n625), .A4(new_n588), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n622), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n616), .B1(new_n619), .B2(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n284), .A2(new_n289), .A3(G244), .A4(new_n286), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT4), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT81), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n326), .A2(G244), .A3(new_n286), .A4(new_n631), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n326), .A2(G250), .A3(G1698), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n633), .A2(new_n634), .A3(new_n499), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n294), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n483), .A2(new_n294), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G257), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n637), .A2(new_n484), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G200), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n551), .A2(new_n552), .A3(G97), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n272), .A2(G97), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n256), .A2(G77), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT6), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT79), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT79), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT6), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n205), .B2(G107), .ZN(new_n650));
  NAND2_X1  g0450(.A1(G97), .A2(G107), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n207), .A2(new_n646), .A3(new_n648), .A4(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n650), .A2(new_n529), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n329), .A2(new_n277), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n654), .A2(new_n417), .B1(new_n429), .B2(new_n430), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n644), .B(new_n653), .C1(new_n655), .C2(new_n206), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n643), .B1(new_n656), .B2(new_n263), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n636), .A2(new_n294), .B1(new_n638), .B2(G257), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n658), .A2(G190), .A3(new_n484), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n641), .A2(new_n642), .A3(new_n657), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n653), .A2(new_n644), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n206), .B1(new_n431), .B2(new_n432), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n263), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n643), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n642), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n640), .A2(new_n366), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n658), .A2(new_n368), .A3(new_n484), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n660), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n628), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n480), .A2(new_n528), .A3(new_n587), .A4(new_n670), .ZN(new_n671));
  XOR2_X1   g0471(.A(new_n671), .B(KEYINPUT90), .Z(G372));
  NAND2_X1  g0472(.A1(new_n371), .A2(KEYINPUT91), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT91), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n367), .A2(new_n674), .A3(new_n369), .A4(new_n370), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n365), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n325), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT92), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n475), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n677), .A2(KEYINPUT92), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n458), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n405), .A2(new_n406), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n681), .A2(new_n682), .B1(new_n393), .B2(new_n380), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT26), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n608), .A2(G200), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n600), .A2(new_n612), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n608), .A2(new_n366), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n617), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n686), .B1(new_n627), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n684), .B1(new_n689), .B2(new_n668), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n624), .A2(new_n626), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n598), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(new_n618), .A3(new_n617), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n693), .A2(KEYINPUT26), .A3(new_n694), .A4(new_n616), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n496), .B1(new_n521), .B2(new_n522), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n697), .A2(KEYINPUT21), .B1(new_n523), .B2(new_n517), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n571), .A2(new_n368), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n385), .B1(new_n581), .B2(new_n582), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n579), .B(new_n699), .C1(new_n700), .C2(new_n556), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n523), .A2(new_n497), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT21), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n698), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n598), .A2(new_n599), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n613), .A2(new_n614), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n706), .B1(G190), .B2(new_n707), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n584), .A2(new_n586), .B1(new_n708), .B2(new_n685), .ZN(new_n709));
  INV_X1    g0509(.A(new_n669), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n705), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n688), .A2(new_n627), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n696), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n480), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n683), .A2(new_n715), .ZN(G369));
  NAND2_X1  g0516(.A1(new_n698), .A2(new_n704), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n216), .A2(new_n267), .A3(G13), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n718), .A2(KEYINPUT27), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(KEYINPUT27), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(G213), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G343), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n724), .B1(new_n522), .B2(new_n521), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT93), .B1(new_n717), .B2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n528), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n726), .B1(new_n727), .B2(new_n725), .ZN(new_n728));
  XOR2_X1   g0528(.A(KEYINPUT94), .B(G330), .Z(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n717), .A2(KEYINPUT93), .A3(new_n725), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n728), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n587), .B1(new_n584), .B2(new_n724), .ZN(new_n733));
  INV_X1    g0533(.A(new_n701), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n723), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n723), .B1(new_n698), .B2(new_n704), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n587), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n734), .A2(new_n724), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n738), .A2(new_n742), .ZN(G399));
  INV_X1    g0543(.A(new_n210), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G41), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n267), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n746), .A2(new_n747), .B1(new_n220), .B2(new_n745), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT28), .Z(new_n749));
  INV_X1    g0549(.A(KEYINPUT30), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n610), .A2(new_n658), .A3(new_n517), .A4(new_n611), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n750), .B1(new_n751), .B2(new_n578), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n658), .A2(new_n517), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n753), .A2(new_n571), .A3(KEYINPUT30), .A4(new_n707), .ZN(new_n754));
  AND3_X1   g0554(.A1(new_n608), .A2(new_n368), .A3(new_n495), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n578), .A2(new_n640), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n752), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n757), .A2(KEYINPUT31), .A3(new_n723), .ZN(new_n758));
  AOI21_X1  g0558(.A(KEYINPUT31), .B1(new_n757), .B2(new_n723), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n670), .A2(new_n528), .A3(new_n587), .A4(new_n724), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n730), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n689), .A2(new_n668), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(KEYINPUT95), .A3(KEYINPUT26), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT95), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n694), .B(new_n616), .C1(new_n627), .C2(new_n619), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n767), .B1(new_n768), .B2(new_n684), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n689), .A2(new_n684), .A3(new_n668), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n766), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n709), .A2(new_n710), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n712), .B1(new_n772), .B2(new_n705), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(KEYINPUT29), .A3(new_n724), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n714), .A2(new_n724), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT29), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n764), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n749), .B1(new_n779), .B2(G1), .ZN(G364));
  AOI21_X1  g0580(.A(new_n217), .B1(G20), .B2(new_n366), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n216), .A2(new_n368), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n782), .A2(new_n341), .A3(new_n401), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n784), .A2(KEYINPUT98), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(KEYINPUT98), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n782), .A2(G190), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G200), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n788), .A2(new_n231), .B1(G58), .B2(new_n790), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n791), .A2(KEYINPUT99), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(KEYINPUT99), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n216), .A2(G190), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G179), .A2(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G159), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT32), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n368), .A2(new_n401), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n794), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n216), .B1(G190), .B2(new_n795), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n801), .A2(new_n257), .B1(new_n802), .B2(new_n205), .ZN(new_n803));
  NOR4_X1   g0603(.A1(new_n277), .A2(new_n341), .A3(new_n401), .A4(G179), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G87), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n401), .A2(G179), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n794), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n326), .B(new_n805), .C1(new_n807), .C2(new_n206), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n789), .A2(new_n401), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n803), .B(new_n808), .C1(G50), .C2(new_n809), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n792), .A2(new_n793), .A3(new_n799), .A4(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT100), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n788), .A2(G311), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n790), .A2(G322), .ZN(new_n815));
  INV_X1    g0615(.A(new_n804), .ZN(new_n816));
  XOR2_X1   g0616(.A(KEYINPUT33), .B(G317), .Z(new_n817));
  OAI221_X1 g0617(.A(new_n329), .B1(new_n816), .B2(new_n489), .C1(new_n801), .C2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G326), .B2(new_n809), .ZN(new_n819));
  INV_X1    g0619(.A(G283), .ZN(new_n820));
  INV_X1    g0620(.A(G329), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n820), .A2(new_n807), .B1(new_n796), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n802), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n822), .B1(G294), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n814), .A2(new_n815), .A3(new_n819), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n813), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n811), .A2(new_n812), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n781), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(G13), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n529), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(G45), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n746), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(G13), .A2(G33), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(G20), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(new_n781), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n326), .A2(new_n210), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(KEYINPUT96), .B2(G355), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(KEYINPUT96), .B2(G355), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(G116), .B2(new_n210), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n254), .A2(G45), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT97), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n744), .A2(new_n326), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n313), .A2(new_n314), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(new_n220), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n842), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n828), .B(new_n833), .C1(new_n838), .C2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n728), .A2(new_n731), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n836), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n732), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(new_n833), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n852), .A2(new_n730), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n850), .A2(new_n854), .B1(new_n857), .B2(new_n858), .ZN(G396));
  NAND4_X1  g0659(.A1(new_n673), .A2(new_n370), .A3(new_n675), .A4(new_n723), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n723), .A2(new_n370), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n359), .A2(new_n360), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n340), .B1(new_n341), .B2(new_n339), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n371), .B(new_n861), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n776), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n361), .A2(new_n371), .A3(new_n724), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n714), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n833), .B1(new_n870), .B2(new_n763), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n763), .B2(new_n870), .ZN(new_n872));
  INV_X1    g0672(.A(new_n781), .ZN(new_n873));
  INV_X1    g0673(.A(new_n801), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n809), .A2(G137), .B1(new_n874), .B2(G150), .ZN(new_n875));
  INV_X1    g0675(.A(G143), .ZN(new_n876));
  INV_X1    g0676(.A(new_n790), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n875), .B1(new_n876), .B2(new_n877), .C1(new_n787), .C2(new_n797), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT34), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n807), .A2(new_n257), .ZN(new_n880));
  OAI221_X1 g0680(.A(new_n326), .B1(new_n816), .B2(new_n202), .C1(new_n222), .C2(new_n802), .ZN(new_n881));
  INV_X1    g0681(.A(new_n796), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n880), .B(new_n881), .C1(G132), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n788), .A2(G116), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n809), .A2(G303), .ZN(new_n886));
  INV_X1    g0686(.A(G87), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n887), .A2(new_n807), .B1(new_n801), .B2(new_n820), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(G311), .B2(new_n882), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n329), .B1(new_n816), .B2(new_n206), .C1(new_n205), .C2(new_n802), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(G294), .B2(new_n790), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n885), .A2(new_n886), .A3(new_n889), .A4(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n873), .B1(new_n884), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n781), .A2(new_n834), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n832), .B(new_n893), .C1(new_n260), .C2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n835), .B2(new_n865), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n872), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(G384));
  NOR2_X1   g0698(.A1(new_n830), .A2(new_n267), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n325), .A2(new_n723), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  INV_X1    g0702(.A(new_n721), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n455), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n477), .A2(KEYINPUT103), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n455), .A2(new_n447), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n472), .A2(new_n473), .A3(new_n450), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT37), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n907), .A2(new_n904), .A3(new_n911), .A4(new_n908), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n906), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT103), .B1(new_n477), .B2(new_n905), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n902), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT104), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n329), .A2(new_n216), .A3(new_n417), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n918), .B(G68), .C1(new_n417), .C2(new_n416), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT16), .B1(new_n919), .B2(new_n415), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n450), .B1(new_n454), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n903), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n447), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n908), .A2(new_n924), .A3(new_n922), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT37), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n477), .A2(new_n923), .B1(new_n926), .B2(new_n912), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT39), .B1(new_n927), .B2(KEYINPUT38), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n916), .A2(new_n917), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n477), .A2(new_n923), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n926), .A2(new_n912), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT38), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT38), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT39), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n917), .B1(new_n916), .B2(new_n928), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n901), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n458), .A2(new_n903), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n371), .A2(new_n723), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n714), .B2(new_n868), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n280), .A2(new_n723), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n325), .A2(new_n365), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n941), .B1(new_n325), .B2(new_n365), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT102), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n932), .B2(new_n933), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n930), .A2(new_n931), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n902), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT38), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n949), .A2(KEYINPUT102), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n938), .B1(new_n945), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n937), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n775), .A2(new_n480), .A3(new_n778), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n683), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n954), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n477), .A2(new_n905), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT103), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(new_n913), .A3(new_n906), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n932), .B1(new_n961), .B2(new_n902), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n865), .B1(new_n942), .B2(new_n943), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  AND4_X1   g0764(.A1(new_n528), .A2(new_n670), .A3(new_n587), .A4(new_n724), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n757), .A2(new_n723), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT31), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n757), .A2(KEYINPUT31), .A3(new_n723), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n964), .B(KEYINPUT40), .C1(new_n965), .C2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n962), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n964), .B1(new_n965), .B2(new_n970), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NOR3_X1   g0774(.A1(new_n932), .A2(new_n933), .A3(new_n946), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT102), .B1(new_n949), .B2(new_n950), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT40), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n972), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n480), .A2(new_n762), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(new_n980), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n981), .A2(new_n730), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n899), .B1(new_n957), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n957), .B2(new_n983), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n650), .A2(new_n652), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT35), .ZN(new_n987));
  OAI211_X1 g0787(.A(G116), .B(new_n218), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(new_n987), .B2(new_n986), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT36), .Z(new_n990));
  AOI211_X1 g0790(.A(new_n219), .B(new_n230), .C1(G58), .C2(G68), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n257), .A2(G50), .ZN(new_n992));
  OAI211_X1 g0792(.A(G1), .B(new_n829), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT101), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n985), .A2(new_n995), .ZN(G367));
  INV_X1    g0796(.A(new_n738), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n665), .A2(new_n723), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n669), .A2(new_n998), .B1(new_n668), .B2(new_n724), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT108), .ZN(new_n1000));
  OAI21_X1  g0800(.A(KEYINPUT107), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT107), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1000), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n738), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  OR3_X1    g0805(.A1(new_n1000), .A2(KEYINPUT42), .A3(new_n740), .ZN(new_n1006));
  OAI21_X1  g0806(.A(KEYINPUT42), .B1(new_n1000), .B2(new_n740), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n694), .B1(new_n1003), .B2(new_n734), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1006), .B(new_n1007), .C1(new_n1008), .C2(new_n723), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n706), .A2(new_n723), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT105), .Z(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n712), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n689), .B2(new_n1011), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(KEYINPUT43), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1009), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1005), .A2(new_n1015), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1013), .A2(KEYINPUT106), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT43), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1013), .A2(KEYINPUT106), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1001), .A2(new_n1014), .A3(new_n1009), .A4(new_n1004), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1016), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1016), .A2(new_n1022), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n1020), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n745), .B(KEYINPUT41), .Z(new_n1026));
  NOR2_X1   g0826(.A1(new_n1000), .A2(new_n742), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT45), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1000), .A2(new_n742), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT44), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n738), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT109), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n855), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n732), .A2(KEYINPUT109), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n736), .A2(new_n739), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1035), .A2(new_n740), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n740), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1039), .A2(new_n1034), .A3(new_n855), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1028), .A2(new_n997), .A3(new_n1031), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1033), .A2(new_n1041), .A3(new_n779), .A4(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1026), .B1(new_n1043), .B2(new_n779), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n831), .A2(G1), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1023), .B(new_n1025), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n837), .B1(new_n210), .B2(new_n342), .C1(new_n246), .C2(new_n846), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n833), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n788), .A2(G50), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n790), .A2(G150), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n326), .B1(new_n816), .B2(new_n222), .C1(new_n807), .C2(new_n230), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G143), .B2(new_n809), .ZN(new_n1052));
  INV_X1    g0852(.A(G137), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n1053), .A2(new_n796), .B1(new_n801), .B2(new_n797), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G68), .B2(new_n823), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n788), .A2(G283), .ZN(new_n1057));
  AND3_X1   g0857(.A1(new_n804), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1058));
  AOI21_X1  g0858(.A(KEYINPUT46), .B1(new_n804), .B2(G116), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n1058), .A2(new_n1059), .A3(new_n326), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G294), .A2(new_n874), .B1(new_n882), .B2(G317), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n807), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1062), .A2(G97), .B1(new_n823), .B2(G107), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1057), .A2(new_n1060), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G303), .A2(new_n790), .B1(new_n809), .B2(G311), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT110), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1056), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT47), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1048), .B1(new_n1068), .B2(new_n781), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1013), .A2(new_n853), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1046), .A2(new_n1071), .ZN(G387));
  INV_X1    g0872(.A(new_n745), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n1041), .B2(new_n779), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n779), .B2(new_n1041), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n737), .A2(new_n836), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n845), .B1(new_n243), .B2(new_n847), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n747), .B2(new_n839), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n350), .A2(G50), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT50), .ZN(new_n1080));
  AOI21_X1  g0880(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1080), .A2(new_n747), .A3(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1078), .A2(new_n1082), .B1(new_n206), .B2(new_n744), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n833), .B1(new_n1083), .B2(new_n838), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n329), .B1(new_n804), .B2(new_n231), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n205), .B2(new_n807), .C1(new_n877), .C2(new_n202), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n809), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1087), .A2(new_n797), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(G150), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n1090), .A2(new_n796), .B1(new_n801), .B2(new_n409), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n802), .A2(new_n342), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1089), .B(new_n1093), .C1(new_n257), .C2(new_n787), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n326), .B1(new_n882), .B2(G326), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n804), .A2(G294), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n802), .B2(new_n820), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n790), .A2(G317), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n809), .A2(G322), .B1(new_n874), .B2(G311), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(new_n787), .C2(new_n489), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT48), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1097), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n1101), .B2(new_n1100), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT49), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1095), .B1(new_n501), .B2(new_n807), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1094), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1084), .B1(new_n1107), .B2(new_n781), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1041), .A2(new_n1045), .B1(new_n1076), .B2(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1075), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(G393));
  NOR2_X1   g0911(.A1(new_n251), .A2(new_n846), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n837), .B1(new_n205), .B2(new_n210), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G150), .A2(new_n809), .B1(new_n790), .B2(G159), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT112), .ZN(new_n1115));
  OR2_X1    g0915(.A1(new_n1115), .A2(KEYINPUT51), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(KEYINPUT51), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n787), .A2(new_n350), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n326), .B1(new_n816), .B2(new_n257), .C1(new_n807), .C2(new_n887), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n874), .A2(G50), .B1(new_n823), .B2(G77), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n876), .B2(new_n796), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1118), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1116), .A2(new_n1117), .A3(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(G311), .A2(new_n790), .B1(new_n809), .B2(G317), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n1124), .B(KEYINPUT52), .Z(new_n1125));
  AOI22_X1  g0925(.A1(new_n874), .A2(G303), .B1(new_n823), .B2(G116), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1126), .B(new_n329), .C1(new_n206), .C2(new_n807), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n788), .B2(G294), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n882), .A2(G322), .B1(G283), .B2(new_n804), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT113), .Z(new_n1130));
  NAND3_X1  g0930(.A1(new_n1125), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1123), .A2(new_n1131), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n833), .B1(new_n1112), .B2(new_n1113), .C1(new_n1132), .C2(new_n873), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n836), .B2(new_n1000), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1033), .A2(KEYINPUT111), .A3(new_n1042), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT111), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1032), .A2(new_n1136), .A3(new_n738), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1134), .B1(new_n1138), .B2(new_n1045), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1041), .A2(new_n779), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1135), .A2(new_n1140), .A3(new_n1137), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT114), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1043), .A2(new_n745), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1144), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT114), .B1(new_n1146), .B2(new_n1141), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1139), .B1(new_n1145), .B2(new_n1147), .ZN(G390));
  INV_X1    g0948(.A(new_n944), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n865), .A2(G330), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1149), .B1(new_n762), .B2(new_n1150), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n729), .B(new_n866), .C1(new_n760), .C2(new_n761), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1151), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n723), .B1(new_n771), .B2(new_n773), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n939), .B1(new_n1154), .B2(new_n865), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n762), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n1152), .B2(new_n1149), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n940), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1153), .A2(new_n1155), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n480), .A2(new_n762), .A3(G330), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(KEYINPUT115), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT115), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n480), .A2(new_n762), .A3(new_n1162), .A4(G330), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1164), .A2(new_n955), .A3(new_n683), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1159), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n962), .A2(new_n901), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1155), .B2(new_n944), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n900), .B1(new_n940), .B2(new_n944), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n916), .A2(new_n928), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(KEYINPUT104), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1169), .A2(new_n1171), .A3(new_n934), .A4(new_n929), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1152), .A2(new_n1149), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1168), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1166), .B(new_n1174), .C1(new_n1175), .C2(new_n1156), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1164), .A2(new_n683), .A3(new_n955), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1151), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1155), .A2(new_n1173), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1177), .A2(new_n1181), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1168), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1156), .B1(new_n1168), .B2(new_n1172), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1176), .A2(new_n1185), .A3(new_n745), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n1045), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT54), .B(G143), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n788), .A2(new_n1190), .B1(G137), .B2(new_n874), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1191), .A2(KEYINPUT116), .B1(G159), .B2(new_n823), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(KEYINPUT116), .B2(new_n1191), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT117), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n804), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT53), .B1(new_n804), .B2(G150), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1197), .A2(new_n329), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n882), .A2(G125), .B1(new_n1062), .B2(G50), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G128), .A2(new_n809), .B1(new_n790), .B2(G132), .ZN(new_n1200));
  AND4_X1   g1000(.A1(new_n1194), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n882), .A2(G294), .B1(new_n823), .B2(G77), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n880), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1202), .A2(new_n329), .A3(new_n805), .A4(new_n1203), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n809), .A2(G283), .B1(new_n874), .B2(G107), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n787), .B2(new_n205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT118), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1204), .B(new_n1207), .C1(G116), .C2(new_n790), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n781), .B1(new_n1201), .B2(new_n1208), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1171), .A2(new_n834), .A3(new_n934), .A4(new_n929), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n832), .B1(new_n409), .B2(new_n894), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1186), .A2(new_n1188), .A3(new_n1212), .ZN(G378));
  INV_X1    g1013(.A(new_n407), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n393), .A2(new_n903), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT121), .Z(new_n1218));
  NAND2_X1  g1018(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1216), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1218), .B1(new_n1216), .B2(new_n1219), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n979), .B2(G330), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n978), .B(new_n963), .C1(new_n761), .C2(new_n760), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n916), .A2(new_n950), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n973), .B1(new_n947), .B2(new_n951), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1227), .B(G330), .C1(new_n1228), .C2(KEYINPUT40), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(new_n1222), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n954), .B1(new_n1224), .B2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n979), .A2(G330), .A3(new_n1223), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1229), .A2(new_n1222), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1232), .A2(new_n937), .A3(new_n1233), .A4(new_n953), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G97), .A2(new_n874), .B1(new_n882), .B2(G283), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n329), .A2(new_n296), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n231), .B2(new_n804), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT119), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1236), .B(new_n1239), .C1(new_n787), .C2(new_n342), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n877), .A2(new_n206), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1062), .A2(G58), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1242), .B1(new_n257), .B2(new_n802), .C1(new_n1087), .C2(new_n501), .ZN(new_n1243));
  OR3_X1    g1043(.A1(new_n1240), .A2(new_n1241), .A3(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT58), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1237), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n823), .A2(G150), .B1(new_n804), .B2(new_n1190), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G132), .B2(new_n874), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(G125), .A2(new_n809), .B1(new_n790), .B2(G128), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1251), .B(new_n1252), .C1(new_n787), .C2(new_n1053), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1253), .A2(KEYINPUT59), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(KEYINPUT59), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n288), .B(new_n296), .C1(new_n807), .C2(new_n797), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(G124), .B2(new_n882), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n1248), .B1(new_n1245), .B2(new_n1244), .C1(new_n1254), .C2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n781), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT120), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1260), .B(new_n1261), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n832), .B(new_n1262), .C1(new_n202), .C2(new_n894), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1222), .A2(new_n834), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n1235), .A2(new_n1045), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1235), .A2(KEYINPUT57), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1165), .B1(new_n1187), .B2(new_n1181), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n745), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT57), .B1(new_n1269), .B2(new_n1235), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1265), .B1(new_n1268), .B2(new_n1270), .ZN(G375));
  NAND2_X1  g1071(.A1(new_n944), .A2(new_n834), .ZN(new_n1272));
  XOR2_X1   g1072(.A(new_n1272), .B(KEYINPUT122), .Z(new_n1273));
  NOR2_X1   g1073(.A1(new_n877), .A2(new_n820), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1092), .B1(G97), .B2(new_n804), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n1275), .B1(new_n501), .B2(new_n801), .C1(new_n489), .C2(new_n796), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n1274), .B(new_n1276), .C1(G294), .C2(new_n809), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n329), .B1(new_n807), .B2(new_n260), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(KEYINPUT123), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n787), .B2(new_n206), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n809), .A2(G132), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n790), .A2(G137), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n329), .B1(new_n804), .B2(G159), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1282), .A2(new_n1283), .A3(new_n1242), .A4(new_n1284), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(G128), .A2(new_n882), .B1(new_n874), .B2(new_n1190), .ZN(new_n1286));
  OAI221_X1 g1086(.A(new_n1286), .B1(new_n202), .B2(new_n802), .C1(new_n787), .C2(new_n1090), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n1278), .A2(new_n1281), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n781), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n832), .B1(new_n257), .B2(new_n894), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1273), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1045), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1291), .B1(new_n1159), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1026), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1182), .A2(new_n1295), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1177), .A2(new_n1181), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1294), .B1(new_n1296), .B2(new_n1297), .ZN(G381));
  INV_X1    g1098(.A(G396), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1110), .A2(new_n1299), .A3(new_n897), .ZN(new_n1300));
  OR3_X1    g1100(.A1(G387), .A2(G381), .A3(new_n1300), .ZN(new_n1301));
  OR4_X1    g1101(.A1(G390), .A2(new_n1301), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1102(.A(G378), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n722), .A2(G213), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  OAI211_X1 g1106(.A(G407), .B(G213), .C1(G375), .C2(new_n1306), .ZN(G409));
  AND2_X1   g1107(.A1(new_n1046), .A2(new_n1071), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(G390), .A2(new_n1308), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1110), .B(G396), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1143), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1146), .A2(KEYINPUT114), .A3(new_n1141), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1313), .A2(G387), .A3(new_n1139), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1309), .A2(new_n1310), .A3(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1310), .B1(new_n1309), .B2(new_n1314), .ZN(new_n1316));
  NOR3_X1   g1116(.A1(new_n1315), .A2(new_n1316), .A3(KEYINPUT61), .ZN(new_n1317));
  NOR3_X1   g1117(.A1(new_n1224), .A2(new_n1230), .A3(new_n954), .ZN(new_n1318));
  AOI22_X1  g1118(.A1(new_n1232), .A2(new_n1233), .B1(new_n937), .B2(new_n953), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1295), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(KEYINPUT124), .B1(new_n1320), .B2(new_n1267), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT124), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1269), .A2(new_n1322), .A3(new_n1295), .A4(new_n1235), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1321), .A2(new_n1265), .A3(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1303), .ZN(new_n1325));
  OAI211_X1 g1125(.A(G378), .B(new_n1265), .C1(new_n1268), .C2(new_n1270), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1305), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT60), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1328), .B1(new_n1177), .B2(new_n1181), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1073), .B1(new_n1177), .B2(new_n1181), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1159), .A2(KEYINPUT60), .A3(new_n1165), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1329), .A2(new_n1330), .A3(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(KEYINPUT125), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT125), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1329), .A2(new_n1330), .A3(new_n1334), .A4(new_n1331), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1333), .A2(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(G384), .B1(new_n1336), .B2(new_n1294), .ZN(new_n1337));
  AOI211_X1 g1137(.A(new_n897), .B(new_n1293), .C1(new_n1333), .C2(new_n1335), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1327), .A2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT63), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1305), .A2(G2897), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1343), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1344), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n745), .B1(new_n1159), .B2(new_n1165), .ZN(new_n1346));
  AOI21_X1  g1146(.A(KEYINPUT60), .B1(new_n1159), .B2(new_n1165), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1334), .B1(new_n1348), .B2(new_n1331), .ZN(new_n1349));
  AND4_X1   g1149(.A1(new_n1334), .A2(new_n1329), .A3(new_n1330), .A4(new_n1331), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1294), .B1(new_n1349), .B2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(new_n897), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1336), .A2(G384), .A3(new_n1294), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1352), .A2(new_n1353), .A3(new_n1343), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1345), .A2(new_n1354), .ZN(new_n1355));
  OR2_X1    g1155(.A1(new_n1327), .A2(new_n1355), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1327), .A2(KEYINPUT63), .A3(new_n1339), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1317), .A2(new_n1342), .A3(new_n1356), .A4(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT62), .ZN(new_n1359));
  AND3_X1   g1159(.A1(new_n1327), .A2(new_n1359), .A3(new_n1339), .ZN(new_n1360));
  XOR2_X1   g1160(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1361));
  OAI21_X1  g1161(.A(new_n1361), .B1(new_n1327), .B2(new_n1355), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1359), .B1(new_n1327), .B2(new_n1339), .ZN(new_n1363));
  NOR3_X1   g1163(.A1(new_n1360), .A2(new_n1362), .A3(new_n1363), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1358), .B1(new_n1364), .B2(new_n1365), .ZN(G405));
  NAND2_X1  g1166(.A1(G375), .A2(new_n1303), .ZN(new_n1367));
  OAI21_X1  g1167(.A(new_n1367), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1326), .A2(KEYINPUT127), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1339), .A2(new_n1303), .A3(G375), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1368), .A2(new_n1369), .A3(new_n1370), .ZN(new_n1371));
  INV_X1    g1171(.A(new_n1371), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1369), .B1(new_n1368), .B2(new_n1370), .ZN(new_n1373));
  OAI22_X1  g1173(.A1(new_n1372), .A2(new_n1373), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1374));
  INV_X1    g1174(.A(new_n1373), .ZN(new_n1375));
  NAND3_X1  g1175(.A1(new_n1375), .A2(new_n1365), .A3(new_n1371), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1374), .A2(new_n1376), .ZN(G402));
endmodule


