

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582;

  INV_X1 U323 ( .A(KEYINPUT92), .ZN(n328) );
  XNOR2_X1 U324 ( .A(n433), .B(n432), .ZN(n434) );
  AND2_X1 U325 ( .A1(G229GAT), .A2(G233GAT), .ZN(n291) );
  XOR2_X1 U326 ( .A(n381), .B(n380), .Z(n520) );
  XNOR2_X1 U327 ( .A(KEYINPUT113), .B(KEYINPUT46), .ZN(n453) );
  XNOR2_X1 U328 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U329 ( .A(KEYINPUT27), .B(KEYINPUT94), .ZN(n342) );
  XNOR2_X1 U330 ( .A(n517), .B(n342), .ZN(n385) );
  XOR2_X1 U331 ( .A(G8GAT), .B(G183GAT), .Z(n325) );
  XNOR2_X1 U332 ( .A(n424), .B(n291), .ZN(n425) );
  XNOR2_X1 U333 ( .A(n426), .B(n425), .ZN(n428) );
  XNOR2_X1 U334 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U335 ( .A(KEYINPUT55), .B(KEYINPUT123), .ZN(n470) );
  XNOR2_X1 U336 ( .A(n331), .B(n330), .ZN(n335) );
  XNOR2_X1 U337 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U338 ( .A(n435), .B(n434), .ZN(n452) );
  XOR2_X1 U339 ( .A(n469), .B(KEYINPUT28), .Z(n530) );
  XNOR2_X1 U340 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U341 ( .A(G36GAT), .B(KEYINPUT104), .ZN(n450) );
  XNOR2_X1 U342 ( .A(n476), .B(n475), .ZN(G1349GAT) );
  XNOR2_X1 U343 ( .A(n451), .B(n450), .ZN(G1329GAT) );
  XNOR2_X1 U344 ( .A(KEYINPUT37), .B(KEYINPUT102), .ZN(n417) );
  XOR2_X1 U345 ( .A(G78GAT), .B(G155GAT), .Z(n293) );
  XNOR2_X1 U346 ( .A(G127GAT), .B(G71GAT), .ZN(n292) );
  XNOR2_X1 U347 ( .A(n293), .B(n292), .ZN(n306) );
  XOR2_X1 U348 ( .A(G57GAT), .B(KEYINPUT13), .Z(n443) );
  XOR2_X1 U349 ( .A(n443), .B(n325), .Z(n295) );
  NAND2_X1 U350 ( .A1(G231GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U351 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U352 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n297) );
  XNOR2_X1 U353 ( .A(KEYINPUT15), .B(KEYINPUT74), .ZN(n296) );
  XNOR2_X1 U354 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U355 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U356 ( .A(G15GAT), .B(G22GAT), .Z(n418) );
  XOR2_X1 U357 ( .A(KEYINPUT12), .B(G64GAT), .Z(n301) );
  XNOR2_X1 U358 ( .A(G1GAT), .B(G211GAT), .ZN(n300) );
  XNOR2_X1 U359 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n418), .B(n302), .ZN(n303) );
  XNOR2_X1 U361 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U362 ( .A(n306), .B(n305), .Z(n459) );
  XNOR2_X1 U363 ( .A(KEYINPUT87), .B(KEYINPUT86), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n307), .B(KEYINPUT3), .ZN(n308) );
  XOR2_X1 U365 ( .A(n308), .B(KEYINPUT2), .Z(n310) );
  XNOR2_X1 U366 ( .A(G141GAT), .B(G155GAT), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n310), .B(n309), .ZN(n358) );
  XOR2_X1 U368 ( .A(KEYINPUT85), .B(G218GAT), .Z(n312) );
  XNOR2_X1 U369 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n311) );
  XNOR2_X1 U370 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U371 ( .A(G197GAT), .B(n313), .Z(n339) );
  XNOR2_X1 U372 ( .A(n358), .B(n339), .ZN(n324) );
  XOR2_X1 U373 ( .A(G50GAT), .B(G162GAT), .Z(n406) );
  XOR2_X1 U374 ( .A(KEYINPUT84), .B(KEYINPUT24), .Z(n315) );
  XNOR2_X1 U375 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U377 ( .A(n406), .B(n316), .Z(n318) );
  NAND2_X1 U378 ( .A1(G228GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U380 ( .A(n319), .B(KEYINPUT22), .Z(n322) );
  XNOR2_X1 U381 ( .A(G106GAT), .B(G78GAT), .ZN(n320) );
  XNOR2_X1 U382 ( .A(n320), .B(G148GAT), .ZN(n440) );
  XNOR2_X1 U383 ( .A(n440), .B(G204GAT), .ZN(n321) );
  XNOR2_X1 U384 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U385 ( .A(n324), .B(n323), .ZN(n469) );
  XOR2_X1 U386 ( .A(n325), .B(KEYINPUT93), .Z(n327) );
  NAND2_X1 U387 ( .A1(G226GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U388 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U389 ( .A(G36GAT), .B(G190GAT), .Z(n405) );
  XNOR2_X1 U390 ( .A(n405), .B(KEYINPUT91), .ZN(n329) );
  XOR2_X1 U391 ( .A(G92GAT), .B(G64GAT), .Z(n333) );
  XNOR2_X1 U392 ( .A(G176GAT), .B(KEYINPUT71), .ZN(n332) );
  XNOR2_X1 U393 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U394 ( .A(G204GAT), .B(n334), .Z(n445) );
  XNOR2_X1 U395 ( .A(n335), .B(n445), .ZN(n341) );
  XOR2_X1 U396 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n337) );
  XNOR2_X1 U397 ( .A(KEYINPUT17), .B(KEYINPUT82), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U399 ( .A(G169GAT), .B(n338), .Z(n377) );
  XOR2_X1 U400 ( .A(n377), .B(n339), .Z(n340) );
  XOR2_X1 U401 ( .A(n341), .B(n340), .Z(n517) );
  XOR2_X1 U402 ( .A(KEYINPUT78), .B(G134GAT), .Z(n344) );
  XNOR2_X1 U403 ( .A(KEYINPUT77), .B(G127GAT), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U405 ( .A(KEYINPUT0), .B(n345), .Z(n381) );
  XOR2_X1 U406 ( .A(KEYINPUT1), .B(G162GAT), .Z(n347) );
  XNOR2_X1 U407 ( .A(G120GAT), .B(G148GAT), .ZN(n346) );
  XNOR2_X1 U408 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U409 ( .A(n348), .B(G85GAT), .Z(n350) );
  XOR2_X1 U410 ( .A(G113GAT), .B(G1GAT), .Z(n419) );
  XNOR2_X1 U411 ( .A(G29GAT), .B(n419), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U413 ( .A(n381), .B(n351), .ZN(n362) );
  XOR2_X1 U414 ( .A(KEYINPUT90), .B(KEYINPUT5), .Z(n353) );
  XNOR2_X1 U415 ( .A(KEYINPUT4), .B(G57GAT), .ZN(n352) );
  XNOR2_X1 U416 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U417 ( .A(KEYINPUT89), .B(n354), .Z(n356) );
  NAND2_X1 U418 ( .A1(G225GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U419 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U420 ( .A(n357), .B(KEYINPUT88), .Z(n360) );
  XNOR2_X1 U421 ( .A(n358), .B(KEYINPUT6), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n362), .B(n361), .ZN(n514) );
  NAND2_X1 U424 ( .A1(n385), .A2(n514), .ZN(n363) );
  XOR2_X1 U425 ( .A(KEYINPUT95), .B(n363), .Z(n527) );
  NOR2_X1 U426 ( .A1(n530), .A2(n527), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n364), .B(KEYINPUT96), .ZN(n382) );
  XOR2_X1 U428 ( .A(KEYINPUT79), .B(G176GAT), .Z(n366) );
  XNOR2_X1 U429 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U431 ( .A(KEYINPUT81), .B(KEYINPUT83), .Z(n368) );
  XNOR2_X1 U432 ( .A(G113GAT), .B(G183GAT), .ZN(n367) );
  XNOR2_X1 U433 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U434 ( .A(n370), .B(n369), .Z(n379) );
  XOR2_X1 U435 ( .A(G120GAT), .B(G71GAT), .Z(n446) );
  XOR2_X1 U436 ( .A(KEYINPUT80), .B(G190GAT), .Z(n372) );
  XNOR2_X1 U437 ( .A(G43GAT), .B(G99GAT), .ZN(n371) );
  XNOR2_X1 U438 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U439 ( .A(n446), .B(n373), .Z(n375) );
  NAND2_X1 U440 ( .A1(G227GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U441 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U442 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n379), .B(n378), .ZN(n380) );
  AND2_X1 U444 ( .A1(n382), .A2(n531), .ZN(n394) );
  NOR2_X1 U445 ( .A1(n520), .A2(n469), .ZN(n383) );
  XOR2_X1 U446 ( .A(KEYINPUT97), .B(n383), .Z(n384) );
  XNOR2_X1 U447 ( .A(KEYINPUT26), .B(n384), .ZN(n565) );
  NAND2_X1 U448 ( .A1(n385), .A2(n565), .ZN(n386) );
  XOR2_X1 U449 ( .A(KEYINPUT98), .B(n386), .Z(n391) );
  NAND2_X1 U450 ( .A1(n517), .A2(n520), .ZN(n387) );
  NAND2_X1 U451 ( .A1(n387), .A2(n469), .ZN(n388) );
  XNOR2_X1 U452 ( .A(n388), .B(KEYINPUT99), .ZN(n389) );
  XOR2_X1 U453 ( .A(KEYINPUT25), .B(n389), .Z(n390) );
  NOR2_X1 U454 ( .A1(n391), .A2(n390), .ZN(n392) );
  NOR2_X1 U455 ( .A1(n514), .A2(n392), .ZN(n393) );
  NOR2_X1 U456 ( .A1(n394), .A2(n393), .ZN(n481) );
  XOR2_X1 U457 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n396) );
  XNOR2_X1 U458 ( .A(KEYINPUT65), .B(KEYINPUT10), .ZN(n395) );
  XNOR2_X1 U459 ( .A(n396), .B(n395), .ZN(n414) );
  XOR2_X1 U460 ( .A(KEYINPUT9), .B(KEYINPUT64), .Z(n398) );
  NAND2_X1 U461 ( .A1(G232GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U462 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U463 ( .A(n399), .B(KEYINPUT73), .Z(n404) );
  XOR2_X1 U464 ( .A(G29GAT), .B(G43GAT), .Z(n401) );
  XNOR2_X1 U465 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n401), .B(n400), .ZN(n429) );
  XNOR2_X1 U467 ( .A(G99GAT), .B(G85GAT), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n402), .B(KEYINPUT70), .ZN(n439) );
  XNOR2_X1 U469 ( .A(n429), .B(n439), .ZN(n403) );
  XNOR2_X1 U470 ( .A(n404), .B(n403), .ZN(n410) );
  XOR2_X1 U471 ( .A(n405), .B(G92GAT), .Z(n408) );
  XNOR2_X1 U472 ( .A(G106GAT), .B(n406), .ZN(n407) );
  XNOR2_X1 U473 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U474 ( .A(n410), .B(n409), .Z(n412) );
  XNOR2_X1 U475 ( .A(G134GAT), .B(G218GAT), .ZN(n411) );
  XNOR2_X1 U476 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U477 ( .A(n414), .B(n413), .ZN(n561) );
  XOR2_X1 U478 ( .A(KEYINPUT36), .B(n561), .Z(n580) );
  NOR2_X1 U479 ( .A1(n481), .A2(n580), .ZN(n415) );
  NAND2_X1 U480 ( .A1(n459), .A2(n415), .ZN(n416) );
  XNOR2_X1 U481 ( .A(n417), .B(n416), .ZN(n511) );
  XOR2_X1 U482 ( .A(G36GAT), .B(G50GAT), .Z(n421) );
  XNOR2_X1 U483 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n426) );
  XOR2_X1 U485 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n423) );
  XNOR2_X1 U486 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n424) );
  INV_X1 U488 ( .A(KEYINPUT66), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n428), .B(n427), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n429), .B(KEYINPUT67), .ZN(n433) );
  XOR2_X1 U491 ( .A(G8GAT), .B(G197GAT), .Z(n431) );
  XNOR2_X1 U492 ( .A(G169GAT), .B(G141GAT), .ZN(n430) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n432) );
  INV_X1 U494 ( .A(n452), .ZN(n558) );
  XOR2_X1 U495 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n437) );
  NAND2_X1 U496 ( .A1(G230GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U498 ( .A(n438), .B(KEYINPUT31), .Z(n442) );
  XNOR2_X1 U499 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U502 ( .A(n446), .B(n445), .Z(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n570) );
  NOR2_X1 U504 ( .A1(n452), .A2(n570), .ZN(n482) );
  NAND2_X1 U505 ( .A1(n511), .A2(n482), .ZN(n449) );
  XOR2_X1 U506 ( .A(KEYINPUT38), .B(n449), .Z(n497) );
  NAND2_X1 U507 ( .A1(n497), .A2(n517), .ZN(n451) );
  INV_X1 U508 ( .A(n520), .ZN(n531) );
  INV_X1 U509 ( .A(n517), .ZN(n466) );
  INV_X1 U510 ( .A(n459), .ZN(n573) );
  XOR2_X1 U511 ( .A(n570), .B(KEYINPUT41), .Z(n550) );
  NAND2_X1 U512 ( .A1(n558), .A2(n550), .ZN(n454) );
  NOR2_X1 U513 ( .A1(n573), .A2(n455), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n456), .B(KEYINPUT114), .ZN(n457) );
  INV_X1 U515 ( .A(n561), .ZN(n477) );
  NAND2_X1 U516 ( .A1(n457), .A2(n477), .ZN(n458) );
  XNOR2_X1 U517 ( .A(n458), .B(KEYINPUT47), .ZN(n464) );
  NOR2_X1 U518 ( .A1(n459), .A2(n580), .ZN(n460) );
  XNOR2_X1 U519 ( .A(n460), .B(KEYINPUT45), .ZN(n461) );
  NAND2_X1 U520 ( .A1(n461), .A2(n452), .ZN(n462) );
  NOR2_X1 U521 ( .A1(n462), .A2(n570), .ZN(n463) );
  NOR2_X1 U522 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n465), .B(KEYINPUT48), .ZN(n528) );
  NOR2_X1 U524 ( .A1(n466), .A2(n528), .ZN(n467) );
  XOR2_X1 U525 ( .A(KEYINPUT54), .B(n467), .Z(n468) );
  NOR2_X1 U526 ( .A1(n514), .A2(n468), .ZN(n566) );
  NAND2_X1 U527 ( .A1(n566), .A2(n469), .ZN(n471) );
  NOR2_X1 U528 ( .A1(n531), .A2(n472), .ZN(n562) );
  XNOR2_X1 U529 ( .A(n550), .B(KEYINPUT106), .ZN(n536) );
  NAND2_X1 U530 ( .A1(n562), .A2(n536), .ZN(n476) );
  XOR2_X1 U531 ( .A(G176GAT), .B(KEYINPUT124), .Z(n474) );
  XNOR2_X1 U532 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n473) );
  NAND2_X1 U533 ( .A1(n573), .A2(n477), .ZN(n478) );
  XNOR2_X1 U534 ( .A(n478), .B(KEYINPUT76), .ZN(n479) );
  XNOR2_X1 U535 ( .A(n479), .B(KEYINPUT16), .ZN(n480) );
  NOR2_X1 U536 ( .A1(n481), .A2(n480), .ZN(n500) );
  AND2_X1 U537 ( .A1(n482), .A2(n500), .ZN(n490) );
  NAND2_X1 U538 ( .A1(n490), .A2(n514), .ZN(n483) );
  XNOR2_X1 U539 ( .A(n483), .B(KEYINPUT34), .ZN(n484) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(n484), .ZN(G1324GAT) );
  NAND2_X1 U541 ( .A1(n517), .A2(n490), .ZN(n485) );
  XNOR2_X1 U542 ( .A(n485), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n487) );
  NAND2_X1 U544 ( .A1(n490), .A2(n520), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(n489) );
  XOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT100), .Z(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(G1326GAT) );
  NAND2_X1 U548 ( .A1(n490), .A2(n530), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n491), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U550 ( .A1(n497), .A2(n514), .ZN(n494) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n492), .B(KEYINPUT103), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U554 ( .A1(n497), .A2(n520), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n495), .B(KEYINPUT40), .ZN(n496) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n496), .ZN(G1330GAT) );
  XOR2_X1 U557 ( .A(G50GAT), .B(KEYINPUT105), .Z(n499) );
  NAND2_X1 U558 ( .A1(n530), .A2(n497), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(G1331GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n503) );
  NAND2_X1 U561 ( .A1(n452), .A2(n536), .ZN(n512) );
  INV_X1 U562 ( .A(n500), .ZN(n501) );
  NOR2_X1 U563 ( .A1(n512), .A2(n501), .ZN(n508) );
  NAND2_X1 U564 ( .A1(n508), .A2(n514), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(n504), .ZN(G1332GAT) );
  NAND2_X1 U567 ( .A1(n517), .A2(n508), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n505), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U569 ( .A1(n508), .A2(n520), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(KEYINPUT108), .ZN(n507) );
  XNOR2_X1 U571 ( .A(G71GAT), .B(n507), .ZN(G1334GAT) );
  XOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U573 ( .A1(n508), .A2(n530), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  XOR2_X1 U575 ( .A(G85GAT), .B(KEYINPUT109), .Z(n516) );
  INV_X1 U576 ( .A(n511), .ZN(n513) );
  NOR2_X1 U577 ( .A1(n513), .A2(n512), .ZN(n522) );
  NAND2_X1 U578 ( .A1(n522), .A2(n514), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n517), .A2(n522), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n518), .B(KEYINPUT110), .ZN(n519) );
  XNOR2_X1 U582 ( .A(G92GAT), .B(n519), .ZN(G1337GAT) );
  NAND2_X1 U583 ( .A1(n522), .A2(n520), .ZN(n521) );
  XNOR2_X1 U584 ( .A(n521), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n526) );
  XOR2_X1 U586 ( .A(KEYINPUT112), .B(KEYINPUT111), .Z(n524) );
  NAND2_X1 U587 ( .A1(n522), .A2(n530), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n526), .B(n525), .ZN(G1339GAT) );
  NOR2_X1 U590 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U591 ( .A(n529), .B(KEYINPUT115), .Z(n546) );
  NOR2_X1 U592 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U593 ( .A1(n546), .A2(n532), .ZN(n533) );
  XOR2_X1 U594 ( .A(KEYINPUT116), .B(n533), .Z(n542) );
  AND2_X1 U595 ( .A1(n542), .A2(n558), .ZN(n535) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(KEYINPUT117), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n535), .B(n534), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n538) );
  NAND2_X1 U599 ( .A1(n542), .A2(n536), .ZN(n537) );
  XNOR2_X1 U600 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n540) );
  NAND2_X1 U602 ( .A1(n542), .A2(n573), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U604 ( .A(G127GAT), .B(n541), .Z(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U606 ( .A1(n542), .A2(n561), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U608 ( .A(G134GAT), .B(n545), .Z(G1343GAT) );
  XOR2_X1 U609 ( .A(G141GAT), .B(KEYINPUT121), .Z(n549) );
  NAND2_X1 U610 ( .A1(n546), .A2(n565), .ZN(n547) );
  XOR2_X1 U611 ( .A(KEYINPUT120), .B(n547), .Z(n556) );
  NAND2_X1 U612 ( .A1(n558), .A2(n556), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n549), .B(n548), .ZN(G1344GAT) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n554) );
  XOR2_X1 U615 ( .A(KEYINPUT122), .B(KEYINPUT52), .Z(n552) );
  NAND2_X1 U616 ( .A1(n550), .A2(n556), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n556), .A2(n573), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n556), .A2(n561), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n557), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U623 ( .A1(n562), .A2(n558), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U625 ( .A1(n573), .A2(n562), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U627 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1351GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n579) );
  NOR2_X1 U631 ( .A1(n452), .A2(n579), .ZN(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n572) );
  INV_X1 U636 ( .A(n579), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n574), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  XOR2_X1 U639 ( .A(G211GAT), .B(KEYINPUT125), .Z(n576) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1354GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n578) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n582) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(n582), .B(n581), .Z(G1355GAT) );
endmodule

