//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n454), .A2(G567), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n457), .A2(KEYINPUT65), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(new_n453), .B2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(KEYINPUT65), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(KEYINPUT66), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n472), .A2(new_n475), .ZN(G160));
  INV_X1    g051(.A(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT3), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n468), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(G2105), .ZN(new_n483));
  AOI22_X1  g058(.A1(G124), .A2(new_n482), .B1(new_n483), .B2(G136), .ZN(new_n484));
  OR2_X1    g059(.A1(new_n468), .A2(G112), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n486), .B1(G100), .B2(G2105), .ZN(new_n487));
  OR3_X1    g062(.A1(new_n486), .A2(G100), .A3(G2105), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n485), .A2(G2104), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n470), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n478), .A2(new_n480), .A3(G126), .ZN(new_n495));
  NAND2_X1  g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n463), .A2(G102), .A3(G2104), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n492), .A2(new_n493), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n468), .A2(new_n469), .A3(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n494), .A2(new_n498), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XOR2_X1   g086(.A(KEYINPUT68), .B(G651), .Z(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g089(.A(new_n514), .B(KEYINPUT69), .Z(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n516), .A2(G543), .A3(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n509), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n516), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(G50), .A2(new_n520), .B1(new_n523), .B2(G88), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n515), .A2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  AND2_X1   g101(.A1(new_n520), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n522), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT70), .ZN(new_n532));
  XOR2_X1   g107(.A(new_n532), .B(KEYINPUT7), .Z(new_n533));
  NOR3_X1   g108(.A1(new_n527), .A2(new_n530), .A3(new_n533), .ZN(G168));
  XNOR2_X1  g109(.A(KEYINPUT71), .B(G90), .ZN(new_n535));
  AOI22_X1  g110(.A1(G52), .A2(new_n520), .B1(new_n523), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT72), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(new_n512), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND2_X1  g116(.A1(new_n523), .A2(G81), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n520), .A2(G43), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n512), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n509), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n523), .A2(G91), .B1(G651), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n519), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n520), .A2(KEYINPUT9), .A3(G53), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n557), .A2(new_n560), .A3(new_n561), .ZN(G299));
  INV_X1    g137(.A(G168), .ZN(G286));
  NAND2_X1  g138(.A1(new_n520), .A2(G49), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n523), .A2(G87), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(G288));
  NAND2_X1  g142(.A1(new_n523), .A2(G86), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n520), .A2(G48), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n521), .A2(KEYINPUT73), .A3(G61), .ZN(new_n570));
  NAND2_X1  g145(.A1(G73), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT73), .ZN(new_n572));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n509), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n570), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(new_n513), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n568), .A2(new_n569), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT74), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT74), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  AND2_X1   g156(.A1(new_n579), .A2(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n512), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n584), .B(KEYINPUT75), .Z(new_n585));
  AOI22_X1  g160(.A1(G47), .A2(new_n520), .B1(new_n523), .B2(G85), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n509), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n520), .A2(G54), .B1(G651), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(G92), .ZN(new_n592));
  OR3_X1    g167(.A1(new_n522), .A2(KEYINPUT10), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(KEYINPUT10), .B1(new_n522), .B2(new_n592), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(G171), .B2(new_n596), .ZN(G284));
  OAI21_X1  g173(.A(new_n597), .B1(G171), .B2(new_n596), .ZN(G321));
  NAND2_X1  g174(.A1(G299), .A2(new_n596), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(G168), .B2(new_n596), .ZN(G297));
  OAI21_X1  g176(.A(new_n600), .B1(G168), .B2(new_n596), .ZN(G280));
  INV_X1    g177(.A(new_n595), .ZN(new_n603));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G860), .ZN(G148));
  OAI21_X1  g180(.A(KEYINPUT76), .B1(new_n547), .B2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n603), .A2(new_n604), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  MUX2_X1   g183(.A(KEYINPUT76), .B(new_n606), .S(new_n608), .Z(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g185(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2100), .ZN(new_n614));
  AOI22_X1  g189(.A1(G123), .A2(new_n482), .B1(new_n483), .B2(G135), .ZN(new_n615));
  OAI221_X1 g190(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n468), .C2(G111), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G2096), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n614), .A2(new_n619), .ZN(G156));
  XOR2_X1   g195(.A(KEYINPUT15), .B(G2435), .Z(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT77), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2427), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT78), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n623), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(KEYINPUT14), .ZN(new_n627));
  XOR2_X1   g202(.A(G2451), .B(G2454), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n627), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT79), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT80), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(G14), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n638), .B1(new_n632), .B2(new_n634), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n635), .A2(new_n636), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n637), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  XNOR2_X1  g218(.A(G2072), .B(G2078), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2067), .B(G2678), .Z(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(KEYINPUT17), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n647), .B1(new_n649), .B2(new_n646), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT81), .Z(new_n651));
  INV_X1    g226(.A(new_n646), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n652), .A2(new_n644), .A3(new_n643), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT18), .Z(new_n654));
  NAND3_X1  g229(.A1(new_n649), .A2(new_n643), .A3(new_n646), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n651), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(new_n618), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(G2100), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G227));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT82), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT19), .Z(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT83), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n663), .A2(new_n664), .ZN(new_n669));
  AOI22_X1  g244(.A1(new_n667), .A2(new_n668), .B1(new_n662), .B2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n669), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(new_n665), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n662), .A2(new_n672), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n670), .B(new_n673), .C1(new_n668), .C2(new_n667), .ZN(new_n674));
  XOR2_X1   g249(.A(G1991), .B(G1996), .Z(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n674), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1981), .B(G1986), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT84), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT85), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(G229));
  INV_X1    g257(.A(KEYINPUT30), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(G28), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(G28), .ZN(new_n685));
  INV_X1    g260(.A(G29), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(new_n617), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(G164), .A2(G29), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G27), .B2(G29), .ZN(new_n690));
  INV_X1    g265(.A(G2078), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G20), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT98), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT23), .ZN(new_n696));
  INV_X1    g271(.A(G299), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n693), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1956), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n690), .A2(new_n691), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(G29), .A2(G32), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n482), .A2(G129), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n483), .A2(G141), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n705));
  NAND3_X1  g280(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT26), .Z(new_n707));
  NAND4_X1  g282(.A1(new_n703), .A2(new_n704), .A3(new_n705), .A4(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n702), .B1(new_n708), .B2(new_n686), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT27), .B(G1996), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT96), .ZN(new_n712));
  INV_X1    g287(.A(G34), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n713), .A2(KEYINPUT24), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(KEYINPUT24), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n686), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G160), .B2(new_n686), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G2084), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n712), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G2072), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n720), .A2(KEYINPUT95), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT93), .B(KEYINPUT25), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n483), .A2(G139), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n468), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT94), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G29), .ZN(new_n730));
  OR2_X1    g305(.A1(G29), .A2(G33), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n721), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n720), .A2(KEYINPUT95), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n730), .A2(KEYINPUT95), .A3(new_n720), .A4(new_n731), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n719), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT97), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI211_X1 g313(.A(KEYINPUT97), .B(new_n719), .C1(new_n734), .C2(new_n735), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n692), .B(new_n701), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n603), .A2(G16), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G4), .B2(G16), .ZN(new_n742));
  INV_X1    g317(.A(G1348), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n547), .A2(G16), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G16), .B2(G19), .ZN(new_n745));
  INV_X1    g320(.A(G1341), .ZN(new_n746));
  OAI22_X1  g321(.A1(new_n742), .A2(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT92), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n686), .A2(G26), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n749), .B(new_n750), .Z(new_n751));
  NAND2_X1  g326(.A1(new_n482), .A2(G128), .ZN(new_n752));
  OAI221_X1 g327(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n468), .C2(G116), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n483), .A2(G140), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n751), .B1(new_n686), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2067), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n693), .A2(G21), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G168), .B2(new_n693), .ZN(new_n760));
  INV_X1    g335(.A(G1966), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G2090), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n686), .A2(G35), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G162), .B2(new_n686), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT29), .Z(new_n766));
  OAI21_X1  g341(.A(new_n762), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  NOR4_X1   g342(.A1(new_n740), .A2(new_n747), .A3(new_n758), .A4(new_n767), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n709), .A2(new_n710), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n745), .B2(new_n746), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n693), .A2(G5), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G171), .B2(new_n693), .ZN(new_n773));
  INV_X1    g348(.A(G1961), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n742), .A2(new_n743), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n768), .A2(new_n771), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  OR2_X1    g352(.A1(G16), .A2(G23), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G288), .B2(new_n693), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT33), .B(G1976), .Z(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n779), .B(new_n781), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n693), .A2(G22), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G303), .B2(G16), .ZN(new_n784));
  INV_X1    g359(.A(G1971), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  OR3_X1    g362(.A1(new_n782), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT32), .B(G1981), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT88), .ZN(new_n790));
  NOR2_X1   g365(.A1(G6), .A2(G16), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n790), .B(new_n792), .C1(G305), .C2(new_n693), .ZN(new_n793));
  INV_X1    g368(.A(new_n790), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n693), .B1(new_n579), .B2(new_n581), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n791), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(KEYINPUT89), .B1(new_n788), .B2(new_n797), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n782), .A2(new_n786), .A3(new_n787), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT89), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n799), .A2(new_n800), .A3(new_n793), .A4(new_n796), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n798), .A2(new_n801), .A3(KEYINPUT34), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT90), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n798), .A2(new_n801), .A3(KEYINPUT90), .A4(KEYINPUT34), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI221_X1 g381(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n468), .C2(G107), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT86), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n482), .A2(G119), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n483), .A2(G131), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  MUX2_X1   g386(.A(G25), .B(new_n811), .S(G29), .Z(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT35), .B(G1991), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT87), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n812), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n798), .A2(new_n801), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n693), .A2(G24), .ZN(new_n819));
  INV_X1    g394(.A(G290), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(new_n693), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(G1986), .Z(new_n822));
  NAND4_X1  g397(.A1(new_n806), .A2(new_n815), .A3(new_n818), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT36), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n804), .A2(new_n805), .B1(new_n817), .B2(new_n816), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n825), .A2(new_n826), .A3(new_n815), .A4(new_n822), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n777), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n766), .A2(new_n763), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n717), .A2(G2084), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT31), .B(G11), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n828), .A2(new_n829), .A3(new_n830), .A4(new_n831), .ZN(G150));
  INV_X1    g407(.A(G150), .ZN(G311));
  NAND2_X1  g408(.A1(new_n523), .A2(G93), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n520), .A2(G55), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n834), .B(new_n835), .C1(new_n512), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G860), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT99), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT37), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n837), .B(new_n546), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n595), .A2(new_n604), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n840), .B1(new_n845), .B2(G860), .ZN(G145));
  XNOR2_X1  g421(.A(new_n490), .B(G160), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(new_n617), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n756), .B(new_n502), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n729), .B(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(new_n708), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n811), .B(new_n612), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n482), .A2(G130), .ZN(new_n853));
  OAI221_X1 g428(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n468), .C2(G118), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n483), .A2(G142), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n852), .B(new_n856), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT100), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n851), .A2(new_n858), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n857), .A2(KEYINPUT100), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n860), .A2(new_n858), .A3(new_n851), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n848), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n859), .A2(new_n848), .A3(new_n861), .ZN(new_n865));
  INV_X1    g440(.A(G37), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g444(.A1(new_n837), .A2(new_n596), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT106), .ZN(new_n871));
  INV_X1    g446(.A(G288), .ZN(new_n872));
  XNOR2_X1  g447(.A(G305), .B(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n820), .ZN(new_n874));
  XOR2_X1   g449(.A(G303), .B(KEYINPUT104), .Z(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n875), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n873), .A2(G290), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n873), .A2(G290), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT42), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n841), .B(new_n607), .Z(new_n883));
  NAND2_X1  g458(.A1(new_n603), .A2(G299), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n697), .A2(new_n595), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  OR3_X1    g462(.A1(new_n883), .A2(KEYINPUT102), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(KEYINPUT102), .B1(new_n883), .B2(new_n887), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(KEYINPUT41), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n697), .A2(KEYINPUT103), .A3(new_n595), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(new_n886), .B2(KEYINPUT103), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n890), .B1(new_n892), .B2(KEYINPUT41), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n883), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n888), .A2(new_n889), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n895), .A2(new_n896), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n882), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(G868), .B1(new_n882), .B2(new_n897), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n871), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n882), .A2(new_n897), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n882), .A2(new_n897), .A3(new_n898), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n902), .A2(KEYINPUT106), .A3(G868), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n901), .A2(new_n904), .ZN(G295));
  NAND2_X1  g480(.A1(new_n901), .A2(new_n904), .ZN(G331));
  NAND2_X1  g481(.A1(G301), .A2(G168), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n537), .A2(G286), .A3(new_n539), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n841), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n910), .A2(KEYINPUT107), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n841), .B1(new_n907), .B2(new_n908), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT107), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n886), .A3(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n910), .A2(new_n912), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n893), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n866), .B1(new_n881), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n914), .A2(new_n916), .A3(KEYINPUT108), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n881), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT43), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n911), .A2(new_n913), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n892), .A2(KEYINPUT41), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n926), .B(KEYINPUT109), .C1(KEYINPUT41), .C2(new_n887), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n925), .B(new_n927), .C1(KEYINPUT109), .C2(new_n926), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n915), .A2(new_n887), .ZN(new_n929));
  AOI22_X1  g504(.A1(new_n928), .A2(new_n929), .B1(new_n876), .B2(new_n880), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n930), .A2(new_n918), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT44), .B1(new_n924), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n919), .B2(new_n923), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n930), .A2(new_n918), .A3(KEYINPUT43), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n933), .B1(new_n936), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g512(.A(KEYINPUT125), .ZN(new_n938));
  INV_X1    g513(.A(G1384), .ZN(new_n939));
  INV_X1    g514(.A(new_n496), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n469), .B2(G126), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n499), .B(new_n501), .C1(new_n941), .C2(new_n463), .ZN(new_n942));
  XNOR2_X1  g517(.A(KEYINPUT66), .B(G2105), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n481), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT4), .B1(new_n944), .B2(G138), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n939), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(G160), .A2(G40), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(G1996), .A3(new_n708), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT111), .ZN(new_n952));
  INV_X1    g527(.A(G2067), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n755), .B(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(G1996), .B2(new_n708), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n952), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n811), .A2(new_n813), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n811), .A2(new_n813), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n950), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(G290), .A2(G1986), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT110), .Z(new_n962));
  INV_X1    g537(.A(G1986), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n962), .B1(new_n963), .B2(new_n820), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n960), .B1(new_n950), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n967), .B(new_n939), .C1(new_n942), .C2(new_n945), .ZN(new_n968));
  INV_X1    g543(.A(G40), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n472), .A2(new_n475), .A3(new_n969), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  AOI211_X1 g546(.A(KEYINPUT113), .B(new_n967), .C1(new_n502), .C2(new_n939), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT113), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(new_n946), .B2(KEYINPUT50), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n971), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT114), .B1(new_n975), .B2(G2090), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n968), .A2(new_n970), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n501), .A2(new_n499), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n463), .B1(new_n495), .B2(new_n496), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n980), .B2(new_n494), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT113), .B1(new_n981), .B2(new_n967), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n946), .A2(new_n973), .A3(KEYINPUT50), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n977), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n985), .A3(new_n763), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n949), .B1(new_n947), .B2(new_n946), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n939), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n981), .A2(KEYINPUT112), .A3(KEYINPUT45), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n987), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n785), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n976), .A2(new_n986), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(G303), .A2(G8), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n997), .B(KEYINPUT55), .Z(new_n998));
  NAND4_X1  g573(.A1(new_n976), .A2(new_n986), .A3(KEYINPUT115), .A4(new_n993), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n996), .A2(G8), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  OR2_X1    g576(.A1(new_n577), .A2(G1981), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n577), .A2(G1981), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT118), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(KEYINPUT49), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1002), .B(new_n1003), .C1(new_n1005), .C2(KEYINPUT49), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(new_n981), .B2(new_n970), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n564), .A2(new_n565), .A3(G1976), .A4(new_n566), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(new_n1015), .A3(new_n1010), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n1017));
  INV_X1    g592(.A(G1976), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1010), .A2(new_n1013), .A3(new_n1018), .A4(G288), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1017), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1021), .A2(new_n1014), .A3(new_n1015), .A4(new_n1010), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1011), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(new_n1018), .A3(new_n872), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n1002), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1001), .A2(new_n1023), .B1(new_n1010), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n998), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n977), .B1(KEYINPUT50), .B2(new_n946), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n992), .A2(new_n785), .B1(new_n1029), .B2(new_n763), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1028), .B1(new_n1009), .B2(new_n1030), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1000), .A2(new_n1023), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n948), .A2(new_n970), .A3(new_n988), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n761), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n975), .B2(G2084), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT122), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(KEYINPUT122), .B(new_n1034), .C1(new_n975), .C2(G2084), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(KEYINPUT51), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G2084), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n984), .A2(new_n1040), .B1(new_n761), .B2(new_n1033), .ZN(new_n1041));
  OAI21_X1  g616(.A(G168), .B1(new_n1041), .B2(KEYINPUT51), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1039), .A2(G8), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1037), .A2(G168), .A3(new_n1038), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n1045), .B2(G8), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT62), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1032), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1045), .A2(G8), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT51), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT62), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1039), .A2(G8), .A3(new_n1042), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(G2078), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n987), .A2(new_n988), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n984), .B2(G1961), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT123), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT123), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1056), .B(new_n1059), .C1(new_n984), .C2(G1961), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1054), .B1(new_n992), .B2(G2078), .ZN(new_n1062));
  AOI21_X1  g637(.A(G301), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1053), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1027), .B1(new_n1048), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT124), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n987), .A2(new_n990), .A3(new_n991), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n1055), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n975), .A2(new_n774), .ZN(new_n1069));
  AND4_X1   g644(.A1(G301), .A2(new_n1068), .A3(new_n1062), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1060), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1059), .B1(new_n1069), .B2(new_n1056), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1062), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1070), .B1(new_n1073), .B2(G171), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1066), .B1(new_n1074), .B2(KEYINPUT54), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n1076));
  OAI211_X1 g651(.A(KEYINPUT124), .B(new_n1076), .C1(new_n1063), .C2(new_n1070), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1000), .A2(new_n1023), .A3(new_n1031), .ZN(new_n1079));
  OAI211_X1 g654(.A(G301), .B(new_n1062), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1068), .A2(new_n1062), .A3(new_n1069), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G171), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1080), .A2(KEYINPUT54), .A3(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1078), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1996), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1067), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n981), .A2(new_n970), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT58), .B(G1341), .Z(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n546), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1092), .B(KEYINPUT59), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1029), .A2(G1956), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT56), .B(G2072), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1067), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n1097));
  XNOR2_X1  g672(.A(G299), .B(new_n1097), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT120), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT61), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(KEYINPUT120), .B(KEYINPUT61), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1093), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1089), .A2(G2067), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n975), .B2(new_n743), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(KEYINPUT119), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n1109));
  AOI211_X1 g684(.A(new_n1109), .B(new_n1106), .C1(new_n975), .C2(new_n743), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT60), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(KEYINPUT121), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT60), .ZN(new_n1113));
  OAI22_X1  g688(.A1(new_n984), .A2(G1348), .B1(G2067), .B2(new_n1089), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1109), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1107), .A2(KEYINPUT119), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1113), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n603), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1111), .A2(KEYINPUT121), .A3(new_n595), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1112), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1122), .A2(KEYINPUT60), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1105), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1122), .A2(new_n1099), .A3(new_n595), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1125), .A2(new_n1100), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1065), .B1(new_n1086), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT63), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1041), .A2(new_n1009), .A3(G286), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1129), .B1(new_n1079), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n996), .A2(G8), .A3(new_n999), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1129), .B1(new_n1133), .B2(new_n1028), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(new_n1000), .A3(new_n1023), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1132), .B1(new_n1135), .B2(new_n1131), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n966), .B1(new_n1128), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n950), .A2(new_n1087), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT46), .ZN(new_n1139));
  INV_X1    g714(.A(new_n954), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n950), .B1(new_n1140), .B2(new_n708), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  XOR2_X1   g717(.A(new_n1142), .B(KEYINPUT47), .Z(new_n1143));
  NAND2_X1  g718(.A1(new_n956), .A2(new_n958), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(G2067), .B2(new_n755), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1143), .B1(new_n1145), .B2(new_n950), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n962), .A2(new_n949), .A3(new_n948), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT48), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1146), .B1(new_n1148), .B2(new_n960), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n938), .B1(new_n1137), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1027), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1064), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1079), .B1(new_n1085), .B2(KEYINPUT62), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1078), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1154), .B(new_n1136), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n965), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1149), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1158), .A2(KEYINPUT125), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1150), .A2(new_n1160), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g736(.A1(G229), .A2(new_n461), .ZN(new_n1163));
  NAND3_X1  g737(.A1(new_n641), .A2(new_n1163), .A3(new_n658), .ZN(new_n1164));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n1165));
  NOR2_X1   g739(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g740(.A(new_n1166), .B1(new_n864), .B2(new_n867), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1168));
  OAI211_X1 g742(.A(new_n1167), .B(new_n1168), .C1(new_n934), .C2(new_n935), .ZN(G225));
  INV_X1    g743(.A(G225), .ZN(G308));
endmodule


