//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n557, new_n558, new_n559, new_n560, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n571, new_n572, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n632,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G221), .A4(G218), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  OR2_X1    g028(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  NAND2_X1  g031(.A1(new_n451), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT68), .B(G2105), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT69), .B(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n468), .A2(new_n469), .B1(new_n471), .B2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n464), .A2(KEYINPUT69), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n473), .A2(new_n475), .A3(KEYINPUT3), .ZN(new_n476));
  AND2_X1   g051(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n476), .A2(G137), .A3(new_n479), .A4(new_n463), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n476), .A2(new_n463), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(new_n479), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT70), .Z(new_n486));
  OAI221_X1 g061(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n479), .C2(G112), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n483), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(G162));
  NAND4_X1  g065(.A1(new_n476), .A2(G138), .A3(new_n479), .A4(new_n463), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  AND2_X1   g067(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n493));
  NOR2_X1   g068(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n463), .B(new_n465), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n469), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n492), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G2105), .ZN(new_n501));
  OR2_X1    g076(.A1(new_n501), .A2(G114), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT71), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n501), .A2(G114), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(new_n503), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n476), .A2(G126), .A3(G2105), .A4(new_n463), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n500), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT74), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT74), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(new_n517), .A3(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(new_n514), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT73), .A2(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(KEYINPUT6), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n519), .A2(new_n523), .A3(G543), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G50), .ZN(new_n526));
  OR2_X1    g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n529), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n521), .A2(new_n522), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n519), .A2(new_n523), .A3(new_n529), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G88), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n526), .A2(new_n533), .A3(new_n535), .ZN(G303));
  INV_X1    g111(.A(G303), .ZN(G166));
  INV_X1    g112(.A(KEYINPUT75), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n527), .A2(new_n528), .ZN(new_n539));
  NAND2_X1  g114(.A1(G63), .A2(G651), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n529), .A2(KEYINPUT75), .A3(G63), .A4(G651), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT76), .B(G51), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n519), .A2(new_n523), .A3(G543), .A4(new_n544), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n519), .A2(new_n523), .A3(G89), .A4(new_n529), .ZN(new_n546));
  NAND3_X1  g121(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n543), .A2(new_n545), .A3(new_n546), .A4(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT77), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n541), .A2(new_n542), .B1(new_n549), .B2(new_n548), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n554), .A2(KEYINPUT77), .A3(new_n545), .A4(new_n546), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n553), .A2(new_n555), .ZN(G168));
  NAND2_X1  g131(.A1(new_n525), .A2(G52), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n529), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n558), .A2(new_n532), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n534), .A2(G90), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(G301));
  INV_X1    g136(.A(G301), .ZN(G171));
  NAND2_X1  g137(.A1(new_n525), .A2(G43), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n529), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n532), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n534), .A2(G81), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  XNOR2_X1  g148(.A(KEYINPUT79), .B(G65), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n529), .A2(new_n574), .B1(G78), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n514), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(G91), .B2(new_n534), .ZN(new_n577));
  AND2_X1   g152(.A1(KEYINPUT78), .A2(G53), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n519), .A2(new_n523), .A3(G543), .A4(new_n578), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT9), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(G299));
  INV_X1    g156(.A(G168), .ZN(G286));
  NAND2_X1  g157(.A1(new_n525), .A2(G49), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n534), .A2(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n529), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(new_n529), .A2(G61), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(KEYINPUT80), .B1(G73), .B2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n527), .B2(new_n528), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n532), .B1(new_n588), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n519), .A2(new_n523), .A3(G86), .A4(new_n529), .ZN(new_n595));
  INV_X1    g170(.A(G48), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n524), .B2(new_n596), .ZN(new_n597));
  NOR3_X1   g172(.A1(new_n593), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n597), .ZN(new_n599));
  INV_X1    g174(.A(new_n592), .ZN(new_n600));
  NAND2_X1  g175(.A1(G73), .A2(G543), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n590), .B2(new_n591), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n531), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(KEYINPUT81), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n598), .A2(new_n604), .ZN(G305));
  XOR2_X1   g180(.A(KEYINPUT82), .B(G47), .Z(new_n606));
  NAND2_X1  g181(.A1(new_n525), .A2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n529), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(new_n532), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n534), .A2(G85), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n607), .A2(new_n609), .A3(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT83), .Z(new_n613));
  NAND4_X1  g188(.A1(new_n519), .A2(new_n523), .A3(G92), .A4(new_n529), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT10), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n524), .A2(KEYINPUT84), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT84), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n519), .A2(new_n523), .A3(new_n617), .A4(G543), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n616), .A2(G54), .A3(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n529), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n620), .A2(new_n514), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT85), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n619), .A2(KEYINPUT85), .A3(new_n621), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n615), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n613), .B1(G868), .B2(new_n626), .ZN(G284));
  OAI21_X1  g202(.A(new_n613), .B1(G868), .B2(new_n626), .ZN(G321));
  NOR2_X1   g203(.A1(G299), .A2(G868), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(G868), .B2(G168), .ZN(G297));
  XNOR2_X1  g205(.A(G297), .B(KEYINPUT86), .ZN(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n626), .B1(new_n632), .B2(G860), .ZN(G148));
  NAND2_X1  g208(.A1(new_n626), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G868), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(G868), .B2(new_n568), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR3_X1   g212(.A1(new_n466), .A2(new_n470), .A3(G2105), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT88), .B(KEYINPUT13), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2100), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n488), .A2(G135), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n484), .A2(G123), .ZN(new_n645));
  OAI221_X1 g220(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n479), .C2(G111), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n647), .A2(G2096), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(G2096), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n643), .A2(new_n648), .A3(new_n649), .ZN(G156));
  XOR2_X1   g225(.A(G2451), .B(G2454), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT14), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n658), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n654), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(G14), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n663), .B2(new_n661), .ZN(G401));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2100), .ZN(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n669), .B2(KEYINPUT18), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2096), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT19), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n681), .A2(new_n682), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n680), .A2(new_n685), .A3(new_n683), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n680), .A2(new_n685), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n688));
  AOI211_X1 g263(.A(new_n684), .B(new_n686), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(new_n687), .B2(new_n688), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  XNOR2_X1  g272(.A(KEYINPUT96), .B(KEYINPUT23), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G20), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G299), .B2(G16), .ZN(new_n702));
  INV_X1    g277(.A(G1956), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(G16), .A2(G19), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n568), .B2(G16), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(G1341), .ZN(new_n707));
  NOR2_X1   g282(.A1(G171), .A2(new_n699), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G5), .B2(new_n699), .ZN(new_n709));
  INV_X1    g284(.A(G1961), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G2078), .ZN(new_n712));
  NAND2_X1  g287(.A1(G164), .A2(G29), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G27), .B2(G29), .ZN(new_n714));
  AOI211_X1 g289(.A(new_n707), .B(new_n711), .C1(new_n712), .C2(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n712), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT24), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(G34), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(G34), .ZN(new_n719));
  AOI21_X1  g294(.A(G29), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n481), .B2(G29), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G2084), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n709), .A2(new_n710), .B1(G1341), .B2(new_n706), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n715), .A2(new_n716), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(G168), .A2(new_n699), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n699), .B2(G21), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  AOI211_X1 g302(.A(new_n704), .B(new_n724), .C1(G1966), .C2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT30), .B(G28), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  OR2_X1    g305(.A1(KEYINPUT31), .A2(G11), .ZN(new_n731));
  NAND2_X1  g306(.A1(KEYINPUT31), .A2(G11), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n729), .A2(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n647), .B2(new_n730), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT95), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n730), .A2(G26), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT28), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n488), .A2(G140), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n484), .A2(G128), .ZN(new_n739));
  OAI221_X1 g314(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n479), .C2(G116), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n737), .B1(new_n742), .B2(new_n730), .ZN(new_n743));
  INV_X1    g318(.A(G2067), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n730), .A2(G33), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n479), .A2(G103), .A3(G2104), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT25), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n488), .A2(G139), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n463), .A2(new_n465), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n751), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n749), .B(new_n750), .C1(new_n479), .C2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT93), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n746), .B1(new_n755), .B2(new_n730), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n745), .B1(new_n756), .B2(G2072), .ZN(new_n757));
  AOI211_X1 g332(.A(new_n735), .B(new_n757), .C1(G2072), .C2(new_n756), .ZN(new_n758));
  NOR2_X1   g333(.A1(G29), .A2(G35), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G162), .B2(G29), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT29), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2090), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n488), .A2(G141), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n484), .A2(G129), .ZN(new_n764));
  NAND3_X1  g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT26), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n471), .A2(G105), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n763), .A2(new_n764), .A3(new_n769), .ZN(new_n770));
  MUX2_X1   g345(.A(G32), .B(new_n770), .S(G29), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT94), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT27), .B(G1996), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G1966), .B2(new_n727), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n762), .A2(new_n775), .ZN(new_n776));
  AND3_X1   g351(.A1(new_n728), .A2(new_n758), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n699), .A2(G22), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G166), .B2(new_n699), .ZN(new_n779));
  INV_X1    g354(.A(G1971), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n699), .A2(G23), .ZN(new_n782));
  INV_X1    g357(.A(G288), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n699), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT33), .B(G1976), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  MUX2_X1   g361(.A(G6), .B(G305), .S(G16), .Z(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT32), .B(G1981), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n781), .B(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n788), .B2(new_n787), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT34), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n730), .A2(G25), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT90), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n488), .A2(G131), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n484), .A2(G119), .ZN(new_n797));
  NOR2_X1   g372(.A1(G95), .A2(G2105), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT91), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G107), .C2(new_n479), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n796), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n795), .B1(new_n802), .B2(new_n730), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT35), .B(G1991), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(G16), .A2(G24), .ZN(new_n806));
  XOR2_X1   g381(.A(G290), .B(KEYINPUT92), .Z(new_n807));
  AOI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(G16), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(G1986), .Z(new_n809));
  NAND4_X1  g384(.A1(new_n792), .A2(new_n793), .A3(new_n805), .A4(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT36), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n699), .A2(G4), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n626), .B2(new_n699), .ZN(new_n813));
  INV_X1    g388(.A(G1348), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n777), .A2(new_n811), .A3(new_n815), .ZN(G150));
  INV_X1    g391(.A(G150), .ZN(G311));
  NAND2_X1  g392(.A1(new_n525), .A2(G55), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n529), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(new_n532), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n534), .A2(G93), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n818), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G860), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT37), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n626), .A2(G559), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT38), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n567), .B(new_n822), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT97), .ZN(new_n831));
  INV_X1    g406(.A(G860), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n828), .B2(new_n829), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n824), .B1(new_n831), .B2(new_n833), .ZN(G145));
  NAND2_X1  g409(.A1(new_n488), .A2(G142), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT98), .Z(new_n836));
  OAI221_X1 g411(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n479), .C2(G118), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n484), .A2(G130), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n801), .B(new_n640), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT99), .ZN(new_n843));
  OR3_X1    g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n841), .B2(new_n842), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n755), .B(new_n770), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n741), .B(new_n512), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n846), .A2(new_n847), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n844), .B(new_n845), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n850), .ZN(new_n852));
  INV_X1    g427(.A(new_n845), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n852), .A2(new_n853), .A3(new_n848), .ZN(new_n854));
  XNOR2_X1  g429(.A(G160), .B(new_n647), .ZN(new_n855));
  XNOR2_X1  g430(.A(G162), .B(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n851), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(G37), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n856), .B1(new_n851), .B2(new_n854), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(KEYINPUT100), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n862));
  AOI211_X1 g437(.A(new_n862), .B(new_n856), .C1(new_n851), .C2(new_n854), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n859), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n866));
  XNOR2_X1  g441(.A(G303), .B(G288), .ZN(new_n867));
  INV_X1    g442(.A(G290), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n598), .B2(new_n604), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n594), .B1(new_n593), .B2(new_n597), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n599), .A2(KEYINPUT81), .A3(new_n603), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n871), .A3(G290), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n867), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n867), .B1(new_n869), .B2(new_n872), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n866), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n869), .A2(new_n872), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n783), .A2(G303), .ZN(new_n878));
  NOR2_X1   g453(.A1(G166), .A2(G288), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(KEYINPUT102), .A3(new_n873), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT42), .ZN(new_n884));
  OR3_X1    g459(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT42), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT103), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n634), .B(new_n827), .ZN(new_n887));
  INV_X1    g462(.A(new_n615), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n619), .A2(KEYINPUT85), .A3(new_n621), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT85), .B1(new_n619), .B2(new_n621), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(G299), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g468(.A(G299), .B(new_n888), .C1(new_n889), .C2(new_n890), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n887), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT101), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n626), .B2(G299), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n891), .A2(KEYINPUT101), .A3(new_n892), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n894), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n901), .B1(new_n626), .B2(G299), .ZN(new_n902));
  AOI22_X1  g477(.A1(new_n900), .A2(new_n901), .B1(new_n893), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n896), .B1(new_n903), .B2(new_n887), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n886), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n884), .A2(KEYINPUT103), .A3(new_n885), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n886), .A2(new_n904), .ZN(new_n908));
  OAI21_X1  g483(.A(G868), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(G868), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n822), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(G295));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n911), .ZN(G331));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n553), .A2(G301), .A3(new_n555), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n567), .B(new_n822), .Z(new_n917));
  AOI21_X1  g492(.A(G301), .B1(new_n553), .B2(new_n555), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n916), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n827), .B1(new_n915), .B2(new_n918), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n895), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n898), .A2(new_n902), .A3(new_n899), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n895), .A2(new_n901), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n921), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n827), .B(KEYINPUT104), .C1(new_n915), .C2(new_n918), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n920), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n923), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT107), .B1(new_n931), .B2(new_n882), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n926), .A2(new_n930), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n933), .B(new_n883), .C1(new_n934), .C2(new_n923), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n928), .A2(new_n895), .A3(new_n920), .A4(new_n929), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n920), .A2(new_n921), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n882), .B(new_n938), .C1(new_n903), .C2(new_n939), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n940), .A2(new_n858), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n936), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n938), .B1(new_n903), .B2(new_n939), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n938), .B(KEYINPUT105), .C1(new_n903), .C2(new_n939), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n883), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n937), .B1(new_n947), .B2(new_n941), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n942), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AOI211_X1 g525(.A(KEYINPUT106), .B(new_n937), .C1(new_n947), .C2(new_n941), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n914), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n936), .A2(KEYINPUT43), .A3(new_n941), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT43), .B1(new_n947), .B2(new_n941), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT44), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(G397));
  XNOR2_X1  g531(.A(new_n741), .B(new_n744), .ZN(new_n957));
  INV_X1    g532(.A(G1996), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n770), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n802), .A2(new_n804), .ZN(new_n961));
  OAI22_X1  g536(.A1(new_n960), .A2(new_n961), .B1(G2067), .B2(new_n741), .ZN(new_n962));
  INV_X1    g537(.A(G1384), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n491), .A2(KEYINPUT4), .B1(new_n496), .B2(new_n498), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n509), .A2(new_n510), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n472), .A2(G40), .A3(new_n480), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n962), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n770), .B1(KEYINPUT46), .B2(new_n958), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n957), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n970), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT46), .B1(new_n970), .B2(new_n958), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n975), .A2(KEYINPUT125), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(KEYINPUT125), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n978), .B(KEYINPUT47), .Z(new_n979));
  INV_X1    g554(.A(new_n960), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n801), .B(new_n804), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n970), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT126), .ZN(new_n984));
  NOR4_X1   g559(.A1(new_n968), .A2(G1986), .A3(G290), .A4(new_n969), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT48), .Z(new_n986));
  AOI211_X1 g561(.A(new_n971), .B(new_n979), .C1(new_n984), .C2(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n472), .A2(G40), .A3(new_n480), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n990));
  AOI21_X1  g565(.A(G1384), .B1(new_n500), .B2(new_n511), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n966), .A2(KEYINPUT108), .A3(KEYINPUT50), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n989), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(KEYINPUT115), .B(G2084), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT116), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n991), .A2(KEYINPUT114), .A3(KEYINPUT45), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n969), .B1(new_n966), .B2(new_n967), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT45), .B(new_n963), .C1(new_n964), .C2(new_n965), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1966), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n995), .A2(new_n1007), .A3(new_n996), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n998), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1009), .A2(G8), .A3(G168), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT63), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n968), .A2(new_n988), .A3(new_n1001), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n780), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n969), .B1(new_n991), .B2(new_n992), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n966), .A2(KEYINPUT108), .A3(KEYINPUT50), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT108), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1014), .B1(new_n1018), .B2(G2090), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT109), .ZN(new_n1020));
  NAND2_X1  g595(.A1(G303), .A2(G8), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1021), .B(KEYINPUT55), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT109), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1024), .B(new_n1014), .C1(new_n1018), .C2(G2090), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1020), .A2(G8), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n966), .A2(new_n969), .ZN(new_n1027));
  INV_X1    g602(.A(G8), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1976), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(new_n1030), .B2(G288), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT52), .B1(G288), .B2(new_n1030), .ZN(new_n1033));
  XOR2_X1   g608(.A(new_n1033), .B(KEYINPUT111), .Z(new_n1034));
  NAND2_X1  g609(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1031), .B1(KEYINPUT110), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1029), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n1040));
  OAI21_X1  g615(.A(G1981), .B1(new_n593), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n599), .A2(new_n603), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT49), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1039), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1043), .A2(KEYINPUT49), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1036), .A2(new_n1038), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1020), .A2(G8), .A3(new_n1025), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n1022), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1012), .A2(new_n1026), .A3(new_n1048), .A4(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n992), .B1(new_n512), .B2(new_n963), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n989), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G2090), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1053), .A2(new_n1054), .B1(new_n1013), .B2(new_n780), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(G8), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1022), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1059), .A2(new_n1048), .A3(new_n1026), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1011), .B1(new_n1060), .B2(new_n1010), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1051), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1008), .A2(new_n1006), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1007), .B1(new_n995), .B2(new_n996), .ZN(new_n1064));
  OAI21_X1  g639(.A(G8), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n1066));
  NAND2_X1  g641(.A1(G286), .A2(G8), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1067), .B(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1065), .A2(new_n1066), .A3(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1069), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT51), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1069), .B1(new_n1009), .B2(G8), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1071), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1059), .A2(new_n1048), .A3(new_n1026), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n968), .A2(new_n712), .A3(new_n988), .A4(new_n1001), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(G2078), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n999), .A2(new_n1000), .A3(new_n1003), .A4(new_n1080), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1079), .B(new_n1081), .C1(new_n995), .C2(G1961), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(G171), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT121), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(new_n1085), .A3(G171), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1075), .A2(KEYINPUT62), .A3(new_n1076), .A4(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(new_n1030), .A3(new_n783), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1042), .A2(G1981), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1039), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1026), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1092), .B1(new_n1093), .B2(new_n1048), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1062), .A2(new_n1088), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT62), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1087), .B(new_n1076), .C1(new_n1075), .C2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(G299), .B(KEYINPUT57), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n703), .B1(new_n989), .B2(new_n1052), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n968), .A2(new_n988), .A3(new_n1001), .A4(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1099), .B1(KEYINPUT117), .B2(new_n1101), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1101), .A2(KEYINPUT117), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1098), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1018), .A2(new_n814), .B1(new_n744), .B2(new_n1027), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1104), .B1(new_n891), .B2(new_n1105), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1101), .A2(KEYINPUT117), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1098), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1101), .A2(KEYINPUT117), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .A4(new_n1099), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1027), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n995), .A2(G1348), .B1(G2067), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT60), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1113), .A2(new_n1114), .A3(new_n626), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n891), .B1(new_n1105), .B2(KEYINPUT60), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT118), .B(G1996), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n968), .A2(new_n988), .A3(new_n1001), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  XOR2_X1   g697(.A(KEYINPUT58), .B(G1341), .Z(new_n1123));
  NAND2_X1  g698(.A1(new_n1112), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n568), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT59), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1129), .B(new_n568), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1118), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1104), .A2(new_n1110), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT61), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1104), .A2(new_n1110), .A3(KEYINPUT61), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1111), .B1(new_n1132), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1018), .A2(new_n710), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n1078), .B(G2078), .C1(new_n988), .C2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n969), .A2(KEYINPUT122), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1141), .A2(new_n1001), .A3(new_n968), .A4(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1139), .A2(new_n1079), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(G171), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT54), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n1082), .B2(G171), .ZN(new_n1148));
  OR3_X1    g723(.A1(new_n1082), .A2(new_n1147), .A3(G171), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1150), .A2(new_n1060), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1138), .A2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1139), .A2(G301), .A3(new_n1079), .A4(new_n1143), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1084), .A2(new_n1086), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1155), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1097), .B1(new_n1152), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1075), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1095), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n982), .ZN(new_n1163));
  XOR2_X1   g738(.A(G290), .B(G1986), .Z(new_n1164));
  AOI211_X1 g739(.A(new_n969), .B(new_n968), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n987), .B1(new_n1162), .B2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g741(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1168));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n1169));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OR2_X1    g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1171));
  AND3_X1   g745(.A1(new_n696), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  OAI211_X1 g746(.A(new_n864), .B(new_n1172), .C1(new_n950), .C2(new_n951), .ZN(G225));
  INV_X1    g747(.A(G225), .ZN(G308));
endmodule


