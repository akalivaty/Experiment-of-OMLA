

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X1 U325 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U326 ( .A(n431), .B(n430), .Z(n293) );
  AND2_X1 U327 ( .A1(G230GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U328 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n295) );
  NAND2_X1 U329 ( .A1(n408), .A2(n565), .ZN(n296) );
  XNOR2_X1 U330 ( .A(KEYINPUT25), .B(KEYINPUT97), .ZN(n406) );
  XNOR2_X1 U331 ( .A(n407), .B(n406), .ZN(n411) );
  XNOR2_X1 U332 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U333 ( .A(n425), .B(n294), .ZN(n427) );
  XNOR2_X1 U334 ( .A(n298), .B(KEYINPUT93), .ZN(n299) );
  XNOR2_X1 U335 ( .A(n388), .B(n387), .ZN(n392) );
  XNOR2_X1 U336 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n465) );
  XNOR2_X1 U337 ( .A(n388), .B(n299), .ZN(n301) );
  XNOR2_X1 U338 ( .A(n432), .B(n293), .ZN(n433) );
  XNOR2_X1 U339 ( .A(n466), .B(n465), .ZN(n527) );
  XNOR2_X1 U340 ( .A(n434), .B(n433), .ZN(n438) );
  NOR2_X1 U341 ( .A1(n496), .A2(n508), .ZN(n452) );
  XNOR2_X1 U342 ( .A(n471), .B(KEYINPUT124), .ZN(n584) );
  INV_X1 U343 ( .A(G106GAT), .ZN(n476) );
  XNOR2_X1 U344 ( .A(n473), .B(G204GAT), .ZN(n474) );
  XNOR2_X1 U345 ( .A(n476), .B(KEYINPUT44), .ZN(n477) );
  XNOR2_X1 U346 ( .A(n453), .B(G92GAT), .ZN(n454) );
  XNOR2_X1 U347 ( .A(n475), .B(n474), .ZN(G1353GAT) );
  XNOR2_X1 U348 ( .A(n455), .B(n454), .ZN(G1337GAT) );
  XNOR2_X1 U349 ( .A(G190GAT), .B(KEYINPUT18), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n295), .B(n297), .ZN(n388) );
  AND2_X1 U351 ( .A1(G226GAT), .A2(G233GAT), .ZN(n298) );
  INV_X1 U352 ( .A(KEYINPUT94), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n306) );
  XOR2_X1 U354 ( .A(G183GAT), .B(G211GAT), .Z(n334) );
  XNOR2_X1 U355 ( .A(n334), .B(KEYINPUT92), .ZN(n304) );
  XNOR2_X1 U356 ( .A(G176GAT), .B(G92GAT), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n302), .B(G64GAT), .ZN(n426) );
  INV_X1 U358 ( .A(n426), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n306), .B(n305), .ZN(n311) );
  XNOR2_X1 U361 ( .A(G169GAT), .B(G36GAT), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n307), .B(G8GAT), .ZN(n445) );
  XOR2_X1 U363 ( .A(G204GAT), .B(KEYINPUT21), .Z(n309) );
  XNOR2_X1 U364 ( .A(G197GAT), .B(G218GAT), .ZN(n308) );
  XNOR2_X1 U365 ( .A(n309), .B(n308), .ZN(n371) );
  XNOR2_X1 U366 ( .A(n445), .B(n371), .ZN(n310) );
  XNOR2_X1 U367 ( .A(n311), .B(n310), .ZN(n513) );
  XOR2_X1 U368 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n313) );
  XNOR2_X1 U369 ( .A(G190GAT), .B(G162GAT), .ZN(n312) );
  XNOR2_X1 U370 ( .A(n313), .B(n312), .ZN(n329) );
  XOR2_X1 U371 ( .A(G106GAT), .B(G218GAT), .Z(n315) );
  XNOR2_X1 U372 ( .A(G134GAT), .B(KEYINPUT73), .ZN(n314) );
  XNOR2_X1 U373 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U374 ( .A(n316), .B(KEYINPUT74), .Z(n318) );
  XOR2_X1 U375 ( .A(G99GAT), .B(G85GAT), .Z(n425) );
  XNOR2_X1 U376 ( .A(G36GAT), .B(n425), .ZN(n317) );
  XNOR2_X1 U377 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U378 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n320) );
  NAND2_X1 U379 ( .A1(G232GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U380 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U381 ( .A(n322), .B(n321), .Z(n327) );
  XOR2_X1 U382 ( .A(KEYINPUT7), .B(G50GAT), .Z(n324) );
  XNOR2_X1 U383 ( .A(G43GAT), .B(G29GAT), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U385 ( .A(KEYINPUT8), .B(n325), .Z(n440) );
  XNOR2_X1 U386 ( .A(n440), .B(G92GAT), .ZN(n326) );
  XNOR2_X1 U387 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U388 ( .A(n329), .B(n328), .Z(n574) );
  XOR2_X1 U389 ( .A(KEYINPUT36), .B(n574), .Z(n585) );
  XNOR2_X1 U390 ( .A(G1GAT), .B(G127GAT), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n330), .B(G57GAT), .ZN(n361) );
  XOR2_X1 U392 ( .A(n361), .B(KEYINPUT75), .Z(n332) );
  NAND2_X1 U393 ( .A1(G231GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U394 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U395 ( .A(n334), .B(n333), .Z(n338) );
  XOR2_X1 U396 ( .A(G15GAT), .B(G22GAT), .Z(n439) );
  XOR2_X1 U397 ( .A(KEYINPUT13), .B(KEYINPUT69), .Z(n336) );
  XNOR2_X1 U398 ( .A(G71GAT), .B(KEYINPUT70), .ZN(n335) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n429) );
  XNOR2_X1 U400 ( .A(n439), .B(n429), .ZN(n337) );
  XNOR2_X1 U401 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U402 ( .A(G64GAT), .B(G78GAT), .Z(n340) );
  XNOR2_X1 U403 ( .A(G8GAT), .B(G155GAT), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U405 ( .A(n342), .B(n341), .Z(n350) );
  XOR2_X1 U406 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n344) );
  XNOR2_X1 U407 ( .A(KEYINPUT12), .B(KEYINPUT80), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U409 ( .A(KEYINPUT76), .B(KEYINPUT15), .Z(n346) );
  XNOR2_X1 U410 ( .A(KEYINPUT79), .B(KEYINPUT77), .ZN(n345) );
  XNOR2_X1 U411 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U412 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U413 ( .A(n350), .B(n349), .Z(n582) );
  XOR2_X1 U414 ( .A(KEYINPUT6), .B(KEYINPUT89), .Z(n352) );
  XNOR2_X1 U415 ( .A(G29GAT), .B(G85GAT), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U417 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n354) );
  XNOR2_X1 U418 ( .A(KEYINPUT90), .B(KEYINPUT5), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U420 ( .A(n356), .B(n355), .Z(n366) );
  XNOR2_X1 U421 ( .A(G155GAT), .B(KEYINPUT87), .ZN(n357) );
  XNOR2_X1 U422 ( .A(n357), .B(KEYINPUT3), .ZN(n358) );
  XOR2_X1 U423 ( .A(n358), .B(KEYINPUT2), .Z(n360) );
  XNOR2_X1 U424 ( .A(G141GAT), .B(G162GAT), .ZN(n359) );
  XNOR2_X1 U425 ( .A(n360), .B(n359), .ZN(n384) );
  XOR2_X1 U426 ( .A(G120GAT), .B(G148GAT), .Z(n435) );
  XOR2_X1 U427 ( .A(n435), .B(n361), .Z(n363) );
  NAND2_X1 U428 ( .A1(G225GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n384), .B(n364), .ZN(n365) );
  XNOR2_X1 U431 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U432 ( .A(KEYINPUT81), .B(G134GAT), .Z(n368) );
  XNOR2_X1 U433 ( .A(KEYINPUT82), .B(KEYINPUT0), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U435 ( .A(G113GAT), .B(n369), .ZN(n393) );
  XNOR2_X1 U436 ( .A(n370), .B(n393), .ZN(n415) );
  XOR2_X1 U437 ( .A(G106GAT), .B(G78GAT), .Z(n436) );
  XOR2_X1 U438 ( .A(n436), .B(n371), .Z(n373) );
  XNOR2_X1 U439 ( .A(G50GAT), .B(KEYINPUT73), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U441 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n375) );
  NAND2_X1 U442 ( .A1(G228GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U443 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U444 ( .A(n377), .B(n376), .Z(n382) );
  XOR2_X1 U445 ( .A(KEYINPUT88), .B(G148GAT), .Z(n379) );
  XNOR2_X1 U446 ( .A(G22GAT), .B(G211GAT), .ZN(n378) );
  XNOR2_X1 U447 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U448 ( .A(n380), .B(KEYINPUT23), .ZN(n381) );
  XNOR2_X1 U449 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U450 ( .A(n384), .B(n383), .ZN(n558) );
  NAND2_X1 U451 ( .A1(G227GAT), .A2(G233GAT), .ZN(n386) );
  INV_X1 U452 ( .A(G99GAT), .ZN(n385) );
  XOR2_X1 U453 ( .A(G71GAT), .B(G176GAT), .Z(n390) );
  XNOR2_X1 U454 ( .A(G169GAT), .B(G183GAT), .ZN(n389) );
  XOR2_X1 U455 ( .A(n390), .B(n389), .Z(n391) );
  XNOR2_X1 U456 ( .A(n392), .B(n391), .ZN(n395) );
  XOR2_X1 U457 ( .A(G43GAT), .B(n393), .Z(n394) );
  XNOR2_X1 U458 ( .A(n395), .B(n394), .ZN(n403) );
  XOR2_X1 U459 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n397) );
  XNOR2_X1 U460 ( .A(G127GAT), .B(KEYINPUT85), .ZN(n396) );
  XNOR2_X1 U461 ( .A(n397), .B(n396), .ZN(n401) );
  XOR2_X1 U462 ( .A(G120GAT), .B(KEYINPUT83), .Z(n399) );
  XNOR2_X1 U463 ( .A(G15GAT), .B(KEYINPUT84), .ZN(n398) );
  XNOR2_X1 U464 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U465 ( .A(n401), .B(n400), .Z(n402) );
  XOR2_X1 U466 ( .A(n403), .B(n402), .Z(n408) );
  INV_X1 U467 ( .A(n408), .ZN(n562) );
  NOR2_X1 U468 ( .A1(n513), .A2(n562), .ZN(n404) );
  XOR2_X1 U469 ( .A(KEYINPUT96), .B(n404), .Z(n405) );
  NAND2_X1 U470 ( .A1(n558), .A2(n405), .ZN(n407) );
  XOR2_X1 U471 ( .A(n513), .B(KEYINPUT27), .Z(n416) );
  NOR2_X1 U472 ( .A1(n558), .A2(n408), .ZN(n409) );
  XNOR2_X1 U473 ( .A(n409), .B(KEYINPUT26), .ZN(n544) );
  NAND2_X1 U474 ( .A1(n416), .A2(n544), .ZN(n410) );
  NAND2_X1 U475 ( .A1(n411), .A2(n410), .ZN(n412) );
  XOR2_X1 U476 ( .A(KEYINPUT98), .B(n412), .Z(n413) );
  NOR2_X1 U477 ( .A1(n415), .A2(n413), .ZN(n414) );
  XNOR2_X1 U478 ( .A(KEYINPUT99), .B(n414), .ZN(n421) );
  XNOR2_X1 U479 ( .A(KEYINPUT91), .B(n415), .ZN(n520) );
  INV_X1 U480 ( .A(n416), .ZN(n417) );
  NOR2_X1 U481 ( .A1(n520), .A2(n417), .ZN(n525) );
  XNOR2_X1 U482 ( .A(KEYINPUT28), .B(n558), .ZN(n529) );
  NAND2_X1 U483 ( .A1(n525), .A2(n529), .ZN(n418) );
  NOR2_X1 U484 ( .A1(n408), .A2(n418), .ZN(n419) );
  XNOR2_X1 U485 ( .A(KEYINPUT95), .B(n419), .ZN(n420) );
  NAND2_X1 U486 ( .A1(n421), .A2(n420), .ZN(n482) );
  NAND2_X1 U487 ( .A1(n582), .A2(n482), .ZN(n422) );
  NOR2_X1 U488 ( .A1(n585), .A2(n422), .ZN(n424) );
  XNOR2_X1 U489 ( .A(KEYINPUT104), .B(KEYINPUT37), .ZN(n423) );
  XNOR2_X1 U490 ( .A(n424), .B(n423), .ZN(n496) );
  XOR2_X1 U491 ( .A(n428), .B(KEYINPUT33), .Z(n434) );
  XNOR2_X1 U492 ( .A(n429), .B(KEYINPUT31), .ZN(n432) );
  XOR2_X1 U493 ( .A(KEYINPUT71), .B(KEYINPUT32), .Z(n431) );
  XNOR2_X1 U494 ( .A(G204GAT), .B(G57GAT), .ZN(n430) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n479) );
  XOR2_X1 U497 ( .A(n479), .B(KEYINPUT41), .Z(n565) );
  XOR2_X1 U498 ( .A(n439), .B(G197GAT), .Z(n442) );
  XNOR2_X1 U499 ( .A(n440), .B(G113GAT), .ZN(n441) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n451) );
  XOR2_X1 U501 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n444) );
  XNOR2_X1 U502 ( .A(G141GAT), .B(G1GAT), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n449) );
  XOR2_X1 U504 ( .A(n445), .B(KEYINPUT29), .Z(n447) );
  NAND2_X1 U505 ( .A1(G229GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U506 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U507 ( .A(n449), .B(n448), .Z(n450) );
  XNOR2_X1 U508 ( .A(n451), .B(n450), .ZN(n577) );
  NAND2_X1 U509 ( .A1(n565), .A2(n577), .ZN(n508) );
  XOR2_X1 U510 ( .A(KEYINPUT110), .B(n452), .Z(n523) );
  NOR2_X1 U511 ( .A1(n513), .A2(n523), .ZN(n455) );
  XNOR2_X1 U512 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n453) );
  XOR2_X1 U513 ( .A(n582), .B(KEYINPUT114), .Z(n571) );
  INV_X1 U514 ( .A(n565), .ZN(n550) );
  NOR2_X1 U515 ( .A1(n577), .A2(n550), .ZN(n456) );
  XNOR2_X1 U516 ( .A(n456), .B(KEYINPUT46), .ZN(n457) );
  NOR2_X1 U517 ( .A1(n571), .A2(n457), .ZN(n458) );
  INV_X1 U518 ( .A(n574), .ZN(n556) );
  NAND2_X1 U519 ( .A1(n458), .A2(n556), .ZN(n459) );
  XNOR2_X1 U520 ( .A(n459), .B(KEYINPUT47), .ZN(n464) );
  NOR2_X1 U521 ( .A1(n585), .A2(n582), .ZN(n460) );
  XNOR2_X1 U522 ( .A(KEYINPUT45), .B(n460), .ZN(n461) );
  XOR2_X1 U523 ( .A(KEYINPUT68), .B(n577), .Z(n563) );
  INV_X1 U524 ( .A(n563), .ZN(n531) );
  NAND2_X1 U525 ( .A1(n461), .A2(n531), .ZN(n462) );
  NOR2_X1 U526 ( .A1(n462), .A2(n479), .ZN(n463) );
  NOR2_X1 U527 ( .A1(n464), .A2(n463), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n513), .B(KEYINPUT122), .ZN(n467) );
  NOR2_X1 U529 ( .A1(n527), .A2(n467), .ZN(n468) );
  XNOR2_X1 U530 ( .A(n468), .B(KEYINPUT54), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n469), .A2(n520), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n470), .B(KEYINPUT65), .ZN(n559) );
  NAND2_X1 U533 ( .A1(n544), .A2(n559), .ZN(n471) );
  INV_X1 U534 ( .A(n584), .ZN(n472) );
  NAND2_X1 U535 ( .A1(n479), .A2(n472), .ZN(n475) );
  XOR2_X1 U536 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n473) );
  NOR2_X1 U537 ( .A1(n529), .A2(n523), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(G1339GAT) );
  NOR2_X1 U539 ( .A1(n531), .A2(n479), .ZN(n480) );
  XOR2_X1 U540 ( .A(KEYINPUT72), .B(n480), .Z(n495) );
  NOR2_X1 U541 ( .A1(n574), .A2(n582), .ZN(n481) );
  XNOR2_X1 U542 ( .A(KEYINPUT16), .B(n481), .ZN(n483) );
  NAND2_X1 U543 ( .A1(n483), .A2(n482), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(KEYINPUT100), .ZN(n509) );
  OR2_X1 U545 ( .A1(n495), .A2(n509), .ZN(n492) );
  NOR2_X1 U546 ( .A1(n520), .A2(n492), .ZN(n486) );
  XNOR2_X1 U547 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(n487), .ZN(G1324GAT) );
  NOR2_X1 U550 ( .A1(n513), .A2(n492), .ZN(n488) );
  XOR2_X1 U551 ( .A(KEYINPUT102), .B(n488), .Z(n489) );
  XNOR2_X1 U552 ( .A(G8GAT), .B(n489), .ZN(G1325GAT) );
  NOR2_X1 U553 ( .A1(n562), .A2(n492), .ZN(n491) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n490) );
  XNOR2_X1 U555 ( .A(n491), .B(n490), .ZN(G1326GAT) );
  NOR2_X1 U556 ( .A1(n529), .A2(n492), .ZN(n494) );
  XNOR2_X1 U557 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n494), .B(n493), .ZN(G1327GAT) );
  XNOR2_X1 U559 ( .A(KEYINPUT38), .B(KEYINPUT105), .ZN(n498) );
  NOR2_X1 U560 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n506) );
  NOR2_X1 U562 ( .A1(n506), .A2(n520), .ZN(n500) );
  XNOR2_X1 U563 ( .A(KEYINPUT106), .B(KEYINPUT39), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U565 ( .A(G29GAT), .B(n501), .ZN(G1328GAT) );
  NOR2_X1 U566 ( .A1(n513), .A2(n506), .ZN(n502) );
  XOR2_X1 U567 ( .A(G36GAT), .B(n502), .Z(G1329GAT) );
  NOR2_X1 U568 ( .A1(n506), .A2(n562), .ZN(n504) );
  XNOR2_X1 U569 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n503) );
  XNOR2_X1 U570 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U571 ( .A(G43GAT), .B(n505), .ZN(G1330GAT) );
  NOR2_X1 U572 ( .A1(n529), .A2(n506), .ZN(n507) );
  XOR2_X1 U573 ( .A(G50GAT), .B(n507), .Z(G1331GAT) );
  NOR2_X1 U574 ( .A1(n509), .A2(n508), .ZN(n510) );
  XOR2_X1 U575 ( .A(KEYINPUT108), .B(n510), .Z(n517) );
  NOR2_X1 U576 ( .A1(n517), .A2(n520), .ZN(n511) );
  XOR2_X1 U577 ( .A(KEYINPUT42), .B(n511), .Z(n512) );
  XNOR2_X1 U578 ( .A(G57GAT), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U579 ( .A1(n513), .A2(n517), .ZN(n514) );
  XOR2_X1 U580 ( .A(G64GAT), .B(n514), .Z(G1333GAT) );
  NOR2_X1 U581 ( .A1(n517), .A2(n562), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(G1334GAT) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n519) );
  NOR2_X1 U585 ( .A1(n529), .A2(n517), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NOR2_X1 U587 ( .A1(n523), .A2(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(G1336GAT) );
  NOR2_X1 U590 ( .A1(n523), .A2(n562), .ZN(n524) );
  XOR2_X1 U591 ( .A(G99GAT), .B(n524), .Z(G1338GAT) );
  INV_X1 U592 ( .A(n525), .ZN(n526) );
  NOR2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n545) );
  NAND2_X1 U594 ( .A1(n408), .A2(n545), .ZN(n528) );
  XNOR2_X1 U595 ( .A(KEYINPUT115), .B(n528), .ZN(n530) );
  NAND2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n539) );
  NOR2_X1 U597 ( .A1(n531), .A2(n539), .ZN(n532) );
  XOR2_X1 U598 ( .A(G113GAT), .B(n532), .Z(G1340GAT) );
  NOR2_X1 U599 ( .A1(n550), .A2(n539), .ZN(n534) );
  XNOR2_X1 U600 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U602 ( .A(G120GAT), .B(n535), .ZN(G1341GAT) );
  INV_X1 U603 ( .A(n539), .ZN(n536) );
  NAND2_X1 U604 ( .A1(n571), .A2(n536), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n537), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  NOR2_X1 U607 ( .A1(n539), .A2(n556), .ZN(n543) );
  XOR2_X1 U608 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n541) );
  XNOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT118), .ZN(n540) );
  XNOR2_X1 U610 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  NAND2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n555) );
  NOR2_X1 U613 ( .A1(n577), .A2(n555), .ZN(n547) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n549) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n548) );
  XNOR2_X1 U618 ( .A(n549), .B(n548), .ZN(n552) );
  NOR2_X1 U619 ( .A1(n550), .A2(n555), .ZN(n551) );
  XOR2_X1 U620 ( .A(n552), .B(n551), .Z(G1345GAT) );
  NOR2_X1 U621 ( .A1(n582), .A2(n555), .ZN(n554) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n553) );
  XNOR2_X1 U623 ( .A(n554), .B(n553), .ZN(G1346GAT) );
  NOR2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U625 ( .A(G162GAT), .B(n557), .Z(G1347GAT) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n561) );
  INV_X1 U627 ( .A(KEYINPUT55), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n566) );
  NOR2_X1 U629 ( .A1(n562), .A2(n566), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n563), .A2(n573), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  OR2_X1 U632 ( .A1(n296), .A2(n566), .ZN(n568) );
  XOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT123), .Z(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n570) );
  XOR2_X1 U635 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1349GAT) );
  NAND2_X1 U637 ( .A1(n571), .A2(n573), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U639 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1351GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n584), .ZN(n581) );
  XOR2_X1 U643 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  OR2_X1 U647 ( .A1(n584), .A2(n582), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n587) );
  NOR2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

