

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729;

  XNOR2_X1 U371 ( .A(n355), .B(KEYINPUT84), .ZN(n592) );
  AND2_X2 U372 ( .A1(n535), .A2(n531), .ZN(n419) );
  NOR2_X2 U373 ( .A1(n649), .A2(n565), .ZN(n509) );
  OR2_X2 U374 ( .A1(n512), .A2(n653), .ZN(n381) );
  XNOR2_X2 U375 ( .A(n431), .B(n421), .ZN(n473) );
  XNOR2_X2 U376 ( .A(n420), .B(G128), .ZN(n431) );
  NOR2_X2 U377 ( .A1(n666), .A2(n518), .ZN(n519) );
  NAND2_X1 U378 ( .A1(n713), .A2(KEYINPUT2), .ZN(n355) );
  XNOR2_X1 U379 ( .A(n401), .B(KEYINPUT114), .ZN(n568) );
  OR2_X1 U380 ( .A1(n564), .A2(n565), .ZN(n401) );
  XNOR2_X1 U381 ( .A(n502), .B(n501), .ZN(n646) );
  XNOR2_X1 U382 ( .A(n608), .B(n607), .ZN(n609) );
  XNOR2_X1 U383 ( .A(KEYINPUT85), .B(KEYINPUT48), .ZN(n581) );
  INV_X1 U384 ( .A(G143), .ZN(n420) );
  INV_X2 U385 ( .A(G953), .ZN(n714) );
  XNOR2_X2 U386 ( .A(KEYINPUT38), .B(n588), .ZN(n637) );
  INV_X2 U387 ( .A(G146), .ZN(n391) );
  NOR2_X1 U388 ( .A1(G902), .A2(n684), .ZN(n485) );
  XNOR2_X2 U389 ( .A(n553), .B(KEYINPUT115), .ZN(n723) );
  XNOR2_X2 U390 ( .A(n463), .B(n390), .ZN(n492) );
  XNOR2_X2 U391 ( .A(n391), .B(G125), .ZN(n463) );
  XNOR2_X1 U392 ( .A(n640), .B(n383), .ZN(n569) );
  INV_X1 U393 ( .A(G134), .ZN(n421) );
  INV_X1 U394 ( .A(KEYINPUT10), .ZN(n390) );
  NOR2_X1 U395 ( .A1(G902), .A2(n606), .ZN(n428) );
  XNOR2_X1 U396 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n474) );
  XNOR2_X1 U397 ( .A(n479), .B(n478), .ZN(n520) );
  NAND2_X1 U398 ( .A1(n381), .A2(n380), .ZN(n379) );
  NOR2_X1 U399 ( .A1(G953), .A2(G237), .ZN(n459) );
  XOR2_X1 U400 ( .A(KEYINPUT67), .B(G140), .Z(n493) );
  XNOR2_X1 U401 ( .A(n463), .B(n359), .ZN(n432) );
  XNOR2_X1 U402 ( .A(n430), .B(n429), .ZN(n359) );
  XNOR2_X1 U403 ( .A(n431), .B(n394), .ZN(n393) );
  XNOR2_X1 U404 ( .A(n395), .B(KEYINPUT18), .ZN(n394) );
  INV_X1 U405 ( .A(KEYINPUT17), .ZN(n395) );
  XNOR2_X1 U406 ( .A(n697), .B(KEYINPUT69), .ZN(n484) );
  XNOR2_X1 U407 ( .A(KEYINPUT66), .B(KEYINPUT0), .ZN(n455) );
  INV_X1 U408 ( .A(n506), .ZN(n521) );
  XNOR2_X1 U409 ( .A(n492), .B(n493), .ZN(n711) );
  XNOR2_X1 U410 ( .A(G137), .B(G119), .ZN(n487) );
  XNOR2_X1 U411 ( .A(n352), .B(n462), .ZN(n466) );
  NOR2_X1 U412 ( .A1(n614), .A2(n561), .ZN(n548) );
  XNOR2_X1 U413 ( .A(n443), .B(n442), .ZN(n444) );
  INV_X1 U414 ( .A(KEYINPUT65), .ZN(n486) );
  BUF_X1 U415 ( .A(n646), .Z(n360) );
  XNOR2_X1 U416 ( .A(n472), .B(n365), .ZN(n477) );
  XNOR2_X1 U417 ( .A(n678), .B(KEYINPUT54), .ZN(n679) );
  XNOR2_X1 U418 ( .A(n400), .B(KEYINPUT47), .ZN(n571) );
  XNOR2_X1 U419 ( .A(n458), .B(n457), .ZN(n497) );
  XNOR2_X1 U420 ( .A(KEYINPUT96), .B(KEYINPUT20), .ZN(n457) );
  XNOR2_X1 U421 ( .A(n507), .B(n367), .ZN(n640) );
  INV_X1 U422 ( .A(KEYINPUT110), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n403), .B(n402), .ZN(n645) );
  XNOR2_X1 U424 ( .A(KEYINPUT98), .B(KEYINPUT21), .ZN(n402) );
  NAND2_X1 U425 ( .A1(n497), .A2(G221), .ZN(n403) );
  INV_X1 U426 ( .A(KEYINPUT5), .ZN(n362) );
  XNOR2_X1 U427 ( .A(G101), .B(G113), .ZN(n423) );
  XOR2_X1 U428 ( .A(KEYINPUT101), .B(G116), .Z(n424) );
  XNOR2_X1 U429 ( .A(n473), .B(n417), .ZN(n710) );
  XNOR2_X1 U430 ( .A(n422), .B(KEYINPUT4), .ZN(n417) );
  XNOR2_X1 U431 ( .A(G131), .B(G137), .ZN(n422) );
  XOR2_X1 U432 ( .A(KEYINPUT3), .B(G119), .Z(n439) );
  XOR2_X1 U433 ( .A(G122), .B(G140), .Z(n461) );
  XNOR2_X1 U434 ( .A(G131), .B(G143), .ZN(n460) );
  XNOR2_X1 U435 ( .A(n368), .B(n405), .ZN(n352) );
  XNOR2_X1 U436 ( .A(n404), .B(KEYINPUT103), .ZN(n368) );
  XNOR2_X1 U437 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n404) );
  XOR2_X1 U438 ( .A(G113), .B(G104), .Z(n464) );
  XNOR2_X1 U439 ( .A(n493), .B(n418), .ZN(n482) );
  XNOR2_X1 U440 ( .A(n710), .B(G146), .ZN(n483) );
  OR2_X1 U441 ( .A1(G237), .A2(G902), .ZN(n446) );
  NAND2_X1 U442 ( .A1(n521), .A2(n520), .ZN(n639) );
  NOR2_X1 U443 ( .A1(n639), .A2(n645), .ZN(n411) );
  OR2_X2 U444 ( .A1(n646), .A2(n645), .ZN(n649) );
  XNOR2_X1 U445 ( .A(n483), .B(n374), .ZN(n606) );
  XNOR2_X1 U446 ( .A(n427), .B(n439), .ZN(n374) );
  XNOR2_X1 U447 ( .A(n425), .B(n361), .ZN(n427) );
  XNOR2_X1 U448 ( .A(n426), .B(n362), .ZN(n361) );
  XNOR2_X1 U449 ( .A(n473), .B(n348), .ZN(n365) );
  XNOR2_X1 U450 ( .A(n483), .B(n384), .ZN(n684) );
  XNOR2_X1 U451 ( .A(n484), .B(n385), .ZN(n384) );
  XNOR2_X1 U452 ( .A(n482), .B(n386), .ZN(n385) );
  XNOR2_X1 U453 ( .A(n617), .B(G104), .ZN(n386) );
  XNOR2_X1 U454 ( .A(n376), .B(n441), .ZN(n677) );
  XNOR2_X1 U455 ( .A(n696), .B(KEYINPUT4), .ZN(n376) );
  XNOR2_X1 U456 ( .A(n432), .B(n393), .ZN(n434) );
  BUF_X1 U457 ( .A(n593), .Z(n705) );
  NOR2_X1 U458 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U459 ( .A(n468), .B(G475), .ZN(n506) );
  XNOR2_X1 U460 ( .A(n369), .B(n467), .ZN(n468) );
  INV_X1 U461 ( .A(KEYINPUT100), .ZN(n510) );
  XNOR2_X1 U462 ( .A(G128), .B(G110), .ZN(n490) );
  XNOR2_X1 U463 ( .A(n599), .B(KEYINPUT59), .ZN(n600) );
  NOR2_X1 U464 ( .A1(n550), .A2(n584), .ZN(n551) );
  XNOR2_X1 U465 ( .A(n529), .B(n354), .ZN(n725) );
  XNOR2_X1 U466 ( .A(n530), .B(KEYINPUT75), .ZN(n354) );
  INV_X1 U467 ( .A(n400), .ZN(n625) );
  NOR2_X1 U468 ( .A1(n506), .A2(n520), .ZN(n630) );
  INV_X1 U469 ( .A(KEYINPUT113), .ZN(n406) );
  INV_X1 U470 ( .A(G107), .ZN(n617) );
  XNOR2_X1 U471 ( .A(n689), .B(n690), .ZN(n353) );
  INV_X1 U472 ( .A(KEYINPUT56), .ZN(n415) );
  NOR2_X1 U473 ( .A1(n675), .A2(G953), .ZN(n412) );
  NAND2_X1 U474 ( .A1(n673), .A2(n414), .ZN(n413) );
  XNOR2_X1 U475 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n348) );
  AND2_X1 U476 ( .A1(n494), .A2(G221), .ZN(n349) );
  NOR2_X1 U477 ( .A1(n713), .A2(KEYINPUT2), .ZN(n350) );
  XNOR2_X1 U478 ( .A(G902), .B(KEYINPUT15), .ZN(n594) );
  INV_X1 U479 ( .A(n594), .ZN(n595) );
  XOR2_X1 U480 ( .A(n686), .B(n685), .Z(n351) );
  XOR2_X1 U481 ( .A(KEYINPUT90), .B(n602), .Z(n683) );
  XNOR2_X1 U482 ( .A(n519), .B(KEYINPUT34), .ZN(n522) );
  XNOR2_X2 U483 ( .A(KEYINPUT35), .B(n523), .ZN(n726) );
  NAND2_X1 U484 ( .A1(n382), .A2(n379), .ZN(n378) );
  XNOR2_X1 U485 ( .A(n711), .B(n349), .ZN(n495) );
  NOR2_X1 U486 ( .A1(n353), .A2(n695), .ZN(G63) );
  AND2_X1 U487 ( .A1(n356), .A2(n683), .ZN(G54) );
  XNOR2_X1 U488 ( .A(n688), .B(n351), .ZN(n356) );
  NOR2_X2 U489 ( .A1(n593), .A2(n592), .ZN(n674) );
  NOR2_X1 U490 ( .A1(n599), .A2(G902), .ZN(n369) );
  NAND2_X1 U491 ( .A1(n371), .A2(n572), .ZN(n370) );
  NOR2_X2 U492 ( .A1(n357), .A2(n674), .ZN(n687) );
  NOR2_X1 U493 ( .A1(n598), .A2(n597), .ZN(n357) );
  XNOR2_X1 U494 ( .A(n550), .B(n447), .ZN(n392) );
  INV_X1 U495 ( .A(G101), .ZN(n375) );
  XNOR2_X1 U496 ( .A(n375), .B(G110), .ZN(n433) );
  XNOR2_X1 U497 ( .A(n358), .B(KEYINPUT39), .ZN(n582) );
  NOR2_X2 U498 ( .A1(n372), .A2(n558), .ZN(n358) );
  NOR2_X2 U499 ( .A1(n726), .A2(n725), .ZN(n535) );
  XNOR2_X2 U500 ( .A(n539), .B(KEYINPUT45), .ZN(n593) );
  INV_X1 U501 ( .A(n387), .ZN(n371) );
  XNOR2_X1 U502 ( .A(n509), .B(KEYINPUT99), .ZN(n387) );
  NOR2_X1 U503 ( .A1(n558), .A2(n370), .ZN(n573) );
  AND2_X2 U504 ( .A1(n515), .A2(n549), .ZN(n517) );
  NAND2_X1 U505 ( .A1(n363), .A2(n533), .ZN(n534) );
  NAND2_X1 U506 ( .A1(n419), .A2(n727), .ZN(n363) );
  NAND2_X1 U507 ( .A1(n527), .A2(n528), .ZN(n529) );
  XNOR2_X1 U508 ( .A(n411), .B(KEYINPUT112), .ZN(n410) );
  XNOR2_X2 U509 ( .A(n364), .B(G122), .ZN(n471) );
  XNOR2_X2 U510 ( .A(G116), .B(G107), .ZN(n364) );
  NOR2_X2 U511 ( .A1(n503), .A2(n653), .ZN(n409) );
  XNOR2_X1 U512 ( .A(n409), .B(n486), .ZN(n408) );
  NAND2_X1 U513 ( .A1(n579), .A2(n366), .ZN(n399) );
  XNOR2_X1 U514 ( .A(n577), .B(n578), .ZN(n366) );
  NAND2_X1 U515 ( .A1(n640), .A2(KEYINPUT47), .ZN(n575) );
  XNOR2_X1 U516 ( .A(n630), .B(KEYINPUT109), .ZN(n583) );
  INV_X1 U517 ( .A(n637), .ZN(n373) );
  OR2_X2 U518 ( .A1(n373), .A2(n387), .ZN(n372) );
  XNOR2_X2 U519 ( .A(n377), .B(n440), .ZN(n696) );
  NAND2_X1 U520 ( .A1(n438), .A2(n437), .ZN(n377) );
  INV_X1 U521 ( .A(n381), .ZN(n618) );
  NAND2_X1 U522 ( .A1(n613), .A2(n378), .ZN(n532) );
  INV_X1 U523 ( .A(n629), .ZN(n380) );
  INV_X1 U524 ( .A(n569), .ZN(n382) );
  INV_X1 U525 ( .A(KEYINPUT79), .ZN(n383) );
  NOR2_X1 U526 ( .A1(n387), .A2(n518), .ZN(n511) );
  NAND2_X1 U527 ( .A1(n388), .A2(n567), .ZN(n580) );
  XNOR2_X1 U528 ( .A(n389), .B(KEYINPUT46), .ZN(n388) );
  NOR2_X2 U529 ( .A1(n729), .A2(n728), .ZN(n389) );
  XNOR2_X1 U530 ( .A(n559), .B(KEYINPUT40), .ZN(n729) );
  NOR2_X2 U531 ( .A1(n392), .A2(n454), .ZN(n456) );
  OR2_X1 U532 ( .A1(n568), .A2(n392), .ZN(n400) );
  NOR2_X2 U533 ( .A1(n677), .A2(n595), .ZN(n445) );
  XNOR2_X1 U534 ( .A(n396), .B(n581), .ZN(n591) );
  NOR2_X1 U535 ( .A1(n580), .A2(n397), .ZN(n396) );
  XNOR2_X1 U536 ( .A(n399), .B(n398), .ZN(n397) );
  INV_X1 U537 ( .A(KEYINPUT71), .ZN(n398) );
  XNOR2_X1 U538 ( .A(n682), .B(n415), .ZN(G51) );
  NAND2_X1 U539 ( .A1(n459), .A2(G214), .ZN(n405) );
  XNOR2_X2 U540 ( .A(n407), .B(n406), .ZN(n727) );
  NAND2_X1 U541 ( .A1(n408), .A2(n360), .ZN(n407) );
  NAND2_X1 U542 ( .A1(n508), .A2(n410), .ZN(n481) );
  NAND2_X1 U543 ( .A1(n413), .A2(n412), .ZN(n676) );
  NOR2_X1 U544 ( .A1(n674), .A2(n350), .ZN(n414) );
  NOR2_X1 U545 ( .A1(n593), .A2(n416), .ZN(n598) );
  NAND2_X1 U546 ( .A1(n713), .A2(n595), .ZN(n416) );
  XNOR2_X1 U547 ( .A(n466), .B(n465), .ZN(n599) );
  NOR2_X2 U548 ( .A1(n591), .A2(n590), .ZN(n713) );
  XNOR2_X2 U549 ( .A(n428), .B(G472), .ZN(n562) );
  AND2_X1 U550 ( .A1(G227), .A2(n714), .ZN(n418) );
  INV_X1 U551 ( .A(KEYINPUT74), .ZN(n429) );
  INV_X1 U552 ( .A(KEYINPUT62), .ZN(n607) );
  INV_X1 U553 ( .A(KEYINPUT77), .ZN(n442) );
  INV_X1 U554 ( .A(KEYINPUT19), .ZN(n447) );
  XNOR2_X1 U555 ( .A(n610), .B(n609), .ZN(n611) );
  INV_X1 U556 ( .A(KEYINPUT60), .ZN(n604) );
  XNOR2_X1 U557 ( .A(n605), .B(n604), .ZN(G60) );
  XNOR2_X1 U558 ( .A(n424), .B(n423), .ZN(n425) );
  NAND2_X1 U559 ( .A1(n459), .A2(G210), .ZN(n426) );
  INV_X1 U560 ( .A(n562), .ZN(n653) );
  NAND2_X1 U561 ( .A1(G224), .A2(n714), .ZN(n430) );
  XNOR2_X1 U562 ( .A(KEYINPUT91), .B(n433), .ZN(n697) );
  XNOR2_X1 U563 ( .A(n484), .B(n434), .ZN(n441) );
  INV_X1 U564 ( .A(n471), .ZN(n435) );
  NAND2_X1 U565 ( .A1(n435), .A2(n464), .ZN(n438) );
  INV_X1 U566 ( .A(n464), .ZN(n436) );
  NAND2_X1 U567 ( .A1(n471), .A2(n436), .ZN(n437) );
  XNOR2_X1 U568 ( .A(n439), .B(KEYINPUT16), .ZN(n440) );
  NAND2_X1 U569 ( .A1(G210), .A2(n446), .ZN(n443) );
  XNOR2_X2 U570 ( .A(n445), .B(n444), .ZN(n574) );
  NAND2_X1 U571 ( .A1(G214), .A2(n446), .ZN(n636) );
  NAND2_X1 U572 ( .A1(n574), .A2(n636), .ZN(n550) );
  NAND2_X1 U573 ( .A1(G234), .A2(G237), .ZN(n448) );
  XNOR2_X1 U574 ( .A(n448), .B(KEYINPUT14), .ZN(n449) );
  XNOR2_X1 U575 ( .A(KEYINPUT72), .B(n449), .ZN(n452) );
  NAND2_X1 U576 ( .A1(G952), .A2(n452), .ZN(n664) );
  NOR2_X1 U577 ( .A1(G953), .A2(n664), .ZN(n450) );
  XNOR2_X1 U578 ( .A(KEYINPUT92), .B(n450), .ZN(n540) );
  XNOR2_X1 U579 ( .A(G898), .B(KEYINPUT93), .ZN(n704) );
  NAND2_X1 U580 ( .A1(n704), .A2(G953), .ZN(n451) );
  XNOR2_X1 U581 ( .A(n451), .B(KEYINPUT94), .ZN(n699) );
  NAND2_X1 U582 ( .A1(G902), .A2(n452), .ZN(n541) );
  NOR2_X1 U583 ( .A1(n699), .A2(n541), .ZN(n453) );
  NOR2_X1 U584 ( .A1(n540), .A2(n453), .ZN(n454) );
  XNOR2_X1 U585 ( .A(n456), .B(n455), .ZN(n508) );
  NAND2_X1 U586 ( .A1(n594), .A2(G234), .ZN(n458) );
  XNOR2_X1 U587 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U588 ( .A(n492), .B(n464), .ZN(n465) );
  XNOR2_X1 U589 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n467) );
  XNOR2_X1 U590 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n469) );
  XNOR2_X1 U591 ( .A(n469), .B(KEYINPUT107), .ZN(n470) );
  XNOR2_X1 U592 ( .A(n471), .B(n470), .ZN(n472) );
  NAND2_X1 U593 ( .A1(n714), .A2(G234), .ZN(n475) );
  XNOR2_X1 U594 ( .A(n475), .B(n474), .ZN(n494) );
  NAND2_X1 U595 ( .A1(G217), .A2(n494), .ZN(n476) );
  XNOR2_X1 U596 ( .A(n477), .B(n476), .ZN(n690) );
  NOR2_X1 U597 ( .A1(G902), .A2(n690), .ZN(n479) );
  XNOR2_X1 U598 ( .A(KEYINPUT108), .B(G478), .ZN(n478) );
  XOR2_X1 U599 ( .A(KEYINPUT22), .B(KEYINPUT70), .Z(n480) );
  XNOR2_X2 U600 ( .A(n481), .B(n480), .ZN(n527) );
  XNOR2_X2 U601 ( .A(G469), .B(n485), .ZN(n565) );
  XNOR2_X2 U602 ( .A(n565), .B(KEYINPUT1), .ZN(n648) );
  NAND2_X1 U603 ( .A1(n527), .A2(n648), .ZN(n503) );
  XOR2_X1 U604 ( .A(KEYINPUT23), .B(KEYINPUT95), .Z(n488) );
  XNOR2_X1 U605 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U606 ( .A(n489), .B(KEYINPUT24), .Z(n491) );
  XNOR2_X1 U607 ( .A(n491), .B(n490), .ZN(n496) );
  XNOR2_X1 U608 ( .A(n495), .B(n496), .ZN(n693) );
  NOR2_X1 U609 ( .A1(G902), .A2(n693), .ZN(n502) );
  XOR2_X1 U610 ( .A(KEYINPUT97), .B(KEYINPUT73), .Z(n499) );
  NAND2_X1 U611 ( .A1(G217), .A2(n497), .ZN(n498) );
  XNOR2_X1 U612 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U613 ( .A(KEYINPUT25), .B(n500), .ZN(n501) );
  NOR2_X1 U614 ( .A1(n360), .A2(n503), .ZN(n505) );
  XNOR2_X1 U615 ( .A(KEYINPUT6), .B(KEYINPUT111), .ZN(n504) );
  XOR2_X1 U616 ( .A(n504), .B(n562), .Z(n549) );
  INV_X1 U617 ( .A(n549), .ZN(n524) );
  NAND2_X1 U618 ( .A1(n505), .A2(n524), .ZN(n613) );
  NAND2_X1 U619 ( .A1(n520), .A2(n506), .ZN(n614) );
  NAND2_X1 U620 ( .A1(n583), .A2(n614), .ZN(n507) );
  INV_X1 U621 ( .A(n508), .ZN(n518) );
  XNOR2_X1 U622 ( .A(n511), .B(n510), .ZN(n512) );
  NOR2_X1 U623 ( .A1(n649), .A2(n648), .ZN(n515) );
  NAND2_X1 U624 ( .A1(n653), .A2(n515), .ZN(n657) );
  NOR2_X1 U625 ( .A1(n518), .A2(n657), .ZN(n514) );
  XOR2_X1 U626 ( .A(KEYINPUT102), .B(KEYINPUT31), .Z(n513) );
  XNOR2_X1 U627 ( .A(n514), .B(n513), .ZN(n629) );
  INV_X1 U628 ( .A(n532), .ZN(n531) );
  XNOR2_X1 U629 ( .A(KEYINPUT88), .B(KEYINPUT33), .ZN(n516) );
  XNOR2_X2 U630 ( .A(n517), .B(n516), .ZN(n666) );
  NOR2_X1 U631 ( .A1(n521), .A2(n520), .ZN(n572) );
  NAND2_X1 U632 ( .A1(n522), .A2(n572), .ZN(n523) );
  XNOR2_X1 U633 ( .A(KEYINPUT64), .B(KEYINPUT32), .ZN(n530) );
  NAND2_X1 U634 ( .A1(n360), .A2(n524), .ZN(n525) );
  NOR2_X1 U635 ( .A1(n648), .A2(n525), .ZN(n526) );
  XNOR2_X1 U636 ( .A(KEYINPUT76), .B(n526), .ZN(n528) );
  OR2_X1 U637 ( .A1(n532), .A2(KEYINPUT44), .ZN(n533) );
  XNOR2_X1 U638 ( .A(n534), .B(KEYINPUT87), .ZN(n538) );
  NAND2_X1 U639 ( .A1(n535), .A2(n727), .ZN(n536) );
  NOR2_X1 U640 ( .A1(n536), .A2(KEYINPUT44), .ZN(n537) );
  NOR2_X2 U641 ( .A1(n538), .A2(n537), .ZN(n539) );
  INV_X1 U642 ( .A(n645), .ZN(n545) );
  INV_X1 U643 ( .A(n540), .ZN(n544) );
  NOR2_X1 U644 ( .A1(G900), .A2(n541), .ZN(n542) );
  NAND2_X1 U645 ( .A1(G953), .A2(n542), .ZN(n543) );
  NAND2_X1 U646 ( .A1(n544), .A2(n543), .ZN(n556) );
  NAND2_X1 U647 ( .A1(n545), .A2(n556), .ZN(n546) );
  XOR2_X1 U648 ( .A(KEYINPUT68), .B(n546), .Z(n547) );
  NAND2_X1 U649 ( .A1(n646), .A2(n547), .ZN(n561) );
  NAND2_X1 U650 ( .A1(n549), .A2(n548), .ZN(n584) );
  XNOR2_X1 U651 ( .A(KEYINPUT36), .B(n551), .ZN(n552) );
  INV_X1 U652 ( .A(n648), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n552), .A2(n585), .ZN(n553) );
  XOR2_X1 U654 ( .A(n723), .B(KEYINPUT86), .Z(n567) );
  INV_X1 U655 ( .A(n636), .ZN(n554) );
  OR2_X1 U656 ( .A1(n562), .A2(n554), .ZN(n555) );
  XOR2_X1 U657 ( .A(KEYINPUT30), .B(n555), .Z(n557) );
  NAND2_X1 U658 ( .A1(n557), .A2(n556), .ZN(n558) );
  INV_X1 U659 ( .A(n574), .ZN(n588) );
  NOR2_X1 U660 ( .A1(n582), .A2(n614), .ZN(n559) );
  NAND2_X1 U661 ( .A1(n637), .A2(n636), .ZN(n641) );
  NOR2_X1 U662 ( .A1(n641), .A2(n639), .ZN(n560) );
  XNOR2_X1 U663 ( .A(n560), .B(KEYINPUT41), .ZN(n667) );
  XOR2_X1 U664 ( .A(KEYINPUT28), .B(n563), .Z(n564) );
  NOR2_X1 U665 ( .A1(n667), .A2(n568), .ZN(n566) );
  XNOR2_X1 U666 ( .A(n566), .B(KEYINPUT42), .ZN(n728) );
  NAND2_X1 U667 ( .A1(n625), .A2(n569), .ZN(n570) );
  NAND2_X1 U668 ( .A1(n571), .A2(n570), .ZN(n579) );
  INV_X1 U669 ( .A(KEYINPUT78), .ZN(n578) );
  NAND2_X1 U670 ( .A1(n574), .A2(n573), .ZN(n624) );
  XNOR2_X1 U671 ( .A(n624), .B(KEYINPUT80), .ZN(n576) );
  NAND2_X1 U672 ( .A1(n576), .A2(n575), .ZN(n577) );
  OR2_X1 U673 ( .A1(n583), .A2(n582), .ZN(n633) );
  NOR2_X1 U674 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U675 ( .A1(n586), .A2(n636), .ZN(n587) );
  XNOR2_X1 U676 ( .A(n587), .B(KEYINPUT43), .ZN(n589) );
  NAND2_X1 U677 ( .A1(n589), .A2(n588), .ZN(n635) );
  NAND2_X1 U678 ( .A1(n633), .A2(n635), .ZN(n590) );
  INV_X1 U679 ( .A(KEYINPUT2), .ZN(n671) );
  XNOR2_X1 U680 ( .A(KEYINPUT83), .B(n595), .ZN(n596) );
  NOR2_X1 U681 ( .A1(n671), .A2(n596), .ZN(n597) );
  NAND2_X1 U682 ( .A1(G475), .A2(n687), .ZN(n601) );
  XNOR2_X1 U683 ( .A(n601), .B(n600), .ZN(n603) );
  NOR2_X1 U684 ( .A1(G952), .A2(n714), .ZN(n602) );
  NAND2_X1 U685 ( .A1(n603), .A2(n683), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n687), .A2(G472), .ZN(n610) );
  XOR2_X1 U687 ( .A(n606), .B(KEYINPUT89), .Z(n608) );
  NAND2_X1 U688 ( .A1(n611), .A2(n683), .ZN(n612) );
  XNOR2_X1 U689 ( .A(n612), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U690 ( .A(G101), .B(n613), .ZN(G3) );
  XNOR2_X1 U691 ( .A(G104), .B(KEYINPUT116), .ZN(n616) );
  INV_X1 U692 ( .A(n614), .ZN(n627) );
  NAND2_X1 U693 ( .A1(n627), .A2(n618), .ZN(n615) );
  XNOR2_X1 U694 ( .A(n616), .B(n615), .ZN(G6) );
  XOR2_X1 U695 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n620) );
  NAND2_X1 U696 ( .A1(n618), .A2(n630), .ZN(n619) );
  XNOR2_X1 U697 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U698 ( .A(G107), .B(n621), .ZN(G9) );
  XOR2_X1 U699 ( .A(G128), .B(KEYINPUT29), .Z(n623) );
  NAND2_X1 U700 ( .A1(n625), .A2(n630), .ZN(n622) );
  XNOR2_X1 U701 ( .A(n623), .B(n622), .ZN(G30) );
  XNOR2_X1 U702 ( .A(n624), .B(G143), .ZN(G45) );
  NAND2_X1 U703 ( .A1(n625), .A2(n627), .ZN(n626) );
  XNOR2_X1 U704 ( .A(n626), .B(G146), .ZN(G48) );
  NAND2_X1 U705 ( .A1(n629), .A2(n627), .ZN(n628) );
  XNOR2_X1 U706 ( .A(n628), .B(G113), .ZN(G15) );
  XOR2_X1 U707 ( .A(G116), .B(KEYINPUT117), .Z(n632) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U709 ( .A(n632), .B(n631), .ZN(G18) );
  XNOR2_X1 U710 ( .A(G134), .B(KEYINPUT118), .ZN(n634) );
  XNOR2_X1 U711 ( .A(n634), .B(n633), .ZN(G36) );
  XNOR2_X1 U712 ( .A(G140), .B(n635), .ZN(G42) );
  NOR2_X1 U713 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n643) );
  NOR2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U716 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U717 ( .A1(n666), .A2(n644), .ZN(n661) );
  NAND2_X1 U718 ( .A1(n360), .A2(n645), .ZN(n647) );
  XOR2_X1 U719 ( .A(KEYINPUT49), .B(n647), .Z(n655) );
  NAND2_X1 U720 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U721 ( .A(n650), .B(KEYINPUT119), .ZN(n651) );
  XNOR2_X1 U722 ( .A(KEYINPUT50), .B(n651), .ZN(n652) );
  NOR2_X1 U723 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U724 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U726 ( .A(KEYINPUT51), .B(n658), .ZN(n659) );
  NOR2_X1 U727 ( .A1(n659), .A2(n667), .ZN(n660) );
  NOR2_X1 U728 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U729 ( .A(n662), .B(KEYINPUT52), .ZN(n663) );
  NOR2_X1 U730 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U731 ( .A(n665), .B(KEYINPUT120), .ZN(n669) );
  NOR2_X1 U732 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U733 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U734 ( .A(n670), .B(KEYINPUT121), .ZN(n675) );
  NAND2_X1 U735 ( .A1(n705), .A2(n671), .ZN(n672) );
  XNOR2_X1 U736 ( .A(n672), .B(KEYINPUT82), .ZN(n673) );
  XOR2_X1 U737 ( .A(KEYINPUT53), .B(n676), .Z(G75) );
  NAND2_X1 U738 ( .A1(G210), .A2(n687), .ZN(n680) );
  XNOR2_X1 U739 ( .A(n677), .B(KEYINPUT55), .ZN(n678) );
  XNOR2_X1 U740 ( .A(n680), .B(n679), .ZN(n681) );
  NAND2_X1 U741 ( .A1(n681), .A2(n683), .ZN(n682) );
  INV_X1 U742 ( .A(n683), .ZN(n695) );
  XOR2_X1 U743 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n686) );
  XNOR2_X1 U744 ( .A(n684), .B(KEYINPUT122), .ZN(n685) );
  BUF_X2 U745 ( .A(n687), .Z(n691) );
  NAND2_X1 U746 ( .A1(n691), .A2(G469), .ZN(n688) );
  NAND2_X1 U747 ( .A1(G478), .A2(n691), .ZN(n689) );
  NAND2_X1 U748 ( .A1(G217), .A2(n691), .ZN(n692) );
  XNOR2_X1 U749 ( .A(n692), .B(n693), .ZN(n694) );
  NOR2_X1 U750 ( .A1(n695), .A2(n694), .ZN(G66) );
  XNOR2_X1 U751 ( .A(n696), .B(KEYINPUT124), .ZN(n698) );
  XNOR2_X1 U752 ( .A(n698), .B(n697), .ZN(n700) );
  NAND2_X1 U753 ( .A1(n700), .A2(n699), .ZN(n709) );
  NAND2_X1 U754 ( .A1(G224), .A2(G953), .ZN(n701) );
  XNOR2_X1 U755 ( .A(n701), .B(KEYINPUT123), .ZN(n702) );
  XNOR2_X1 U756 ( .A(n702), .B(KEYINPUT61), .ZN(n703) );
  NOR2_X1 U757 ( .A1(n704), .A2(n703), .ZN(n707) );
  NOR2_X1 U758 ( .A1(G953), .A2(n705), .ZN(n706) );
  NOR2_X1 U759 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U760 ( .A(n709), .B(n708), .ZN(G69) );
  XNOR2_X1 U761 ( .A(KEYINPUT125), .B(n710), .ZN(n712) );
  XNOR2_X1 U762 ( .A(n711), .B(n712), .ZN(n716) );
  XOR2_X1 U763 ( .A(n713), .B(n716), .Z(n715) );
  NAND2_X1 U764 ( .A1(n715), .A2(n714), .ZN(n722) );
  XNOR2_X1 U765 ( .A(n716), .B(KEYINPUT126), .ZN(n717) );
  XNOR2_X1 U766 ( .A(G227), .B(n717), .ZN(n718) );
  NAND2_X1 U767 ( .A1(G900), .A2(n718), .ZN(n719) );
  NAND2_X1 U768 ( .A1(G953), .A2(n719), .ZN(n720) );
  XOR2_X1 U769 ( .A(KEYINPUT127), .B(n720), .Z(n721) );
  NAND2_X1 U770 ( .A1(n722), .A2(n721), .ZN(G72) );
  XNOR2_X1 U771 ( .A(G125), .B(n723), .ZN(n724) );
  XNOR2_X1 U772 ( .A(n724), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U773 ( .A(n725), .B(G119), .Z(G21) );
  XOR2_X1 U774 ( .A(G122), .B(n726), .Z(G24) );
  XNOR2_X1 U775 ( .A(G110), .B(n727), .ZN(G12) );
  XOR2_X1 U776 ( .A(G137), .B(n728), .Z(G39) );
  XOR2_X1 U777 ( .A(n729), .B(G131), .Z(G33) );
endmodule

