//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960;
  INV_X1    g000(.A(KEYINPUT22), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(KEYINPUT71), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(KEYINPUT71), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G169gat), .ZN(new_n212));
  INV_X1    g011(.A(G176gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT26), .ZN(new_n214));
  INV_X1    g013(.A(G183gat), .ZN(new_n215));
  INV_X1    g014(.A(G190gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n212), .A2(new_n213), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT26), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(G169gat), .B2(G176gat), .ZN(new_n219));
  OAI221_X1 g018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT27), .B(G183gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(new_n216), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT67), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT28), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n220), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n222), .B(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(new_n224), .A3(new_n225), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT25), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT23), .B1(new_n212), .B2(new_n213), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT64), .B(G176gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n212), .A2(KEYINPUT23), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(new_n215), .B2(new_n216), .ZN(new_n238));
  NAND3_X1  g037(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n231), .B1(new_n236), .B2(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n239), .B(KEYINPUT65), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n238), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT23), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n243), .A2(KEYINPUT25), .A3(new_n233), .A4(new_n244), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n227), .A2(new_n230), .B1(new_n241), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G226gat), .ZN(new_n247));
  INV_X1    g046(.A(G233gat), .ZN(new_n248));
  OAI22_X1  g047(.A1(new_n246), .A2(KEYINPUT29), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT72), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n227), .A2(new_n230), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n245), .A2(new_n241), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n247), .A2(new_n248), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT72), .B1(new_n249), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n211), .B1(new_n251), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n249), .A2(new_n256), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n259), .A2(new_n211), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G8gat), .B(G36gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(G64gat), .B(G92gat), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n263), .B(new_n264), .Z(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n258), .A2(new_n261), .A3(KEYINPUT30), .A4(new_n265), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n258), .A2(new_n265), .A3(new_n261), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT73), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT30), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n270), .B1(new_n269), .B2(new_n271), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n267), .B(new_n268), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT39), .ZN(new_n276));
  XNOR2_X1  g075(.A(G127gat), .B(G134gat), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n277), .B(KEYINPUT68), .Z(new_n278));
  XNOR2_X1  g077(.A(G113gat), .B(G120gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT1), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(new_n280), .B2(new_n279), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n277), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n286));
  INV_X1    g085(.A(new_n279), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(new_n286), .B2(new_n287), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G148gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(G141gat), .ZN(new_n292));
  INV_X1    g091(.A(G141gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G148gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n292), .A2(new_n294), .B1(new_n295), .B2(KEYINPUT2), .ZN(new_n296));
  NAND2_X1  g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT74), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n295), .A2(G155gat), .A3(G162gat), .ZN(new_n299));
  INV_X1    g098(.A(G155gat), .ZN(new_n300));
  INV_X1    g099(.A(G162gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n298), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n296), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n297), .B1(new_n302), .B2(KEYINPUT2), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n292), .A2(KEYINPUT75), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n292), .A2(KEYINPUT75), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(new_n294), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n304), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n290), .B(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n276), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n283), .A2(new_n289), .A3(new_n309), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(KEYINPUT4), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n309), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT3), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n309), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n290), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n313), .A2(KEYINPUT4), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n315), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n312), .B1(new_n323), .B2(new_n311), .ZN(new_n324));
  XOR2_X1   g123(.A(G1gat), .B(G29gat), .Z(new_n325));
  XNOR2_X1  g124(.A(G57gat), .B(G85gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n322), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n314), .B1(new_n331), .B2(new_n320), .ZN(new_n332));
  INV_X1    g131(.A(new_n311), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n276), .A3(new_n333), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n324), .A2(KEYINPUT40), .A3(new_n330), .A4(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(new_n335), .B(KEYINPUT81), .Z(new_n336));
  AND3_X1   g135(.A1(new_n324), .A2(new_n330), .A3(new_n334), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n337), .A2(KEYINPUT40), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n332), .A2(new_n333), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n341), .B1(new_n310), .B2(new_n311), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n323), .A2(new_n311), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n345), .A2(KEYINPUT78), .A3(new_n341), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n347), .B1(new_n339), .B2(new_n340), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n344), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n338), .B1(new_n329), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n275), .A2(new_n336), .A3(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(G78gat), .B(G106gat), .Z(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT79), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(G22gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n318), .B1(new_n211), .B2(KEYINPUT29), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n316), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT29), .B1(new_n309), .B2(new_n318), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT80), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n211), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n358), .A2(KEYINPUT80), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(G228gat), .A3(G233gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(G228gat), .A2(G233gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n211), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n357), .B(new_n364), .C1(new_n365), .C2(new_n358), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT31), .B(G50gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n363), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n368), .B1(new_n363), .B2(new_n366), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n355), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n363), .A2(new_n366), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n367), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(new_n354), .A3(new_n369), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT6), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT78), .B1(new_n345), .B2(new_n341), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n339), .A2(new_n347), .A3(new_n340), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n343), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n378), .B1(new_n381), .B2(new_n330), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n344), .B(new_n330), .C1(new_n346), .C2(new_n348), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT82), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n349), .A2(KEYINPUT6), .A3(new_n329), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n349), .A2(new_n329), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT82), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n378), .A4(new_n383), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n385), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT72), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n259), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n392), .A2(new_n365), .A3(new_n250), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT83), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n259), .A2(new_n211), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n393), .A2(KEYINPUT83), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT37), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n266), .A2(KEYINPUT37), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT38), .B1(new_n267), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n262), .A2(KEYINPUT37), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n266), .B1(new_n262), .B2(KEYINPUT37), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT38), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n401), .A2(new_n404), .A3(new_n269), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n351), .B(new_n377), .C1(new_n390), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n267), .A2(new_n268), .ZN(new_n407));
  INV_X1    g206(.A(new_n274), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n407), .B1(new_n408), .B2(new_n272), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n386), .B1(new_n382), .B2(new_n384), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n283), .A2(new_n289), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n254), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G227gat), .A2(G233gat), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n246), .A2(new_n290), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n413), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n417), .A2(KEYINPUT32), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n413), .A2(new_n416), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n414), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT34), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT34), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n419), .A2(new_n422), .A3(new_n414), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT33), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  XOR2_X1   g225(.A(G15gat), .B(G43gat), .Z(new_n427));
  XNOR2_X1  g226(.A(G71gat), .B(G99gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n427), .B(new_n428), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n429), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n432), .A2(new_n421), .A3(new_n423), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n418), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n431), .A2(new_n418), .A3(new_n433), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(KEYINPUT36), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT36), .ZN(new_n438));
  INV_X1    g237(.A(new_n436), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n438), .B1(new_n439), .B2(new_n434), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n411), .A2(new_n376), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n406), .A2(new_n441), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n439), .A2(new_n376), .A3(new_n434), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(new_n409), .A3(new_n410), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT35), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT35), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n390), .A2(new_n446), .A3(new_n409), .A4(new_n443), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n450));
  NOR4_X1   g249(.A1(KEYINPUT86), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT86), .ZN(new_n452));
  NOR2_X1   g251(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n453));
  INV_X1    g252(.A(G36gat), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n450), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(G43gat), .B(G50gat), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n457), .A2(KEYINPUT15), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n457), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n456), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT14), .ZN(new_n461));
  INV_X1    g260(.A(G29gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n462), .A3(new_n454), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n450), .ZN(new_n464));
  NAND2_X1  g263(.A1(G29gat), .A2(G36gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(G50gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(G43gat), .ZN(new_n468));
  INV_X1    g267(.A(G43gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(G50gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n470), .A3(KEYINPUT15), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT85), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n463), .A2(new_n450), .B1(G29gat), .B2(G36gat), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT85), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n474), .A2(new_n475), .A3(new_n471), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n460), .B(KEYINPUT17), .C1(new_n473), .C2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G15gat), .B(G22gat), .ZN(new_n478));
  INV_X1    g277(.A(G1gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT16), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n478), .A2(G1gat), .ZN(new_n482));
  OAI21_X1  g281(.A(G8gat), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n478), .A2(new_n480), .ZN(new_n484));
  INV_X1    g283(.A(G8gat), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n484), .B(new_n485), .C1(G1gat), .C2(new_n478), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n475), .B1(new_n474), .B2(new_n471), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n466), .A2(KEYINPUT85), .A3(new_n472), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n471), .A2(new_n465), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n457), .A2(KEYINPUT15), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n488), .A2(new_n489), .B1(new_n492), .B2(new_n456), .ZN(new_n493));
  XOR2_X1   g292(.A(KEYINPUT87), .B(KEYINPUT17), .Z(new_n494));
  OAI211_X1 g293(.A(new_n477), .B(new_n487), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(G229gat), .A2(G233gat), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n460), .B1(new_n473), .B2(new_n476), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n483), .A2(new_n486), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n495), .A2(KEYINPUT18), .A3(new_n496), .A4(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(new_n496), .B(KEYINPUT13), .Z(new_n501));
  INV_X1    g300(.A(new_n499), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n497), .A2(new_n498), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G113gat), .B(G141gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT84), .B(G197gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT11), .B(G169gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT12), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n495), .A2(new_n496), .A3(new_n499), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT18), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(KEYINPUT89), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n514), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT89), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n512), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n513), .A2(KEYINPUT88), .A3(new_n514), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT88), .B1(new_n513), .B2(new_n514), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n520), .A2(new_n521), .A3(new_n505), .ZN(new_n522));
  INV_X1    g321(.A(new_n511), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n449), .A2(KEYINPUT90), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT90), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n406), .A2(new_n441), .B1(new_n445), .B2(new_n447), .ZN(new_n527));
  INV_X1    g326(.A(new_n524), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G230gat), .A2(G233gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(G85gat), .A2(G92gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NOR2_X1   g331(.A1(G85gat), .A2(G92gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(G99gat), .A2(G106gat), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n533), .B1(KEYINPUT8), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G99gat), .B(G106gat), .Z(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n537), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n539), .A2(new_n532), .A3(new_n535), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G71gat), .A2(G78gat), .ZN(new_n543));
  OR2_X1    g342(.A1(G71gat), .A2(G78gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT9), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G57gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT92), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(G57gat), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n550), .A3(G64gat), .ZN(new_n551));
  INV_X1    g350(.A(G64gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(G57gat), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n551), .A2(KEYINPUT93), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT93), .B1(new_n551), .B2(new_n553), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n546), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT94), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(KEYINPUT94), .B(new_n546), .C1(new_n554), .C2(new_n555), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n544), .A2(new_n543), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT91), .ZN(new_n562));
  XNOR2_X1  g361(.A(G57gat), .B(G64gat), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n561), .B(new_n562), .C1(new_n545), .C2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n547), .A2(G64gat), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n545), .B1(new_n553), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n544), .A2(new_n543), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT91), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n542), .B1(new_n560), .B2(new_n570), .ZN(new_n571));
  AOI211_X1 g370(.A(new_n569), .B(new_n541), .C1(new_n558), .C2(new_n559), .ZN(new_n572));
  NOR3_X1   g371(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT10), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n569), .B1(new_n558), .B2(new_n559), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(KEYINPUT10), .A3(new_n542), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n530), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n551), .A2(new_n553), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT93), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n551), .A2(KEYINPUT93), .A3(new_n553), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT94), .B1(new_n582), .B2(new_n546), .ZN(new_n583));
  INV_X1    g382(.A(new_n559), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n570), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(new_n541), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n574), .A2(new_n542), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n530), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G120gat), .B(G148gat), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT98), .ZN(new_n591));
  XNOR2_X1  g390(.A(G176gat), .B(G204gat), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n591), .B(new_n592), .Z(new_n593));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  INV_X1    g394(.A(new_n530), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT10), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n586), .A2(new_n597), .A3(new_n587), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n596), .B1(new_n598), .B2(new_n575), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n595), .B1(new_n599), .B2(new_n588), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n525), .A2(new_n529), .A3(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G183gat), .B(G211gat), .Z(new_n604));
  OAI211_X1 g403(.A(G231gat), .B(G233gat), .C1(new_n574), .C2(KEYINPUT21), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n585), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT20), .Z(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n609), .A2(new_n611), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n604), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n614), .ZN(new_n616));
  INV_X1    g415(.A(new_n604), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n617), .A3(new_n612), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n487), .B1(new_n585), .B2(new_n606), .ZN(new_n620));
  XOR2_X1   g419(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n615), .A2(new_n618), .A3(new_n622), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n542), .A2(new_n497), .ZN(new_n628));
  NAND2_X1  g427(.A1(G232gat), .A2(G233gat), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT41), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n628), .A2(KEYINPUT96), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT96), .B1(new_n628), .B2(new_n632), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n477), .B(new_n541), .C1(new_n493), .C2(new_n494), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(new_n630), .A3(new_n629), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n629), .A2(new_n630), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n636), .A2(new_n640), .A3(new_n637), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G190gat), .B(G218gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT97), .ZN(new_n644));
  XOR2_X1   g443(.A(G134gat), .B(G162gat), .Z(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n639), .A2(new_n641), .A3(new_n646), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n627), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n603), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(new_n410), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(new_n479), .ZN(G1324gat));
  AND2_X1   g453(.A1(new_n603), .A2(new_n651), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n485), .B1(new_n655), .B2(new_n275), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT16), .B(G8gat), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n652), .A2(new_n409), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT42), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n658), .A2(KEYINPUT42), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(G1325gat));
  NAND2_X1  g460(.A1(new_n440), .A2(new_n437), .ZN(new_n662));
  OAI21_X1  g461(.A(G15gat), .B1(new_n652), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n439), .A2(new_n434), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n665), .A2(G15gat), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n663), .B1(new_n652), .B2(new_n666), .ZN(G1326gat));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n377), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT43), .B(G22gat), .Z(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1327gat));
  XOR2_X1   g469(.A(new_n601), .B(KEYINPUT100), .Z(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(new_n528), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n648), .A2(new_n649), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n674), .B1(new_n442), .B2(new_n448), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n673), .B1(new_n675), .B2(KEYINPUT101), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n677));
  NOR4_X1   g476(.A1(new_n527), .A2(new_n677), .A3(KEYINPUT44), .A4(new_n674), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n627), .B(new_n672), .C1(new_n676), .C2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(G29gat), .B1(new_n679), .B2(new_n410), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n626), .A2(new_n674), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n525), .A2(new_n529), .A3(new_n602), .A4(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n410), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n462), .ZN(new_n684));
  OR3_X1    g483(.A1(new_n682), .A2(KEYINPUT99), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT45), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT99), .B1(new_n682), .B2(new_n684), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n686), .B1(new_n685), .B2(new_n687), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n680), .B1(new_n688), .B2(new_n689), .ZN(G1328gat));
  NOR3_X1   g489(.A1(new_n682), .A2(G36gat), .A3(new_n409), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT46), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(G36gat), .B1(new_n679), .B2(new_n409), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n692), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(G1329gat));
  OAI21_X1  g495(.A(new_n469), .B1(new_n682), .B2(new_n665), .ZN(new_n697));
  INV_X1    g496(.A(new_n662), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(G43gat), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n697), .B1(new_n679), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g500(.A(G50gat), .B1(new_n679), .B2(new_n377), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n603), .A2(new_n467), .A3(new_n376), .A4(new_n681), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT48), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n704), .B1(new_n702), .B2(new_n703), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(G1331gat));
  INV_X1    g506(.A(new_n671), .ZN(new_n708));
  NOR4_X1   g507(.A1(new_n708), .A2(new_n627), .A3(new_n650), .A4(new_n524), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n449), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n410), .B(KEYINPUT102), .Z(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n548), .A2(new_n550), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n712), .B(new_n713), .Z(G1332gat));
  INV_X1    g513(.A(new_n710), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n409), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT103), .ZN(new_n718));
  NOR2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1333gat));
  NOR3_X1   g519(.A1(new_n710), .A2(G71gat), .A3(new_n665), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n715), .A2(new_n698), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(G71gat), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT104), .B(KEYINPUT50), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1334gat));
  NAND2_X1  g524(.A1(new_n715), .A2(new_n376), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g526(.A1(new_n602), .A2(new_n524), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n627), .B(new_n728), .C1(new_n676), .C2(new_n678), .ZN(new_n729));
  OAI21_X1  g528(.A(G85gat), .B1(new_n729), .B2(new_n410), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n626), .A2(new_n524), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n732), .B1(new_n675), .B2(KEYINPUT105), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n527), .B2(new_n674), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n733), .A2(KEYINPUT51), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT51), .B1(new_n733), .B2(new_n735), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n601), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n410), .A2(G85gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n730), .B1(new_n738), .B2(new_n739), .ZN(G1336gat));
  NOR2_X1   g539(.A1(new_n409), .A2(G92gat), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n671), .B(new_n741), .C1(new_n736), .C2(new_n737), .ZN(new_n742));
  OAI21_X1  g541(.A(G92gat), .B1(new_n729), .B2(new_n409), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT52), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n742), .A2(new_n743), .A3(new_n744), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(G1337gat));
  OAI21_X1  g548(.A(G99gat), .B1(new_n729), .B2(new_n662), .ZN(new_n750));
  OR2_X1    g549(.A1(new_n665), .A2(G99gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n738), .B2(new_n751), .ZN(G1338gat));
  OAI21_X1  g551(.A(KEYINPUT107), .B1(new_n729), .B2(new_n377), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n449), .A2(KEYINPUT101), .A3(new_n650), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT44), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n675), .A2(KEYINPUT101), .A3(new_n673), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n626), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n757), .A2(new_n758), .A3(new_n376), .A4(new_n728), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n753), .A2(new_n759), .A3(G106gat), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n449), .A2(KEYINPUT105), .A3(new_n650), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n761), .A2(new_n735), .A3(new_n731), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n733), .A2(KEYINPUT51), .A3(new_n735), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n708), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n377), .A2(G106gat), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT53), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n760), .A2(new_n768), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n671), .B(new_n767), .C1(new_n736), .C2(new_n737), .ZN(new_n770));
  OAI21_X1  g569(.A(G106gat), .B1(new_n729), .B2(new_n377), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT53), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n769), .A2(new_n773), .ZN(G1339gat));
  NAND2_X1  g573(.A1(new_n575), .A2(new_n596), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT54), .B1(new_n573), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT55), .B1(new_n776), .B2(new_n599), .ZN(new_n777));
  XOR2_X1   g576(.A(KEYINPUT108), .B(KEYINPUT54), .Z(new_n778));
  OAI211_X1 g577(.A(new_n530), .B(new_n778), .C1(new_n573), .C2(new_n576), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n595), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n594), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT109), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n593), .B1(new_n599), .B2(new_n778), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n530), .B1(new_n572), .B2(KEYINPUT10), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n784), .B1(new_n598), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n577), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n783), .A2(new_n787), .A3(KEYINPUT55), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n789), .A3(new_n594), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT55), .B1(new_n783), .B2(new_n787), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n782), .A2(new_n524), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n495), .A2(new_n499), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(G229gat), .A3(G233gat), .ZN(new_n795));
  OR3_X1    g594(.A1(new_n502), .A2(new_n503), .A3(new_n501), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n510), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n518), .A2(new_n515), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n797), .B1(new_n798), .B2(new_n512), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n601), .A2(new_n799), .A3(KEYINPUT110), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT110), .B1(new_n601), .B2(new_n799), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n650), .B1(new_n793), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n791), .B1(new_n781), .B2(KEYINPUT109), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n804), .A2(new_n650), .A3(new_n799), .A4(new_n790), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n627), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  AND4_X1   g606(.A1(new_n626), .A2(new_n674), .A3(new_n528), .A4(new_n602), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n711), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n810), .A2(new_n409), .A3(new_n443), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT111), .Z(new_n812));
  NOR2_X1   g611(.A1(new_n528), .A2(G113gat), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(KEYINPUT112), .Z(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n376), .B1(new_n807), .B2(new_n809), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n816), .A2(new_n683), .A3(new_n409), .A4(new_n664), .ZN(new_n817));
  OAI21_X1  g616(.A(G113gat), .B1(new_n817), .B2(new_n528), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n818), .ZN(G1340gat));
  INV_X1    g618(.A(G120gat), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n812), .A2(new_n820), .A3(new_n601), .ZN(new_n821));
  OAI21_X1  g620(.A(G120gat), .B1(new_n817), .B2(new_n708), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1341gat));
  OAI21_X1  g622(.A(G127gat), .B1(new_n817), .B2(new_n627), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n627), .A2(G127gat), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n811), .B2(new_n825), .ZN(G1342gat));
  OR3_X1    g625(.A1(new_n811), .A2(G134gat), .A3(new_n674), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n827), .A2(KEYINPUT56), .ZN(new_n828));
  OAI21_X1  g627(.A(G134gat), .B1(new_n817), .B2(new_n674), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(KEYINPUT56), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(G1343gat));
  NOR3_X1   g630(.A1(new_n698), .A2(new_n410), .A3(new_n275), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n528), .A2(new_n293), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n601), .A2(new_n799), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n788), .A2(new_n524), .A3(new_n594), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n779), .B(new_n595), .C1(new_n776), .C2(new_n599), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT113), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT113), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n783), .A2(new_n787), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n835), .B1(new_n836), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n805), .B1(new_n843), .B2(new_n650), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n808), .B1(new_n844), .B2(new_n627), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n376), .A2(KEYINPUT57), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n834), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n846), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n788), .A2(new_n524), .A3(new_n594), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT55), .B1(new_n837), .B2(KEYINPUT113), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n841), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n674), .B1(new_n851), .B2(new_n835), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n626), .B1(new_n852), .B2(new_n805), .ZN(new_n853));
  OAI211_X1 g652(.A(KEYINPUT114), .B(new_n848), .C1(new_n853), .C2(new_n808), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n807), .A2(new_n809), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT57), .B1(new_n856), .B2(new_n376), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n832), .B(new_n833), .C1(new_n855), .C2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n377), .B1(new_n440), .B2(new_n437), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(new_n409), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n810), .A2(new_n524), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n293), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT116), .B1(new_n858), .B2(new_n862), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n865), .B(KEYINPUT58), .C1(new_n864), .C2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n863), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT58), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(KEYINPUT115), .A3(new_n871), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n867), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n868), .B1(new_n867), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(G1344gat));
  NAND2_X1  g674(.A1(new_n810), .A2(new_n860), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT59), .B1(new_n876), .B2(new_n602), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n291), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n855), .A2(new_n857), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n832), .A2(new_n601), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(KEYINPUT59), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n804), .A2(new_n650), .A3(new_n790), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n799), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n626), .B1(new_n887), .B2(new_n852), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n376), .B1(new_n888), .B2(new_n808), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n890));
  AOI22_X1  g689(.A1(new_n889), .A2(new_n890), .B1(new_n856), .B2(new_n848), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n880), .ZN(new_n892));
  NAND2_X1  g691(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n878), .B(new_n882), .C1(new_n892), .C2(new_n893), .ZN(G1345gat));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n832), .ZN(new_n895));
  OAI21_X1  g694(.A(G155gat), .B1(new_n895), .B2(new_n627), .ZN(new_n896));
  INV_X1    g695(.A(new_n876), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(new_n300), .A3(new_n626), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(G1346gat));
  NAND3_X1  g698(.A1(new_n897), .A2(new_n301), .A3(new_n650), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT119), .ZN(new_n901));
  OAI21_X1  g700(.A(G162gat), .B1(new_n895), .B2(new_n674), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1347gat));
  INV_X1    g702(.A(new_n711), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(new_n409), .A3(new_n665), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n816), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n906), .A2(new_n212), .A3(new_n528), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n443), .A2(new_n275), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n908), .B(KEYINPUT120), .Z(new_n909));
  AOI21_X1  g708(.A(new_n683), .B1(new_n807), .B2(new_n809), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(G169gat), .B1(new_n912), .B2(new_n524), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n907), .A2(new_n913), .ZN(G1348gat));
  NAND4_X1  g713(.A1(new_n905), .A2(new_n234), .A3(new_n671), .A4(new_n816), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n915), .A2(KEYINPUT121), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(KEYINPUT121), .ZN(new_n917));
  AOI21_X1  g716(.A(G176gat), .B1(new_n912), .B2(new_n601), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(G1349gat));
  OAI21_X1  g718(.A(G183gat), .B1(new_n906), .B2(new_n627), .ZN(new_n920));
  NAND2_X1  g719(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n626), .A2(new_n221), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n920), .B(new_n921), .C1(new_n911), .C2(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n924));
  XOR2_X1   g723(.A(new_n923), .B(new_n924), .Z(G1350gat));
  OAI21_X1  g724(.A(G190gat), .B1(new_n906), .B2(new_n674), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT61), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n912), .A2(new_n216), .A3(new_n650), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1351gat));
  NAND2_X1  g728(.A1(new_n859), .A2(new_n275), .ZN(new_n930));
  XOR2_X1   g729(.A(new_n930), .B(KEYINPUT123), .Z(new_n931));
  AND2_X1   g730(.A1(new_n931), .A2(new_n910), .ZN(new_n932));
  AOI21_X1  g731(.A(G197gat), .B1(new_n932), .B2(new_n524), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n711), .A2(new_n275), .A3(new_n662), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n891), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n524), .A2(G197gat), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(G1352gat));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n938));
  AOI21_X1  g737(.A(G204gat), .B1(new_n938), .B2(KEYINPUT62), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n932), .A2(new_n601), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n938), .A2(KEYINPUT62), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n940), .B(new_n941), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n891), .A2(new_n708), .A3(new_n934), .ZN(new_n943));
  INV_X1    g742(.A(G204gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(G1353gat));
  NAND2_X1  g744(.A1(new_n935), .A2(new_n626), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G211gat), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n947), .A2(KEYINPUT63), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(KEYINPUT63), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n932), .A2(new_n203), .A3(new_n626), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT125), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(G1354gat));
  NAND3_X1  g751(.A1(new_n931), .A2(new_n650), .A3(new_n910), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n204), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT126), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n935), .A2(G218gat), .A3(new_n650), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n955), .A2(KEYINPUT127), .A3(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1355gat));
endmodule


