//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n188), .A2(KEYINPUT64), .A3(G143), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n192), .A2(new_n193), .A3(G128), .A4(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  OAI21_X1  g011(.A(G128), .B1(new_n197), .B2(new_n193), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n198), .B1(new_n197), .B2(new_n190), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT11), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT65), .A2(G134), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT65), .A2(G134), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G131), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n201), .A2(KEYINPUT11), .A3(G134), .ZN(new_n211));
  OR2_X1    g025(.A1(new_n201), .A2(KEYINPUT11), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n205), .A2(new_n210), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n201), .B1(new_n203), .B2(new_n204), .ZN(new_n214));
  NAND2_X1  g028(.A1(G134), .A2(G137), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(G131), .A3(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n200), .A2(new_n213), .A3(new_n216), .ZN(new_n217));
  OR2_X1    g031(.A1(KEYINPUT65), .A2(G134), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT65), .A2(G134), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n218), .A2(new_n219), .B1(KEYINPUT11), .B2(new_n201), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n211), .B1(KEYINPUT11), .B2(new_n201), .ZN(new_n221));
  OAI21_X1  g035(.A(G131), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n213), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n191), .B1(new_n196), .B2(G146), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n194), .B(new_n225), .C1(new_n226), .C2(new_n197), .ZN(new_n227));
  OR2_X1    g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n224), .B(new_n228), .C1(new_n197), .C2(new_n190), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n223), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n217), .A2(new_n231), .A3(KEYINPUT30), .ZN(new_n232));
  NAND3_X1  g046(.A1(KEYINPUT69), .A2(KEYINPUT2), .A3(G113), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(KEYINPUT69), .B1(KEYINPUT2), .B2(G113), .ZN(new_n235));
  OAI22_X1  g049(.A1(new_n234), .A2(new_n235), .B1(KEYINPUT2), .B2(G113), .ZN(new_n236));
  INV_X1    g050(.A(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G116), .ZN(new_n238));
  INV_X1    g052(.A(G116), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G119), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT70), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(KEYINPUT2), .A2(G113), .ZN(new_n243));
  NAND2_X1  g057(.A1(KEYINPUT2), .A2(G113), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n243), .B1(new_n246), .B2(new_n233), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n248));
  XNOR2_X1  g062(.A(G116), .B(G119), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n242), .A2(new_n250), .B1(new_n236), .B2(new_n241), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n231), .A2(KEYINPUT67), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n223), .A2(new_n254), .A3(new_n230), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n213), .A2(KEYINPUT68), .A3(new_n216), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT68), .B1(new_n213), .B2(new_n216), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n253), .A2(new_n255), .B1(new_n258), .B2(new_n200), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n232), .B(new_n252), .C1(new_n259), .C2(KEYINPUT30), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n217), .A2(new_n231), .A3(new_n251), .ZN(new_n261));
  INV_X1    g075(.A(G237), .ZN(new_n262));
  INV_X1    g076(.A(G953), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n263), .A3(G210), .ZN(new_n264));
  XOR2_X1   g078(.A(new_n264), .B(KEYINPUT27), .Z(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(KEYINPUT26), .ZN(new_n266));
  INV_X1    g080(.A(G101), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n260), .A2(new_n261), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT31), .ZN(new_n270));
  INV_X1    g084(.A(new_n257), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n213), .A2(KEYINPUT68), .A3(new_n216), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n200), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n255), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n254), .B1(new_n223), .B2(new_n230), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n261), .A2(KEYINPUT28), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n217), .A2(new_n231), .A3(new_n251), .A4(new_n278), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n276), .A2(new_n252), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  OR2_X1    g094(.A1(new_n280), .A2(new_n268), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT31), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n260), .A2(new_n282), .A3(new_n261), .A4(new_n268), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n270), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(G472), .A2(G902), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n284), .A2(KEYINPUT71), .A3(new_n285), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT32), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n284), .A2(KEYINPUT32), .A3(new_n285), .ZN(new_n291));
  INV_X1    g105(.A(new_n268), .ZN(new_n292));
  INV_X1    g106(.A(new_n260), .ZN(new_n293));
  INV_X1    g107(.A(new_n261), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n280), .A2(new_n268), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT72), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n276), .A2(new_n252), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n277), .A2(new_n279), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT72), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n268), .A4(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n295), .A2(new_n297), .A3(new_n298), .A4(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n292), .A2(new_n298), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n251), .B1(new_n217), .B2(new_n231), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n305), .B1(new_n277), .B2(new_n279), .ZN(new_n306));
  AOI21_X1  g120(.A(G902), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G472), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n291), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n187), .B1(new_n290), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT32), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n284), .A2(KEYINPUT71), .A3(new_n285), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT71), .B1(new_n284), .B2(new_n285), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n291), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n309), .B1(new_n303), .B2(new_n307), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n318), .A3(KEYINPUT73), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n311), .A2(new_n319), .ZN(new_n320));
  XOR2_X1   g134(.A(KEYINPUT9), .B(G234), .Z(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(G221), .B1(new_n322), .B2(G902), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G469), .ZN(new_n325));
  INV_X1    g139(.A(G902), .ZN(new_n326));
  INV_X1    g140(.A(G104), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G107), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n327), .A2(G107), .ZN(new_n330));
  OAI21_X1  g144(.A(G101), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT3), .B1(new_n327), .B2(G107), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n333));
  INV_X1    g147(.A(G107), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(G104), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n332), .A2(new_n335), .A3(new_n267), .A4(new_n328), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n200), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n192), .A2(new_n194), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n198), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n337), .B1(new_n341), .B2(new_n195), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n223), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT12), .B1(new_n223), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n343), .B(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n332), .A2(new_n335), .A3(new_n328), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G101), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(KEYINPUT4), .A3(new_n336), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n347), .A2(new_n350), .A3(G101), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n230), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n200), .A2(new_n338), .A3(KEYINPUT10), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n352), .B(new_n353), .C1(new_n342), .C2(KEYINPUT10), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n354), .A2(new_n223), .ZN(new_n355));
  XNOR2_X1  g169(.A(G110), .B(G140), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n263), .A2(G227), .ZN(new_n357));
  XOR2_X1   g171(.A(new_n356), .B(new_n357), .Z(new_n358));
  AND3_X1   g172(.A1(new_n346), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n354), .A2(new_n223), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n358), .B1(new_n355), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n325), .B(new_n326), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n361), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n346), .A2(new_n355), .A3(new_n358), .ZN(new_n366));
  AOI21_X1  g180(.A(G902), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(KEYINPUT81), .A3(new_n325), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n358), .B1(new_n346), .B2(new_n355), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n355), .A2(new_n358), .A3(new_n360), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(G469), .B1(new_n372), .B2(G902), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n324), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(G214), .B1(G237), .B2(G902), .ZN(new_n375));
  XOR2_X1   g189(.A(new_n375), .B(KEYINPUT82), .Z(new_n376));
  OAI21_X1  g190(.A(G113), .B1(new_n238), .B2(KEYINPUT5), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT86), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n380));
  OAI211_X1 g194(.A(KEYINPUT86), .B(G113), .C1(new_n238), .C2(KEYINPUT5), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n236), .A2(KEYINPUT70), .A3(new_n241), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n248), .B1(new_n247), .B2(new_n249), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT87), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n242), .A2(new_n250), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT87), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(new_n382), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(new_n338), .A3(new_n389), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n380), .B(G113), .C1(KEYINPUT5), .C2(new_n238), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(new_n337), .A3(new_n391), .ZN(new_n392));
  XOR2_X1   g206(.A(G110), .B(G122), .Z(new_n393));
  XOR2_X1   g207(.A(KEYINPUT85), .B(KEYINPUT8), .Z(new_n394));
  XNOR2_X1  g208(.A(new_n393), .B(new_n394), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n390), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n387), .A2(new_n338), .A3(new_n391), .ZN(new_n397));
  INV_X1    g211(.A(new_n393), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n349), .A2(new_n351), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n397), .B(new_n398), .C1(new_n399), .C2(new_n251), .ZN(new_n400));
  INV_X1    g214(.A(G125), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n200), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n230), .A2(G125), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n263), .A2(G224), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n404), .B(KEYINPUT83), .Z(new_n405));
  AND4_X1   g219(.A1(KEYINPUT7), .A2(new_n402), .A3(new_n403), .A4(new_n405), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n402), .A2(new_n403), .B1(KEYINPUT7), .B2(new_n405), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n400), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n326), .B1(new_n396), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT88), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n402), .A2(new_n403), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT84), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n411), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n405), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n411), .B(KEYINPUT84), .ZN(new_n415));
  INV_X1    g229(.A(new_n405), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n397), .B1(new_n251), .B2(new_n399), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT6), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n393), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n393), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(KEYINPUT6), .A3(new_n400), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n414), .A2(new_n417), .A3(new_n420), .A4(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT88), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n424), .B(new_n326), .C1(new_n396), .C2(new_n408), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n410), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G210), .B1(G237), .B2(G902), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(KEYINPUT89), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n428), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT89), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n410), .A2(new_n423), .A3(new_n427), .A4(new_n425), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n374), .A2(new_n376), .A3(new_n429), .A4(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G217), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(G234), .B2(new_n326), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT78), .ZN(new_n439));
  INV_X1    g253(.A(G128), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G119), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT23), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n237), .A2(G128), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n440), .A2(KEYINPUT23), .A3(G119), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G110), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT24), .B(G110), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(KEYINPUT74), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n444), .A2(new_n441), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT76), .ZN(new_n452));
  INV_X1    g266(.A(G140), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G125), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n401), .A2(G140), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT75), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n453), .A2(KEYINPUT75), .A3(G125), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n452), .B1(new_n459), .B2(KEYINPUT16), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT16), .ZN(new_n461));
  AOI211_X1 g275(.A(KEYINPUT76), .B(new_n461), .C1(new_n457), .C2(new_n458), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n461), .A2(new_n453), .A3(G125), .ZN(new_n464));
  AOI21_X1  g278(.A(G146), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n453), .A2(KEYINPUT75), .A3(G125), .ZN(new_n466));
  XNOR2_X1  g280(.A(G125), .B(G140), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n466), .B1(new_n467), .B2(new_n456), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT76), .B1(new_n468), .B2(new_n461), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n459), .A2(new_n452), .A3(KEYINPUT16), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n469), .A2(G146), .A3(new_n464), .A4(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n447), .B(new_n451), .C1(new_n465), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n467), .A2(new_n188), .ZN(new_n474));
  OAI22_X1  g288(.A1(new_n449), .A2(new_n450), .B1(G110), .B2(new_n446), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n471), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n263), .A2(G221), .A3(G234), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT22), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(new_n201), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n201), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT77), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT77), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n480), .A2(new_n201), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n485), .B1(new_n486), .B2(new_n481), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n439), .B1(new_n478), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n488), .ZN(new_n490));
  AOI211_X1 g304(.A(KEYINPUT78), .B(new_n490), .C1(new_n473), .C2(new_n477), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n473), .A2(new_n477), .A3(new_n482), .A4(new_n483), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n492), .A2(KEYINPUT25), .A3(new_n326), .A4(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n451), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n469), .A2(new_n464), .A3(new_n470), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n188), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n495), .B1(new_n497), .B2(new_n471), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n476), .B1(new_n498), .B2(new_n447), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT78), .B1(new_n499), .B2(new_n490), .ZN(new_n500));
  INV_X1    g314(.A(new_n447), .ZN(new_n501));
  AOI211_X1 g315(.A(new_n501), .B(new_n495), .C1(new_n497), .C2(new_n471), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n439), .B(new_n488), .C1(new_n502), .C2(new_n476), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n500), .A2(new_n326), .A3(new_n493), .A4(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT25), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n438), .B1(new_n494), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n437), .A2(G902), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT79), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n492), .A2(new_n509), .A3(new_n493), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G475), .ZN(new_n512));
  XOR2_X1   g326(.A(G113), .B(G122), .Z(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT92), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(new_n327), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT90), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n454), .A2(new_n455), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n517), .B1(new_n518), .B2(KEYINPUT19), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT19), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n519), .B1(new_n459), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n468), .A2(new_n517), .A3(KEYINPUT19), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n522), .A3(new_n188), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n471), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n262), .A2(new_n263), .A3(G214), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(G143), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n210), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n210), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n471), .A2(KEYINPUT91), .A3(new_n523), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n526), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(KEYINPUT18), .A2(G131), .ZN(new_n536));
  XOR2_X1   g350(.A(new_n528), .B(new_n536), .Z(new_n537));
  OAI21_X1  g351(.A(new_n474), .B1(new_n459), .B2(new_n188), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n516), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n531), .A2(new_n532), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n529), .A2(KEYINPUT17), .A3(new_n530), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n497), .A2(new_n471), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n516), .A3(new_n539), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n512), .B(new_n326), .C1(new_n540), .C2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT20), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n534), .A2(new_n533), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT91), .B1(new_n471), .B2(new_n523), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n539), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n515), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n545), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n554), .A2(KEYINPUT20), .A3(new_n512), .A4(new_n326), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n196), .A2(G128), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n440), .A2(G143), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT93), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT93), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n559), .A2(new_n560), .B1(new_n218), .B2(new_n219), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT13), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n557), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n556), .A2(new_n563), .ZN(new_n566));
  OAI21_X1  g380(.A(G134), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G122), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G116), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n239), .A2(G122), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(new_n334), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n562), .A2(new_n567), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(KEYINPUT14), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n569), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n570), .A2(KEYINPUT14), .ZN(new_n576));
  OAI21_X1  g390(.A(G107), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT94), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n571), .A2(new_n334), .ZN(new_n579));
  INV_X1    g393(.A(new_n560), .ZN(new_n580));
  NOR4_X1   g394(.A1(new_n580), .A2(new_n558), .A3(new_n204), .A4(new_n203), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n579), .B1(new_n581), .B2(new_n561), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n573), .B1(new_n578), .B2(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n322), .A2(new_n436), .A3(G953), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n573), .B(new_n584), .C1(new_n578), .C2(new_n582), .ZN(new_n587));
  AOI21_X1  g401(.A(G902), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(G478), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(KEYINPUT15), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n588), .B(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n516), .B1(new_n544), .B2(new_n539), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n326), .B1(new_n546), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G475), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n549), .A2(new_n555), .A3(new_n591), .A4(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(G952), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(G953), .ZN(new_n597));
  NAND2_X1  g411(.A1(G234), .A2(G237), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT21), .B(G898), .Z(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n598), .A2(G902), .A3(G953), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n600), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n595), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n320), .A2(new_n435), .A3(new_n511), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  AOI21_X1  g422(.A(new_n309), .B1(new_n284), .B2(new_n326), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n288), .B2(new_n289), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(new_n374), .A3(new_n511), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT95), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT95), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n610), .A2(new_n374), .A3(new_n511), .A4(new_n613), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n430), .A2(new_n432), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n615), .A2(new_n375), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n586), .A2(new_n587), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n586), .A2(KEYINPUT33), .A3(new_n587), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n620), .A2(new_n621), .A3(G478), .A4(new_n326), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n588), .A2(G478), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n622), .B1(KEYINPUT96), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n624), .B1(KEYINPUT96), .B2(new_n622), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n549), .A2(new_n594), .A3(new_n555), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(new_n605), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n617), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  OR2_X1    g445(.A1(new_n626), .A2(new_n591), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n605), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT97), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n617), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G107), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  INV_X1    g452(.A(KEYINPUT98), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n488), .A2(KEYINPUT36), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n478), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n509), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n639), .B1(new_n507), .B2(new_n643), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n504), .A2(new_n505), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n504), .A2(new_n505), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n437), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(KEYINPUT98), .A3(new_n642), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n606), .ZN(new_n650));
  INV_X1    g464(.A(new_n609), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n651), .B1(new_n313), .B2(new_n314), .ZN(new_n652));
  NOR4_X1   g466(.A1(new_n434), .A2(new_n649), .A3(new_n650), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT37), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G110), .ZN(G12));
  INV_X1    g469(.A(new_n649), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT99), .B(G900), .Z(new_n657));
  AOI21_X1  g471(.A(new_n600), .B1(new_n604), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n632), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n374), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n616), .A2(new_n375), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n320), .A2(new_n656), .A3(new_n659), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  NAND2_X1  g478(.A1(new_n433), .A2(new_n429), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT38), .ZN(new_n666));
  INV_X1    g480(.A(new_n591), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n626), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n649), .A2(new_n375), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT100), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n292), .B1(new_n305), .B2(new_n294), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n269), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(G472), .B1(new_n674), .B2(G902), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n315), .A2(new_n291), .A3(new_n675), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n672), .B(new_n676), .C1(new_n671), .C2(new_n670), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n658), .B(KEYINPUT39), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n660), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT40), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n679), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G143), .ZN(G45));
  INV_X1    g499(.A(new_n658), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n625), .A2(new_n626), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT102), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n320), .A2(new_n656), .A3(new_n662), .A4(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT103), .B(G146), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G48));
  INV_X1    g505(.A(new_n511), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n311), .B2(new_n319), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n359), .A2(new_n361), .ZN(new_n694));
  OAI211_X1 g508(.A(KEYINPUT104), .B(G469), .C1(new_n694), .C2(G902), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n696), .B1(new_n367), .B2(new_n325), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n323), .A3(new_n369), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n661), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n693), .A2(new_n628), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT41), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G113), .ZN(G15));
  NAND3_X1  g517(.A1(new_n635), .A2(new_n693), .A3(new_n700), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  AND3_X1   g519(.A1(new_n644), .A2(new_n648), .A3(new_n606), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n315), .A2(new_n318), .A3(KEYINPUT73), .ZN(new_n707));
  AOI21_X1  g521(.A(KEYINPUT73), .B1(new_n315), .B2(new_n318), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n706), .B(new_n700), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT105), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n320), .A2(new_n711), .A3(new_n706), .A4(new_n700), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G119), .ZN(G21));
  NOR2_X1   g528(.A1(new_n306), .A2(new_n268), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n269), .B2(KEYINPUT31), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n716), .A2(KEYINPUT106), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n283), .B1(new_n716), .B2(KEYINPUT106), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n285), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n719), .A2(new_n651), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n720), .A2(new_n511), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n668), .A2(new_n605), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n700), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G122), .ZN(G24));
  NAND4_X1  g538(.A1(new_n688), .A2(new_n656), .A3(new_n700), .A4(new_n720), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G125), .ZN(G27));
  INV_X1    g540(.A(KEYINPUT42), .ZN(new_n727));
  INV_X1    g541(.A(new_n375), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n433), .B2(new_n429), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n729), .A2(KEYINPUT107), .A3(new_n374), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT107), .B1(new_n729), .B2(new_n374), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n688), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n511), .B1(new_n707), .B2(new_n708), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n727), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT32), .B1(new_n284), .B2(new_n285), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n511), .B1(new_n310), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n727), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n737), .B(new_n688), .C1(new_n731), .C2(new_n730), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G131), .ZN(G33));
  OR2_X1    g554(.A1(new_n730), .A2(new_n731), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n693), .A3(new_n659), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  OAI21_X1  g557(.A(G469), .B1(new_n372), .B2(KEYINPUT45), .ZN(new_n744));
  XOR2_X1   g558(.A(new_n744), .B(KEYINPUT108), .Z(new_n745));
  NAND2_X1  g559(.A1(new_n372), .A2(KEYINPUT45), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(G469), .A2(G902), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT46), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n749), .A2(KEYINPUT109), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n747), .A2(KEYINPUT46), .A3(new_n748), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(KEYINPUT109), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n750), .A2(new_n369), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n323), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n681), .ZN(new_n755));
  INV_X1    g569(.A(new_n729), .ZN(new_n756));
  INV_X1    g570(.A(new_n625), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(new_n626), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT43), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n759), .A2(new_n652), .A3(new_n656), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n756), .B1(new_n760), .B2(KEYINPUT44), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n755), .B(new_n761), .C1(KEYINPUT44), .C2(new_n760), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  NAND2_X1  g577(.A1(new_n754), .A2(KEYINPUT47), .ZN(new_n764));
  INV_X1    g578(.A(new_n688), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n765), .A2(new_n320), .A3(new_n511), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT47), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n753), .A2(new_n767), .A3(new_n323), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n764), .A2(new_n729), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  AND2_X1   g584(.A1(new_n759), .A2(new_n600), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n771), .A2(new_n721), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n764), .A2(new_n768), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n698), .A2(new_n369), .ZN(new_n774));
  XOR2_X1   g588(.A(new_n774), .B(KEYINPUT110), .Z(new_n775));
  AND2_X1   g589(.A1(new_n775), .A2(new_n324), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n729), .B(new_n772), .C1(new_n773), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n676), .A2(new_n692), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n756), .A2(new_n699), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n779), .A3(new_n600), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n780), .A2(new_n626), .A3(new_n625), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n774), .A2(new_n323), .A3(new_n728), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n782), .A2(KEYINPUT117), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(KEYINPUT117), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n772), .A2(new_n666), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n781), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n771), .A2(new_n656), .A3(new_n720), .A4(new_n779), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n777), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n771), .A2(new_n779), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT118), .B1(new_n794), .B2(new_n736), .ZN(new_n795));
  OAI221_X1 g609(.A(new_n597), .B1(new_n627), .B2(new_n780), .C1(new_n795), .C2(KEYINPUT48), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT48), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n794), .A2(new_n736), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n796), .B1(new_n800), .B2(new_n795), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n777), .A2(new_n789), .A3(KEYINPUT51), .A4(new_n790), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n793), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n435), .A2(new_n706), .A3(new_n610), .ZN(new_n804));
  INV_X1    g618(.A(new_n605), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n632), .A2(new_n627), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n612), .A2(new_n805), .A3(new_n614), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n376), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n665), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n607), .B(new_n804), .C1(new_n807), .C2(new_n810), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n741), .A2(new_n693), .A3(new_n659), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n688), .B(new_n720), .C1(new_n730), .C2(new_n731), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n814), .B1(new_n595), .B2(new_n658), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n374), .A2(new_n665), .A3(new_n375), .A4(new_n815), .ZN(new_n816));
  OR3_X1    g630(.A1(new_n595), .A2(new_n814), .A3(new_n658), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n816), .B(new_n817), .C1(new_n707), .C2(new_n708), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n649), .B1(new_n813), .B2(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n811), .A2(new_n812), .A3(new_n819), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n693), .B(new_n700), .C1(new_n635), .C2(new_n628), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n713), .A2(new_n723), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n820), .A2(new_n822), .A3(new_n823), .A4(new_n739), .ZN(new_n824));
  INV_X1    g638(.A(new_n723), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(new_n710), .B2(new_n712), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n739), .A3(new_n821), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n813), .A2(new_n818), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n656), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n692), .B(new_n650), .C1(new_n311), .C2(new_n319), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n653), .B1(new_n830), .B2(new_n435), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n615), .A2(new_n809), .A3(new_n805), .A4(new_n806), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n829), .A2(new_n831), .A3(new_n832), .A4(new_n742), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT112), .B1(new_n827), .B2(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n507), .A2(new_n643), .A3(new_n658), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT113), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n668), .B1(new_n835), .B2(new_n836), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n662), .A3(new_n676), .A4(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n663), .A2(new_n689), .A3(new_n839), .A4(new_n725), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n824), .A2(new_n834), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n845), .A2(KEYINPUT114), .A3(new_n846), .ZN(new_n847));
  OR3_X1    g661(.A1(new_n843), .A2(KEYINPUT114), .A3(new_n844), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(KEYINPUT54), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n772), .A2(new_n700), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n851), .A2(new_n713), .A3(new_n723), .A4(new_n821), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n851), .B1(new_n826), .B2(new_n821), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n739), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT116), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n833), .A2(new_n844), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n856), .A2(new_n842), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n858), .B(new_n739), .C1(new_n852), .C2(new_n853), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n855), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(new_n846), .A3(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n803), .A2(new_n849), .A3(new_n850), .A4(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(G952), .B2(G953), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n775), .B(KEYINPUT49), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n676), .A2(new_n692), .A3(new_n324), .A4(new_n808), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n865), .A2(new_n666), .A3(new_n758), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n864), .A2(new_n867), .ZN(G75));
  AOI21_X1  g682(.A(new_n326), .B1(new_n860), .B2(new_n846), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT56), .B1(new_n869), .B2(G210), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n414), .A2(new_n417), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n422), .A2(new_n420), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n423), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT55), .Z(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n876), .B1(KEYINPUT119), .B2(new_n877), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n870), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n596), .A2(G953), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n870), .A2(new_n878), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(G51));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n748), .B(KEYINPUT57), .Z(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n860), .A2(new_n846), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(KEYINPUT54), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n885), .B1(new_n887), .B2(new_n862), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n883), .B1(new_n888), .B2(new_n694), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n869), .A2(new_n746), .A3(new_n745), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n860), .A2(new_n846), .A3(new_n861), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n861), .B1(new_n860), .B2(new_n846), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n884), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n694), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(KEYINPUT120), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n889), .A2(new_n890), .A3(new_n895), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n896), .A2(new_n880), .ZN(G54));
  NAND3_X1  g711(.A1(new_n869), .A2(KEYINPUT58), .A3(G475), .ZN(new_n898));
  INV_X1    g712(.A(new_n554), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n900), .A2(new_n880), .A3(new_n901), .ZN(G60));
  AND2_X1   g716(.A1(new_n620), .A2(new_n621), .ZN(new_n903));
  NAND2_X1  g717(.A1(G478), .A2(G902), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT59), .Z(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n903), .B(new_n906), .C1(new_n891), .C2(new_n892), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n905), .B1(new_n849), .B2(new_n862), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n880), .B(new_n907), .C1(new_n908), .C2(new_n903), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(G63));
  XNOR2_X1  g724(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n436), .A2(new_n326), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n860), .B2(new_n846), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n641), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT122), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n492), .A2(new_n493), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n917), .A2(KEYINPUT61), .A3(new_n880), .A4(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n916), .A2(KEYINPUT122), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n915), .B2(new_n641), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n880), .B(new_n919), .C1(new_n921), .C2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n920), .A2(new_n926), .ZN(G66));
  INV_X1    g741(.A(G224), .ZN(new_n928));
  OAI21_X1  g742(.A(G953), .B1(new_n602), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n822), .A2(new_n832), .A3(new_n831), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n929), .B1(new_n931), .B2(G953), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n872), .B1(G898), .B2(new_n263), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT123), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n932), .B(new_n934), .ZN(G69));
  NOR3_X1   g749(.A1(new_n736), .A2(new_n661), .A3(new_n668), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n755), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n762), .A2(new_n739), .A3(new_n769), .A4(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n663), .A2(new_n689), .A3(new_n725), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT124), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n742), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n263), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n263), .A2(G900), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT125), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n232), .B1(new_n259), .B2(KEYINPUT30), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n521), .A2(new_n522), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n684), .A2(new_n940), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT62), .Z(new_n951));
  AND2_X1   g765(.A1(new_n762), .A2(new_n769), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n693), .A2(new_n682), .A3(new_n729), .A4(new_n806), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n954), .A2(new_n263), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n949), .B1(new_n955), .B2(new_n948), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n948), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(G227), .A2(G900), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n958), .A2(G953), .A3(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n956), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n960), .B(new_n949), .C1(new_n955), .C2(new_n948), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(G72));
  NAND2_X1  g778(.A1(new_n260), .A2(new_n261), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT127), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n938), .A2(new_n930), .A3(new_n941), .ZN(new_n967));
  NAND2_X1  g781(.A1(G472), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT63), .Z(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n292), .B(new_n966), .C1(new_n967), .C2(new_n970), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n951), .A2(new_n931), .A3(new_n952), .A4(new_n953), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n969), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n268), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n880), .B(new_n971), .C1(new_n974), .C2(new_n966), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n847), .A2(new_n848), .ZN(new_n976));
  AOI211_X1 g790(.A(new_n970), .B(new_n976), .C1(new_n269), .C2(new_n295), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n975), .A2(new_n977), .ZN(G57));
endmodule


