

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599;

  AND2_X1 U326 ( .A1(G226GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U327 ( .A(n350), .B(KEYINPUT98), .ZN(n351) );
  XNOR2_X1 U328 ( .A(n473), .B(KEYINPUT110), .ZN(n474) );
  INV_X1 U329 ( .A(KEYINPUT32), .ZN(n423) );
  XNOR2_X1 U330 ( .A(n475), .B(n474), .ZN(n478) );
  XNOR2_X1 U331 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U332 ( .A(n403), .B(n294), .ZN(n338) );
  XNOR2_X1 U333 ( .A(n426), .B(n425), .ZN(n429) );
  XNOR2_X1 U334 ( .A(n437), .B(n338), .ZN(n339) );
  XNOR2_X1 U335 ( .A(KEYINPUT114), .B(KEYINPUT48), .ZN(n483) );
  XNOR2_X1 U336 ( .A(n341), .B(KEYINPUT96), .ZN(n342) );
  XNOR2_X1 U337 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U338 ( .A(n484), .B(n483), .ZN(n538) );
  XNOR2_X1 U339 ( .A(n343), .B(n342), .ZN(n345) );
  XNOR2_X1 U340 ( .A(n436), .B(n435), .ZN(n440) );
  NOR2_X1 U341 ( .A1(n517), .A2(n486), .ZN(n582) );
  XNOR2_X1 U342 ( .A(n444), .B(n443), .ZN(n589) );
  INV_X1 U343 ( .A(G190GAT), .ZN(n490) );
  XNOR2_X1 U344 ( .A(n465), .B(n464), .ZN(n512) );
  XNOR2_X1 U345 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U346 ( .A(n466), .B(G43GAT), .ZN(n467) );
  XNOR2_X1 U347 ( .A(n493), .B(n492), .ZN(G1351GAT) );
  XNOR2_X1 U348 ( .A(n468), .B(n467), .ZN(G1330GAT) );
  XOR2_X1 U349 ( .A(KEYINPUT104), .B(KEYINPUT38), .Z(n465) );
  XOR2_X1 U350 ( .A(KEYINPUT37), .B(KEYINPUT103), .Z(n422) );
  XOR2_X1 U351 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n296) );
  XNOR2_X1 U352 ( .A(KEYINPUT18), .B(G169GAT), .ZN(n295) );
  XNOR2_X1 U353 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U354 ( .A(KEYINPUT84), .B(n297), .ZN(n346) );
  XOR2_X1 U355 ( .A(G176GAT), .B(G71GAT), .Z(n299) );
  XNOR2_X1 U356 ( .A(G120GAT), .B(G15GAT), .ZN(n298) );
  XNOR2_X1 U357 ( .A(n299), .B(n298), .ZN(n314) );
  XOR2_X1 U358 ( .A(KEYINPUT82), .B(G190GAT), .Z(n301) );
  XNOR2_X1 U359 ( .A(G127GAT), .B(G99GAT), .ZN(n300) );
  XNOR2_X1 U360 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U361 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n303) );
  XNOR2_X1 U362 ( .A(G183GAT), .B(KEYINPUT81), .ZN(n302) );
  XNOR2_X1 U363 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U364 ( .A(n305), .B(n304), .Z(n312) );
  XOR2_X1 U365 ( .A(G113GAT), .B(KEYINPUT0), .Z(n307) );
  XNOR2_X1 U366 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n306) );
  XNOR2_X1 U367 ( .A(n307), .B(n306), .ZN(n361) );
  XOR2_X1 U368 ( .A(G43GAT), .B(G134GAT), .Z(n309) );
  NAND2_X1 U369 ( .A1(G227GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U370 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n361), .B(n310), .ZN(n311) );
  XNOR2_X1 U372 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U373 ( .A(n314), .B(n313), .Z(n315) );
  XOR2_X1 U374 ( .A(n346), .B(n315), .Z(n532) );
  INV_X1 U375 ( .A(n532), .ZN(n541) );
  XOR2_X1 U376 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n317) );
  XNOR2_X1 U377 ( .A(G155GAT), .B(G204GAT), .ZN(n316) );
  XNOR2_X1 U378 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U379 ( .A(G106GAT), .B(G78GAT), .Z(n433) );
  XOR2_X1 U380 ( .A(n318), .B(n433), .Z(n320) );
  XNOR2_X1 U381 ( .A(G148GAT), .B(G22GAT), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n320), .B(n319), .ZN(n325) );
  XNOR2_X1 U383 ( .A(G211GAT), .B(G197GAT), .ZN(n321) );
  XNOR2_X1 U384 ( .A(n321), .B(KEYINPUT21), .ZN(n340) );
  XOR2_X1 U385 ( .A(G218GAT), .B(G50GAT), .Z(n402) );
  XOR2_X1 U386 ( .A(n340), .B(n402), .Z(n323) );
  NAND2_X1 U387 ( .A1(G228GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U388 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U389 ( .A(n325), .B(n324), .Z(n334) );
  XNOR2_X1 U390 ( .A(KEYINPUT87), .B(KEYINPUT88), .ZN(n326) );
  XNOR2_X1 U391 ( .A(n326), .B(KEYINPUT2), .ZN(n327) );
  XOR2_X1 U392 ( .A(n327), .B(KEYINPUT3), .Z(n329) );
  XNOR2_X1 U393 ( .A(G141GAT), .B(G162GAT), .ZN(n328) );
  XNOR2_X1 U394 ( .A(n329), .B(n328), .ZN(n371) );
  XOR2_X1 U395 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n331) );
  XNOR2_X1 U396 ( .A(KEYINPUT89), .B(KEYINPUT85), .ZN(n330) );
  XNOR2_X1 U397 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U398 ( .A(n371), .B(n332), .ZN(n333) );
  XNOR2_X1 U399 ( .A(n334), .B(n333), .ZN(n487) );
  NOR2_X1 U400 ( .A1(n541), .A2(n487), .ZN(n335) );
  XOR2_X1 U401 ( .A(KEYINPUT26), .B(n335), .Z(n555) );
  INV_X1 U402 ( .A(n555), .ZN(n581) );
  XOR2_X1 U403 ( .A(G204GAT), .B(G176GAT), .Z(n337) );
  XNOR2_X1 U404 ( .A(G92GAT), .B(G64GAT), .ZN(n336) );
  XNOR2_X1 U405 ( .A(n337), .B(n336), .ZN(n437) );
  XOR2_X1 U406 ( .A(G190GAT), .B(G36GAT), .Z(n403) );
  XOR2_X1 U407 ( .A(n339), .B(KEYINPUT95), .Z(n343) );
  XNOR2_X1 U408 ( .A(n340), .B(KEYINPUT94), .ZN(n341) );
  XOR2_X1 U409 ( .A(G183GAT), .B(G8GAT), .Z(n385) );
  XOR2_X1 U410 ( .A(G218GAT), .B(n385), .Z(n344) );
  XNOR2_X1 U411 ( .A(n345), .B(n344), .ZN(n347) );
  XNOR2_X1 U412 ( .A(n347), .B(n346), .ZN(n349) );
  INV_X1 U413 ( .A(n349), .ZN(n530) );
  XOR2_X1 U414 ( .A(KEYINPUT27), .B(KEYINPUT97), .Z(n348) );
  XOR2_X1 U415 ( .A(n530), .B(n348), .Z(n374) );
  NAND2_X1 U416 ( .A1(n581), .A2(n374), .ZN(n354) );
  NAND2_X1 U417 ( .A1(n349), .A2(n541), .ZN(n350) );
  NAND2_X1 U418 ( .A1(n351), .A2(n487), .ZN(n352) );
  XOR2_X1 U419 ( .A(KEYINPUT25), .B(n352), .Z(n353) );
  NAND2_X1 U420 ( .A1(n354), .A2(n353), .ZN(n372) );
  XOR2_X1 U421 ( .A(KEYINPUT5), .B(KEYINPUT91), .Z(n356) );
  XNOR2_X1 U422 ( .A(G85GAT), .B(KEYINPUT6), .ZN(n355) );
  XNOR2_X1 U423 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U424 ( .A(KEYINPUT92), .B(KEYINPUT4), .Z(n358) );
  XNOR2_X1 U425 ( .A(KEYINPUT1), .B(KEYINPUT90), .ZN(n357) );
  XNOR2_X1 U426 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U427 ( .A(n360), .B(n359), .Z(n369) );
  XOR2_X1 U428 ( .A(n361), .B(G57GAT), .Z(n363) );
  NAND2_X1 U429 ( .A1(G225GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U430 ( .A(n363), .B(n362), .ZN(n367) );
  XNOR2_X1 U431 ( .A(G29GAT), .B(G134GAT), .ZN(n417) );
  XOR2_X1 U432 ( .A(G120GAT), .B(G148GAT), .Z(n432) );
  XOR2_X1 U433 ( .A(n417), .B(n432), .Z(n365) );
  XNOR2_X1 U434 ( .A(G127GAT), .B(G155GAT), .ZN(n364) );
  XNOR2_X1 U435 ( .A(n364), .B(G1GAT), .ZN(n387) );
  XNOR2_X1 U436 ( .A(n365), .B(n387), .ZN(n366) );
  XNOR2_X1 U437 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U438 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U439 ( .A(n371), .B(n370), .ZN(n373) );
  NAND2_X1 U440 ( .A1(n372), .A2(n373), .ZN(n377) );
  XOR2_X1 U441 ( .A(KEYINPUT93), .B(n373), .Z(n528) );
  INV_X1 U442 ( .A(n528), .ZN(n517) );
  AND2_X1 U443 ( .A1(n374), .A2(n517), .ZN(n539) );
  XNOR2_X1 U444 ( .A(n487), .B(KEYINPUT28), .ZN(n535) );
  INV_X1 U445 ( .A(n535), .ZN(n540) );
  NOR2_X1 U446 ( .A1(n540), .A2(n541), .ZN(n375) );
  NAND2_X1 U447 ( .A1(n539), .A2(n375), .ZN(n376) );
  NAND2_X1 U448 ( .A1(n377), .A2(n376), .ZN(n378) );
  XOR2_X1 U449 ( .A(KEYINPUT99), .B(n378), .Z(n497) );
  XOR2_X1 U450 ( .A(G15GAT), .B(G22GAT), .Z(n448) );
  INV_X1 U451 ( .A(KEYINPUT67), .ZN(n379) );
  NAND2_X1 U452 ( .A1(n379), .A2(KEYINPUT13), .ZN(n382) );
  INV_X1 U453 ( .A(KEYINPUT13), .ZN(n380) );
  NAND2_X1 U454 ( .A1(n380), .A2(KEYINPUT67), .ZN(n381) );
  NAND2_X1 U455 ( .A1(n382), .A2(n381), .ZN(n384) );
  XNOR2_X1 U456 ( .A(G57GAT), .B(G71GAT), .ZN(n383) );
  XNOR2_X1 U457 ( .A(n384), .B(n383), .ZN(n426) );
  XNOR2_X1 U458 ( .A(n448), .B(n426), .ZN(n386) );
  XNOR2_X1 U459 ( .A(n386), .B(n385), .ZN(n391) );
  XOR2_X1 U460 ( .A(n387), .B(G64GAT), .Z(n389) );
  NAND2_X1 U461 ( .A1(G231GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U462 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U463 ( .A(n391), .B(n390), .Z(n399) );
  XOR2_X1 U464 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n393) );
  XNOR2_X1 U465 ( .A(G211GAT), .B(G78GAT), .ZN(n392) );
  XNOR2_X1 U466 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U467 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n395) );
  XNOR2_X1 U468 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n394) );
  XNOR2_X1 U469 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U470 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U471 ( .A(n399), .B(n398), .Z(n592) );
  INV_X1 U472 ( .A(n592), .ZN(n400) );
  AND2_X1 U473 ( .A1(n497), .A2(n400), .ZN(n401) );
  XNOR2_X1 U474 ( .A(n401), .B(KEYINPUT102), .ZN(n420) );
  INV_X1 U475 ( .A(KEYINPUT36), .ZN(n419) );
  XOR2_X1 U476 ( .A(n403), .B(n402), .Z(n405) );
  NAND2_X1 U477 ( .A1(G232GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U478 ( .A(n405), .B(n404), .ZN(n416) );
  XOR2_X1 U479 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n411) );
  XOR2_X1 U480 ( .A(KEYINPUT11), .B(KEYINPUT73), .Z(n407) );
  XNOR2_X1 U481 ( .A(G162GAT), .B(G92GAT), .ZN(n406) );
  XNOR2_X1 U482 ( .A(n407), .B(n406), .ZN(n409) );
  XNOR2_X1 U483 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n408) );
  XNOR2_X1 U484 ( .A(n408), .B(KEYINPUT7), .ZN(n452) );
  XNOR2_X1 U485 ( .A(n409), .B(n452), .ZN(n410) );
  XNOR2_X1 U486 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U487 ( .A(G85GAT), .B(G99GAT), .Z(n438) );
  XOR2_X1 U488 ( .A(n412), .B(n438), .Z(n414) );
  XNOR2_X1 U489 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n413) );
  XNOR2_X1 U490 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U491 ( .A(n416), .B(n415), .ZN(n418) );
  XOR2_X1 U492 ( .A(n418), .B(n417), .Z(n494) );
  XNOR2_X1 U493 ( .A(n419), .B(n494), .ZN(n595) );
  NAND2_X1 U494 ( .A1(n420), .A2(n595), .ZN(n421) );
  XNOR2_X1 U495 ( .A(n422), .B(n421), .ZN(n527) );
  NAND2_X1 U496 ( .A1(G230GAT), .A2(G233GAT), .ZN(n424) );
  INV_X1 U497 ( .A(n429), .ZN(n428) );
  INV_X1 U498 ( .A(KEYINPUT71), .ZN(n427) );
  NAND2_X1 U499 ( .A1(n428), .A2(n427), .ZN(n431) );
  NAND2_X1 U500 ( .A1(n429), .A2(KEYINPUT71), .ZN(n430) );
  NAND2_X1 U501 ( .A1(n431), .A2(n430), .ZN(n436) );
  XOR2_X1 U502 ( .A(n432), .B(KEYINPUT68), .Z(n434) );
  XOR2_X1 U503 ( .A(n438), .B(n437), .Z(n439) );
  XNOR2_X1 U504 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U505 ( .A(KEYINPUT70), .B(KEYINPUT31), .Z(n442) );
  XNOR2_X1 U506 ( .A(KEYINPUT33), .B(KEYINPUT69), .ZN(n441) );
  XNOR2_X1 U507 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U508 ( .A(G36GAT), .B(G50GAT), .Z(n446) );
  XNOR2_X1 U509 ( .A(G29GAT), .B(G113GAT), .ZN(n445) );
  XNOR2_X1 U510 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U511 ( .A(n448), .B(n447), .Z(n450) );
  NAND2_X1 U512 ( .A1(G229GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U513 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U514 ( .A(n451), .B(KEYINPUT30), .Z(n454) );
  XNOR2_X1 U515 ( .A(n452), .B(KEYINPUT29), .ZN(n453) );
  XNOR2_X1 U516 ( .A(n454), .B(n453), .ZN(n462) );
  XOR2_X1 U517 ( .A(G197GAT), .B(G169GAT), .Z(n456) );
  XNOR2_X1 U518 ( .A(G141GAT), .B(G1GAT), .ZN(n455) );
  XNOR2_X1 U519 ( .A(n456), .B(n455), .ZN(n460) );
  XOR2_X1 U520 ( .A(KEYINPUT64), .B(KEYINPUT66), .Z(n458) );
  XNOR2_X1 U521 ( .A(G8GAT), .B(KEYINPUT65), .ZN(n457) );
  XNOR2_X1 U522 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U523 ( .A(n460), .B(n459), .Z(n461) );
  XOR2_X1 U524 ( .A(n462), .B(n461), .Z(n558) );
  INV_X1 U525 ( .A(n558), .ZN(n583) );
  NOR2_X1 U526 ( .A1(n589), .A2(n583), .ZN(n463) );
  XNOR2_X1 U527 ( .A(n463), .B(KEYINPUT72), .ZN(n499) );
  NAND2_X1 U528 ( .A1(n527), .A2(n499), .ZN(n464) );
  NAND2_X1 U529 ( .A1(n512), .A2(n541), .ZN(n468) );
  XOR2_X1 U530 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n466) );
  NAND2_X1 U531 ( .A1(n595), .A2(n592), .ZN(n469) );
  XOR2_X1 U532 ( .A(KEYINPUT45), .B(n469), .Z(n470) );
  NAND2_X1 U533 ( .A1(n470), .A2(n583), .ZN(n471) );
  NOR2_X1 U534 ( .A1(n589), .A2(n471), .ZN(n472) );
  XNOR2_X1 U535 ( .A(KEYINPUT113), .B(n472), .ZN(n482) );
  XNOR2_X1 U536 ( .A(KEYINPUT41), .B(n589), .ZN(n514) );
  NOR2_X1 U537 ( .A1(n514), .A2(n583), .ZN(n475) );
  XNOR2_X1 U538 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n473) );
  INV_X1 U539 ( .A(n494), .ZN(n568) );
  XNOR2_X1 U540 ( .A(n592), .B(KEYINPUT109), .ZN(n579) );
  INV_X1 U541 ( .A(n579), .ZN(n476) );
  NOR2_X1 U542 ( .A1(n568), .A2(n476), .ZN(n477) );
  AND2_X1 U543 ( .A1(n478), .A2(n477), .ZN(n480) );
  XNOR2_X1 U544 ( .A(KEYINPUT47), .B(KEYINPUT112), .ZN(n479) );
  XNOR2_X1 U545 ( .A(n480), .B(n479), .ZN(n481) );
  NAND2_X1 U546 ( .A1(n482), .A2(n481), .ZN(n484) );
  NAND2_X1 U547 ( .A1(n349), .A2(n538), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n485), .B(KEYINPUT54), .ZN(n486) );
  NAND2_X1 U549 ( .A1(n487), .A2(n582), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n488), .B(KEYINPUT55), .ZN(n489) );
  NAND2_X1 U551 ( .A1(n489), .A2(n541), .ZN(n578) );
  NOR2_X1 U552 ( .A1(n578), .A2(n494), .ZN(n493) );
  XNOR2_X1 U553 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n491) );
  XNOR2_X1 U554 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n502) );
  XOR2_X1 U555 ( .A(KEYINPUT16), .B(KEYINPUT78), .Z(n496) );
  NAND2_X1 U556 ( .A1(n494), .A2(n592), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(n498) );
  AND2_X1 U558 ( .A1(n498), .A2(n497), .ZN(n515) );
  NAND2_X1 U559 ( .A1(n515), .A2(n499), .ZN(n500) );
  XOR2_X1 U560 ( .A(KEYINPUT100), .B(n500), .Z(n506) );
  NAND2_X1 U561 ( .A1(n517), .A2(n506), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(G1324GAT) );
  NAND2_X1 U563 ( .A1(n506), .A2(n349), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n503), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U565 ( .A(G15GAT), .B(KEYINPUT35), .Z(n505) );
  NAND2_X1 U566 ( .A1(n541), .A2(n506), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(G1326GAT) );
  XOR2_X1 U568 ( .A(G22GAT), .B(KEYINPUT101), .Z(n508) );
  NAND2_X1 U569 ( .A1(n540), .A2(n506), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n508), .B(n507), .ZN(G1327GAT) );
  XOR2_X1 U571 ( .A(G29GAT), .B(KEYINPUT39), .Z(n510) );
  NAND2_X1 U572 ( .A1(n512), .A2(n517), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(G1328GAT) );
  NAND2_X1 U574 ( .A1(n512), .A2(n349), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U576 ( .A1(n512), .A2(n540), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n513), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U578 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n519) );
  XNOR2_X1 U579 ( .A(n514), .B(KEYINPUT106), .ZN(n572) );
  NOR2_X1 U580 ( .A1(n558), .A2(n572), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n515), .A2(n526), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n516), .B(KEYINPUT107), .ZN(n523) );
  NAND2_X1 U583 ( .A1(n517), .A2(n523), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(G1332GAT) );
  NAND2_X1 U585 ( .A1(n523), .A2(n349), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n520), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U587 ( .A1(n523), .A2(n541), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(KEYINPUT108), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G71GAT), .B(n522), .ZN(G1334GAT) );
  XOR2_X1 U590 ( .A(G78GAT), .B(KEYINPUT43), .Z(n525) );
  NAND2_X1 U591 ( .A1(n523), .A2(n540), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(G1335GAT) );
  NAND2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n534) );
  NOR2_X1 U594 ( .A1(n528), .A2(n534), .ZN(n529) );
  XOR2_X1 U595 ( .A(G85GAT), .B(n529), .Z(G1336GAT) );
  NOR2_X1 U596 ( .A1(n530), .A2(n534), .ZN(n531) );
  XOR2_X1 U597 ( .A(G92GAT), .B(n531), .Z(G1337GAT) );
  NOR2_X1 U598 ( .A1(n532), .A2(n534), .ZN(n533) );
  XOR2_X1 U599 ( .A(G99GAT), .B(n533), .Z(G1338GAT) );
  NOR2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U601 ( .A(G106GAT), .B(n536), .Z(n537) );
  XNOR2_X1 U602 ( .A(KEYINPUT44), .B(n537), .ZN(G1339GAT) );
  NAND2_X1 U603 ( .A1(n539), .A2(n538), .ZN(n556) );
  NOR2_X1 U604 ( .A1(n540), .A2(n556), .ZN(n542) );
  NAND2_X1 U605 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U606 ( .A(n543), .B(KEYINPUT115), .Z(n547) );
  INV_X1 U607 ( .A(n547), .ZN(n551) );
  NAND2_X1 U608 ( .A1(n551), .A2(n558), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n544), .B(G113GAT), .ZN(G1340GAT) );
  NOR2_X1 U610 ( .A1(n572), .A2(n547), .ZN(n546) );
  XNOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1341GAT) );
  NOR2_X1 U613 ( .A1(n579), .A2(n547), .ZN(n549) );
  XNOR2_X1 U614 ( .A(KEYINPUT116), .B(KEYINPUT50), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U616 ( .A(G127GAT), .B(n550), .Z(G1342GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n553) );
  NAND2_X1 U618 ( .A1(n551), .A2(n568), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U620 ( .A(G134GAT), .B(n554), .Z(G1343GAT) );
  XOR2_X1 U621 ( .A(G141GAT), .B(KEYINPUT119), .Z(n560) );
  NOR2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U623 ( .A(n557), .B(KEYINPUT118), .Z(n563) );
  INV_X1 U624 ( .A(n563), .ZN(n569) );
  NAND2_X1 U625 ( .A1(n558), .A2(n569), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1344GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n562) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n565) );
  NOR2_X1 U630 ( .A1(n514), .A2(n563), .ZN(n564) );
  XOR2_X1 U631 ( .A(n565), .B(n564), .Z(G1345GAT) );
  XOR2_X1 U632 ( .A(G155GAT), .B(KEYINPUT121), .Z(n567) );
  NAND2_X1 U633 ( .A1(n569), .A2(n592), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G1346GAT) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U637 ( .A1(n583), .A2(n578), .ZN(n571) );
  XOR2_X1 U638 ( .A(G169GAT), .B(n571), .Z(G1348GAT) );
  NOR2_X1 U639 ( .A1(n578), .A2(n572), .ZN(n577) );
  XOR2_X1 U640 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n574) );
  XNOR2_X1 U641 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n573) );
  XNOR2_X1 U642 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U643 ( .A(KEYINPUT56), .B(n575), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n577), .B(n576), .ZN(G1349GAT) );
  NOR2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U646 ( .A(G183GAT), .B(n580), .Z(G1350GAT) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n588) );
  NOR2_X1 U648 ( .A1(n588), .A2(n583), .ZN(n587) );
  XOR2_X1 U649 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n585) );
  XNOR2_X1 U650 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1352GAT) );
  XOR2_X1 U653 ( .A(G204GAT), .B(KEYINPUT61), .Z(n591) );
  INV_X1 U654 ( .A(n588), .ZN(n596) );
  NAND2_X1 U655 ( .A1(n596), .A2(n589), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n591), .B(n590), .ZN(G1353GAT) );
  NAND2_X1 U657 ( .A1(n592), .A2(n596), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n593), .B(KEYINPUT126), .ZN(n594) );
  XNOR2_X1 U659 ( .A(G211GAT), .B(n594), .ZN(G1354GAT) );
  XOR2_X1 U660 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n598) );
  NAND2_X1 U661 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U662 ( .A(n598), .B(n597), .ZN(n599) );
  XNOR2_X1 U663 ( .A(G218GAT), .B(n599), .ZN(G1355GAT) );
endmodule

