//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G210), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT27), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(KEYINPUT1), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  OAI22_X1  g011(.A1(new_n193), .A2(new_n195), .B1(new_n197), .B2(G128), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G143), .B(G146), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT64), .B1(new_n200), .B2(new_n193), .ZN(new_n201));
  AND4_X1   g015(.A1(KEYINPUT64), .A2(new_n193), .A3(new_n195), .A4(new_n197), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n199), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G137), .ZN(new_n206));
  INV_X1    g020(.A(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT11), .A3(G134), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(G137), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n206), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n205), .A2(G137), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n207), .A2(G134), .ZN(new_n213));
  OAI21_X1  g027(.A(G131), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n203), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n218));
  NOR3_X1   g032(.A1(new_n218), .A2(KEYINPUT2), .A3(G113), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT2), .ZN(new_n220));
  INV_X1    g034(.A(G113), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT65), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI22_X1  g036(.A1(new_n219), .A2(new_n222), .B1(new_n220), .B2(new_n221), .ZN(new_n223));
  XNOR2_X1  g037(.A(G116), .B(G119), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  OAI221_X1 g040(.A(new_n224), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n219), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n206), .A2(new_n208), .A3(new_n210), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G131), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n211), .ZN(new_n232));
  AND2_X1   g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n195), .A2(new_n197), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT0), .B(G128), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n234), .B1(new_n200), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n217), .A2(new_n229), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n217), .A2(new_n238), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(new_n228), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n193), .A2(new_n195), .A3(new_n197), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n200), .A2(KEYINPUT64), .A3(new_n193), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n215), .B1(new_n247), .B2(new_n199), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n236), .B1(new_n211), .B2(new_n231), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n240), .B(new_n228), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n239), .B1(new_n242), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT28), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT28), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n239), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n191), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n257));
  INV_X1    g071(.A(new_n239), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT30), .B1(new_n248), .B2(new_n249), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT30), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n217), .A2(new_n260), .A3(new_n238), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n258), .B1(new_n262), .B2(new_n228), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n257), .B1(new_n263), .B2(new_n191), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n229), .B1(new_n259), .B2(new_n261), .ZN(new_n265));
  INV_X1    g079(.A(new_n191), .ZN(new_n266));
  NOR4_X1   g080(.A1(new_n265), .A2(new_n258), .A3(KEYINPUT66), .A4(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT31), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n260), .B1(new_n217), .B2(new_n238), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n248), .A2(new_n249), .A3(KEYINPUT30), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n228), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(new_n239), .A3(new_n191), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n256), .B1(new_n268), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(G472), .A2(G902), .ZN(new_n276));
  XOR2_X1   g090(.A(new_n276), .B(KEYINPUT68), .Z(new_n277));
  OAI21_X1  g091(.A(KEYINPUT32), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n253), .A2(new_n255), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n266), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n272), .A2(KEYINPUT66), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n263), .A2(new_n257), .A3(new_n191), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n273), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n274), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n280), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT32), .ZN(new_n286));
  INV_X1    g100(.A(new_n277), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n266), .B1(new_n265), .B2(new_n258), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT29), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n289), .B(new_n290), .C1(new_n279), .C2(new_n266), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n241), .A2(new_n228), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n254), .B1(new_n292), .B2(new_n239), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT69), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT69), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n255), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n294), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n266), .A2(new_n290), .ZN(new_n298));
  AOI21_X1  g112(.A(G902), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n291), .A2(new_n299), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n278), .A2(new_n288), .B1(G472), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G217), .ZN(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n302), .B1(G234), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT80), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n308));
  INV_X1    g122(.A(G119), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n308), .B1(new_n309), .B2(G128), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(G128), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(KEYINPUT23), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT23), .B1(new_n192), .B2(G119), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT72), .B1(new_n192), .B2(G119), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n315), .A3(KEYINPUT73), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G110), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT73), .B1(new_n312), .B2(new_n315), .ZN(new_n318));
  OR2_X1    g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(G125), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n322), .B1(new_n326), .B2(new_n320), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n196), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n329));
  OAI211_X1 g143(.A(G146), .B(new_n322), .C1(new_n326), .C2(new_n320), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT70), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n332), .B1(new_n309), .B2(G128), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n192), .A2(KEYINPUT70), .A3(G119), .ZN(new_n334));
  OAI22_X1  g148(.A1(new_n333), .A2(new_n334), .B1(new_n309), .B2(G128), .ZN(new_n335));
  INV_X1    g149(.A(G110), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT24), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT24), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G110), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT71), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n337), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n340), .B1(new_n337), .B2(new_n339), .ZN(new_n342));
  OR3_X1    g156(.A1(new_n335), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n327), .A2(KEYINPUT74), .A3(new_n196), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n319), .A2(new_n331), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n312), .A2(new_n315), .A3(new_n336), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT75), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n335), .B1(new_n341), .B2(new_n342), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n312), .A2(new_n315), .A3(KEYINPUT75), .A4(new_n336), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n327), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n353));
  AOI21_X1  g167(.A(G146), .B1(new_n326), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G125), .B(G140), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT76), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n352), .A2(G146), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n351), .A2(KEYINPUT77), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT77), .B1(new_n351), .B2(new_n357), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n345), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT22), .B(G137), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(KEYINPUT78), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT79), .ZN(new_n363));
  INV_X1    g177(.A(G953), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n364), .A2(G221), .A3(G234), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n361), .A2(KEYINPUT78), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n361), .A2(KEYINPUT78), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n363), .A2(new_n365), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n365), .B1(new_n363), .B2(new_n369), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n360), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n372), .B(new_n345), .C1(new_n359), .C2(new_n358), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(G902), .B1(new_n305), .B2(new_n306), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n307), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n377), .ZN(new_n379));
  INV_X1    g193(.A(new_n307), .ZN(new_n380));
  AOI211_X1 g194(.A(new_n379), .B(new_n380), .C1(new_n374), .C2(new_n375), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n304), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(KEYINPUT81), .B(new_n304), .C1(new_n378), .C2(new_n381), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n304), .A2(G902), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n376), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n301), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G221), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT9), .B(G234), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n390), .B1(new_n392), .B2(new_n303), .ZN(new_n393));
  INV_X1    g207(.A(G469), .ZN(new_n394));
  INV_X1    g208(.A(G104), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT3), .B1(new_n395), .B2(G107), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n397));
  INV_X1    g211(.A(G107), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(G104), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(G107), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT82), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n396), .A2(new_n399), .A3(new_n403), .A4(new_n400), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(G101), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G101), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n396), .A2(new_n399), .A3(new_n406), .A4(new_n400), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(KEYINPUT4), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n402), .A2(new_n409), .A3(G101), .A4(new_n404), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n237), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n198), .B1(new_n245), .B2(new_n246), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n395), .A2(G107), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n398), .A2(G104), .ZN(new_n414));
  OAI21_X1  g228(.A(G101), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n407), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT10), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT10), .ZN(new_n418));
  INV_X1    g232(.A(new_n416), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n203), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n232), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n411), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G140), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n364), .A2(G227), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n203), .A2(new_n419), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n412), .A2(new_n416), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n232), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT12), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n430), .A2(new_n431), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n423), .B(new_n427), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n411), .A2(new_n421), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n232), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n427), .B1(new_n436), .B2(new_n423), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT83), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n434), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n411), .A2(new_n421), .A3(new_n422), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n422), .B1(new_n411), .B2(new_n421), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n438), .B(new_n426), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n394), .B(new_n303), .C1(new_n439), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT84), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n426), .B1(new_n440), .B2(new_n441), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT83), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n442), .A3(new_n434), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT84), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n394), .A4(new_n303), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n430), .B(new_n431), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n423), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n426), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n440), .A2(new_n426), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n436), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n394), .B1(new_n457), .B2(new_n303), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n393), .B1(new_n451), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(G214), .B1(G237), .B2(G902), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n463));
  INV_X1    g277(.A(G116), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(G119), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT5), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n221), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n309), .A2(G116), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(G119), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT5), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n467), .A2(KEYINPUT85), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT85), .B1(new_n467), .B2(new_n470), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n419), .B(new_n227), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n228), .A2(new_n410), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n407), .A2(KEYINPUT4), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n406), .B1(new_n401), .B2(KEYINPUT82), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n477), .B2(new_n404), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n474), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(G110), .B(G122), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n463), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n408), .A2(new_n228), .A3(new_n410), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n480), .A3(new_n474), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n234), .B(G125), .C1(new_n200), .C2(new_n235), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n412), .B2(G125), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT87), .B(G224), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n364), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n487), .B(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n480), .B1(new_n483), .B2(new_n474), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT86), .B1(new_n491), .B2(new_n463), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n479), .A2(KEYINPUT86), .A3(new_n463), .A4(new_n481), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n485), .B(new_n490), .C1(new_n492), .C2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n480), .B(KEYINPUT8), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n467), .A2(new_n470), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT85), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n471), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n419), .B1(new_n500), .B2(new_n227), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n419), .A2(new_n227), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n470), .A2(KEYINPUT88), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n467), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n470), .A2(KEYINPUT88), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n496), .B1(new_n501), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n489), .A2(KEYINPUT7), .ZN(new_n509));
  NAND2_X1  g323(.A1(KEYINPUT89), .A2(KEYINPUT7), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(new_n487), .B2(new_n510), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n487), .A2(new_n509), .A3(new_n510), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n484), .B(new_n508), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n513), .A2(new_n303), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n495), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT90), .ZN(new_n516));
  OAI21_X1  g330(.A(G210), .B1(G237), .B2(G902), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT90), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n495), .A2(new_n514), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n516), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n495), .A2(new_n514), .A3(new_n517), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n462), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(G113), .B(G122), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(new_n395), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n196), .B1(new_n355), .B2(KEYINPUT76), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n326), .A2(new_n353), .ZN(new_n527));
  OAI22_X1  g341(.A1(new_n526), .A2(new_n527), .B1(new_n196), .B2(new_n355), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n187), .A2(G214), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n194), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n531));
  NAND2_X1  g345(.A1(KEYINPUT18), .A2(G131), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n530), .A2(new_n531), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(KEYINPUT18), .A3(G131), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n528), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n331), .A2(new_n344), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n209), .B1(new_n530), .B2(new_n531), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT17), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n534), .A2(G131), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n530), .A2(new_n209), .A3(new_n531), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n539), .B1(new_n542), .B2(KEYINPUT17), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n525), .B(new_n536), .C1(new_n537), .C2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n355), .B2(KEYINPUT76), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT19), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n353), .B1(new_n547), .B2(KEYINPUT91), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n546), .A2(new_n547), .B1(new_n355), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(G146), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n530), .A2(new_n209), .A3(new_n531), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n330), .B1(new_n551), .B2(new_n538), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n536), .B(KEYINPUT92), .C1(new_n550), .C2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n525), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n542), .B(new_n330), .C1(G146), .C2(new_n549), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT92), .B1(new_n556), .B2(new_n536), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n544), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT93), .ZN(new_n559));
  NOR2_X1   g373(.A1(G475), .A2(G902), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT93), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n544), .B(new_n561), .C1(new_n555), .C2(new_n557), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT20), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT20), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n558), .A2(new_n565), .A3(new_n560), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n536), .B1(new_n537), .B2(new_n543), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n554), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n544), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n303), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n572), .A2(G475), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n391), .A2(new_n302), .A3(G953), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT94), .ZN(new_n577));
  INV_X1    g391(.A(G122), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n577), .B1(new_n578), .B2(G116), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n464), .A2(KEYINPUT94), .A3(G122), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(G116), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n398), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n194), .A2(G128), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n192), .A2(G143), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n205), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n584), .A2(new_n585), .A3(G134), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n581), .A2(KEYINPUT14), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT14), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n579), .A2(new_n591), .A3(new_n580), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n590), .A2(new_n582), .A3(new_n592), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n583), .B(new_n589), .C1(new_n593), .C2(new_n398), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT95), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT13), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n585), .A2(new_n596), .A3(G134), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n587), .A2(new_n588), .A3(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n584), .A2(new_n585), .A3(new_n596), .A4(G134), .ZN(new_n599));
  INV_X1    g413(.A(new_n583), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n398), .B1(new_n581), .B2(new_n582), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n598), .B(new_n599), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n594), .A2(new_n595), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n595), .B1(new_n594), .B2(new_n602), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n576), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n594), .A2(new_n602), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT95), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n594), .A2(new_n595), .A3(new_n602), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n575), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n605), .A2(new_n609), .A3(new_n303), .ZN(new_n610));
  INV_X1    g424(.A(G478), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(KEYINPUT15), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n612), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n605), .A2(new_n609), .A3(new_n303), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(G234), .A2(G237), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(G952), .A3(new_n364), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT21), .B(G898), .Z(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(G902), .A3(G953), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(new_n620), .B(KEYINPUT96), .Z(new_n621));
  AND3_X1   g435(.A1(new_n613), .A2(new_n615), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n568), .A2(new_n574), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT97), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n566), .B1(new_n563), .B2(KEYINPUT20), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(new_n573), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n622), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n389), .A2(new_n460), .A3(new_n523), .A4(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT98), .B(G101), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT99), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n630), .B(new_n632), .ZN(G3));
  INV_X1    g447(.A(new_n388), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n285), .A2(new_n303), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n635), .A2(G472), .B1(new_n287), .B2(new_n285), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n460), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n621), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n611), .A2(G902), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n605), .A2(new_n609), .A3(KEYINPUT33), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT33), .B1(new_n605), .B2(new_n609), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n610), .A2(new_n611), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n645), .B1(new_n625), .B2(new_n573), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n517), .B1(new_n495), .B2(new_n514), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT100), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n461), .B(new_n522), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n513), .A2(new_n303), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n479), .A2(new_n463), .A3(new_n481), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT86), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n653), .A2(new_n493), .B1(new_n484), .B2(new_n482), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n650), .B1(new_n654), .B2(new_n490), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n655), .A2(KEYINPUT100), .A3(new_n461), .A4(new_n517), .ZN(new_n656));
  AOI211_X1 g470(.A(new_n639), .B(new_n646), .C1(new_n649), .C2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n638), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT34), .B(G104), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  AOI21_X1  g474(.A(new_n639), .B1(new_n649), .B2(new_n656), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n559), .A2(new_n565), .A3(new_n560), .A4(new_n562), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n573), .B1(new_n564), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n613), .A2(new_n615), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n661), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n666), .B1(new_n661), .B2(new_n665), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n638), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT35), .B(G107), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G9));
  NOR2_X1   g485(.A1(new_n372), .A2(KEYINPUT36), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(new_n360), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n386), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n384), .A2(new_n385), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n636), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n677), .A2(new_n460), .A3(new_n523), .A4(new_n629), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  AND3_X1   g494(.A1(new_n384), .A2(new_n385), .A3(new_n674), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n301), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n649), .A2(new_n656), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n619), .A2(G900), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n617), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n663), .A2(new_n664), .A3(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n682), .A2(new_n460), .A3(new_n683), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G128), .ZN(G30));
  OAI21_X1  g502(.A(new_n664), .B1(new_n625), .B2(new_n573), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n681), .A2(new_n461), .A3(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n692));
  OR2_X1    g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n278), .A2(new_n288), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n281), .A2(new_n282), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n191), .B1(new_n292), .B2(new_n239), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT102), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n303), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G472), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n691), .A2(new_n692), .B1(new_n694), .B2(new_n699), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n521), .A2(new_n522), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n701), .B(KEYINPUT38), .Z(new_n702));
  NAND3_X1  g516(.A1(new_n693), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT104), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT104), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n693), .A2(new_n700), .A3(new_n702), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n685), .B(KEYINPUT39), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n460), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT40), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n704), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G143), .ZN(G45));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n300), .A2(G472), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n275), .A2(KEYINPUT32), .A3(new_n277), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n286), .B1(new_n285), .B2(new_n287), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n683), .A3(new_n675), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n451), .A2(new_n459), .ZN(new_n718));
  INV_X1    g532(.A(new_n393), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n645), .B(new_n685), .C1(new_n625), .C2(new_n573), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n712), .B1(new_n717), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n458), .B1(new_n445), .B2(new_n450), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n724), .A2(new_n393), .A3(new_n720), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n682), .A2(KEYINPUT105), .A3(new_n725), .A4(new_n683), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G146), .ZN(G48));
  AOI22_X1  g542(.A1(new_n446), .A2(KEYINPUT83), .B1(new_n455), .B2(new_n452), .ZN(new_n729));
  AOI21_X1  g543(.A(G902), .B1(new_n729), .B2(new_n442), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n719), .B1(new_n730), .B2(new_n394), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n450), .B2(new_n445), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n657), .A2(new_n389), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT41), .B(G113), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G15));
  OAI211_X1 g549(.A(new_n389), .B(new_n732), .C1(new_n667), .C2(new_n668), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G116), .ZN(G18));
  INV_X1    g551(.A(new_n731), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n683), .A2(new_n738), .A3(new_n451), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n732), .A2(KEYINPUT106), .A3(new_n683), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n629), .A3(new_n682), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G119), .ZN(G21));
  OAI22_X1  g559(.A1(new_n283), .A2(new_n284), .B1(new_n191), .B2(new_n297), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n277), .B(KEYINPUT107), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n635), .A2(G472), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n388), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n689), .B1(new_n649), .B2(new_n656), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(new_n621), .A3(new_n732), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G122), .ZN(G24));
  NAND3_X1  g567(.A1(new_n748), .A2(new_n721), .A3(new_n675), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n754), .B1(new_n741), .B2(new_n742), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT108), .B(G125), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G27));
  AOI21_X1  g571(.A(new_n462), .B1(new_n655), .B2(new_n517), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n518), .B1(new_n655), .B2(new_n519), .ZN(new_n759));
  INV_X1    g573(.A(new_n520), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n719), .B(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(G469), .A2(G902), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n763), .B(KEYINPUT109), .Z(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n765), .B1(new_n457), .B2(new_n394), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n449), .B1(new_n730), .B2(new_n394), .ZN(new_n768));
  INV_X1    g582(.A(new_n450), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT110), .B1(new_n762), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n766), .B1(new_n445), .B2(new_n450), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n772), .A2(new_n761), .A3(new_n773), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(KEYINPUT111), .A2(KEYINPUT42), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n775), .A2(new_n389), .A3(new_n721), .A4(new_n777), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n389), .B(new_n721), .C1(new_n771), .C2(new_n774), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n776), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G131), .ZN(G33));
  OAI211_X1 g596(.A(new_n389), .B(new_n686), .C1(new_n771), .C2(new_n774), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  NAND2_X1  g598(.A1(new_n626), .A2(new_n645), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT43), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n681), .A2(new_n636), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT112), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n394), .B1(new_n457), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(new_n793), .B2(new_n457), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n765), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(KEYINPUT46), .A3(new_n765), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n451), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n521), .A2(new_n758), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n800), .A2(new_n719), .A3(new_n707), .A4(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n790), .B2(new_n789), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n792), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G137), .ZN(G39));
  NAND2_X1  g620(.A1(new_n800), .A2(new_n719), .ZN(new_n807));
  XOR2_X1   g621(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(KEYINPUT113), .A2(KEYINPUT47), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n810), .B1(new_n800), .B2(new_n719), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n716), .A2(new_n634), .A3(new_n720), .A4(new_n801), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G140), .ZN(G42));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n816));
  INV_X1    g630(.A(new_n750), .ZN(new_n817));
  INV_X1    g631(.A(new_n617), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n787), .A2(new_n818), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n819), .A2(KEYINPUT117), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(KEYINPUT117), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n817), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n702), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n822), .A2(new_n462), .A3(new_n823), .A4(new_n732), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT50), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n451), .B1(new_n394), .B2(new_n730), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n719), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n822), .B(new_n802), .C1(new_n812), .C2(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n699), .B1(new_n714), .B2(new_n715), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n388), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n826), .A2(new_n761), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n830), .A2(new_n831), .A3(new_n818), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n832), .A2(new_n573), .A3(new_n625), .A4(new_n645), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n831), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n820), .B2(new_n821), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n749), .A2(new_n681), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n836), .A2(KEYINPUT118), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT118), .B1(new_n836), .B2(new_n837), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n828), .B(new_n834), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n816), .B1(new_n825), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT50), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n824), .B(new_n842), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n838), .A2(new_n839), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n828), .A2(new_n834), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .A4(KEYINPUT51), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n822), .A2(new_n743), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT119), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT48), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n836), .A2(new_n849), .A3(new_n389), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n849), .B1(new_n836), .B2(new_n389), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g666(.A(G952), .B(new_n364), .C1(new_n832), .C2(new_n646), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n848), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n841), .A2(new_n846), .A3(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n663), .A2(new_n613), .A3(new_n615), .A4(new_n685), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n801), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n682), .A2(new_n857), .A3(new_n460), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n748), .A2(new_n721), .A3(new_n675), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n859), .B1(new_n771), .B2(new_n774), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n783), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n778), .B2(new_n780), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT114), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n629), .A2(new_n460), .A3(new_n523), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n716), .A2(new_n634), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n626), .A2(new_n664), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n646), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n523), .A3(new_n621), .ZN(new_n868));
  OAI22_X1  g682(.A1(new_n864), .A2(new_n865), .B1(new_n637), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n864), .A2(new_n676), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n863), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n636), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n388), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n639), .B1(new_n866), .B2(new_n646), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n873), .A2(new_n460), .A3(new_n523), .A4(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(new_n630), .A3(new_n678), .A4(KEYINPUT114), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n744), .A2(new_n736), .A3(new_n733), .A4(new_n752), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n862), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n685), .A2(KEYINPUT115), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n685), .A2(KEYINPUT115), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n881), .A2(new_n882), .A3(new_n393), .ZN(new_n883));
  AND4_X1   g697(.A1(new_n384), .A2(new_n385), .A3(new_n674), .A4(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n829), .A2(new_n884), .A3(new_n751), .A4(new_n770), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n460), .A2(new_n686), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n885), .B1(new_n717), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n755), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT52), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n888), .A2(new_n889), .A3(new_n727), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n889), .B1(new_n888), .B2(new_n727), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT116), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n723), .A2(new_n726), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT106), .B1(new_n732), .B2(new_n683), .ZN(new_n894));
  AND4_X1   g708(.A1(KEYINPUT106), .A2(new_n683), .A3(new_n738), .A4(new_n451), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n859), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n687), .A3(new_n885), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT52), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT116), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n888), .A2(new_n889), .A3(new_n727), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n880), .A2(new_n892), .A3(KEYINPUT53), .A4(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n878), .B1(new_n871), .B2(new_n876), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(new_n862), .A3(new_n900), .A4(new_n898), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT54), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n880), .A2(KEYINPUT53), .A3(new_n900), .A4(new_n898), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n890), .A2(new_n891), .A3(KEYINPUT116), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n899), .B1(new_n898), .B2(new_n900), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n862), .A2(new_n877), .A3(new_n879), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n909), .B(new_n910), .C1(new_n914), .C2(KEYINPUT53), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n908), .A2(new_n915), .ZN(new_n916));
  OAI22_X1  g730(.A1(new_n855), .A2(new_n916), .B1(G952), .B2(G953), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n826), .B(KEYINPUT49), .Z(new_n918));
  NOR3_X1   g732(.A1(new_n785), .A2(new_n393), .A3(new_n462), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n830), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n917), .B1(new_n702), .B2(new_n920), .ZN(G75));
  NAND3_X1  g735(.A1(new_n880), .A2(new_n892), .A3(new_n901), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n905), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n910), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT122), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n924), .A2(new_n925), .A3(G210), .A4(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n490), .B(KEYINPUT121), .Z(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT55), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n654), .B(KEYINPUT120), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT56), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n303), .B1(new_n923), .B2(new_n910), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n925), .B1(new_n934), .B2(G210), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n364), .A2(G952), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT123), .Z(new_n938));
  AOI21_X1  g752(.A(KEYINPUT56), .B1(new_n934), .B2(G210), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n938), .B1(new_n939), .B2(new_n930), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n936), .A2(new_n940), .ZN(G51));
  INV_X1    g755(.A(new_n938), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n764), .B(KEYINPUT57), .ZN(new_n943));
  INV_X1    g757(.A(new_n915), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n909), .B1(new_n923), .B2(new_n910), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n448), .ZN(new_n947));
  INV_X1    g761(.A(new_n934), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n948), .A2(new_n795), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n942), .B1(new_n947), .B2(new_n949), .ZN(G54));
  NAND3_X1  g764(.A1(new_n934), .A2(KEYINPUT58), .A3(G475), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n559), .A3(new_n562), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n559), .A2(new_n562), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n934), .A2(KEYINPUT58), .A3(G475), .A4(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n942), .B1(new_n952), .B2(new_n954), .ZN(G60));
  NAND2_X1  g769(.A1(G478), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT59), .Z(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n908), .B2(new_n915), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n641), .A2(new_n642), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n938), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n959), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n961), .A2(new_n957), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n944), .B2(new_n945), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT124), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT124), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n965), .B(new_n962), .C1(new_n944), .C2(new_n945), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n960), .B1(new_n964), .B2(new_n966), .ZN(G63));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT60), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n923), .B2(new_n910), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n673), .ZN(new_n971));
  AOI21_X1  g785(.A(KEYINPUT61), .B1(new_n971), .B2(KEYINPUT125), .ZN(new_n972));
  INV_X1    g786(.A(new_n376), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n904), .A2(new_n905), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n905), .B2(new_n922), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n973), .B1(new_n975), .B2(new_n969), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(new_n971), .A3(new_n938), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n972), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n942), .B1(new_n970), .B2(new_n673), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT125), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(new_n970), .B2(new_n673), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n976), .B(new_n979), .C1(new_n981), .C2(KEYINPUT61), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n978), .A2(new_n982), .ZN(G66));
  NAND2_X1  g797(.A1(new_n618), .A2(new_n488), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(G953), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n903), .B2(G953), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n929), .B1(G898), .B2(new_n364), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(G69));
  XNOR2_X1  g802(.A(new_n262), .B(new_n549), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n389), .A2(new_n802), .A3(new_n867), .ZN(new_n990));
  AOI22_X1  g804(.A1(new_n812), .A2(new_n813), .B1(new_n708), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n805), .A2(new_n991), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n727), .A2(new_n687), .A3(new_n896), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n710), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT62), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n710), .A2(KEYINPUT62), .A3(new_n993), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n992), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n989), .B1(new_n998), .B2(G953), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n364), .B1(G227), .B2(G900), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n989), .B1(G900), .B2(G953), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n389), .A2(new_n751), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n1003), .A2(new_n719), .A3(new_n707), .A4(new_n800), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n814), .A2(new_n783), .A3(new_n1004), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n1005), .A2(new_n781), .A3(new_n805), .A4(new_n993), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1002), .B1(new_n1006), .B2(G953), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n999), .A2(new_n1001), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT126), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT127), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n999), .A2(new_n1007), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1012), .B1(new_n1013), .B2(new_n1000), .ZN(new_n1014));
  AOI211_X1 g828(.A(KEYINPUT127), .B(new_n1001), .C1(new_n999), .C2(new_n1007), .ZN(new_n1015));
  OAI22_X1  g829(.A1(new_n1010), .A2(new_n1011), .B1(new_n1014), .B2(new_n1015), .ZN(G72));
  NAND2_X1  g830(.A1(new_n998), .A2(new_n903), .ZN(new_n1017));
  NAND2_X1  g831(.A1(G472), .A2(G902), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT63), .Z(new_n1019));
  AOI211_X1 g833(.A(new_n266), .B(new_n263), .C1(new_n1017), .C2(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(new_n903), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1019), .B1(new_n1006), .B2(new_n1021), .ZN(new_n1022));
  AND3_X1   g836(.A1(new_n1022), .A2(new_n266), .A3(new_n263), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n281), .A2(new_n282), .A3(new_n289), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n907), .A2(new_n1019), .A3(new_n1024), .ZN(new_n1025));
  NOR4_X1   g839(.A1(new_n1020), .A2(new_n1023), .A3(new_n942), .A4(new_n1025), .ZN(G57));
endmodule


