//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT5), .ZN(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G148gat), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G141gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n209), .A2(new_n211), .B1(KEYINPUT2), .B2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT80), .B1(G155gat), .B2(G162gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT80), .ZN(new_n215));
  INV_X1    g014(.A(G155gat), .ZN(new_n216));
  INV_X1    g015(.A(G162gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT79), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n219), .B1(G155gat), .B2(G162gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n212), .A2(KEYINPUT79), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n214), .B(new_n218), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT81), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n213), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n218), .A2(new_n214), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n225), .B(KEYINPUT81), .C1(new_n220), .C2(new_n221), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(G141gat), .A3(new_n229), .ZN(new_n230));
  OR3_X1    g029(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n230), .A2(new_n209), .B1(new_n231), .B2(new_n212), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G113gat), .B(G120gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(KEYINPUT1), .ZN(new_n236));
  XNOR2_X1  g035(.A(G127gat), .B(G134gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n237), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(KEYINPUT1), .B2(new_n235), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n234), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n233), .A3(new_n241), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G225gat), .A2(G233gat), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n207), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT4), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n232), .B1(new_n224), .B2(new_n226), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(KEYINPUT4), .A3(new_n241), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n234), .A2(KEYINPUT83), .A3(KEYINPUT3), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT83), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n255), .B1(new_n251), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n227), .A2(new_n256), .A3(new_n233), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n242), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n253), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n248), .B1(new_n262), .B2(new_n246), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n260), .B1(new_n257), .B2(new_n254), .ZN(new_n264));
  NOR4_X1   g063(.A1(new_n264), .A2(new_n253), .A3(new_n207), .A4(new_n247), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n206), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT6), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n258), .A2(new_n261), .ZN(new_n268));
  INV_X1    g067(.A(new_n253), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT5), .A4(new_n246), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n205), .B(KEYINPUT87), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n264), .A2(new_n247), .A3(new_n253), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n270), .B(new_n272), .C1(new_n273), .C2(new_n248), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n266), .A2(new_n267), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n248), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n268), .A2(new_n269), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n276), .B1(new_n277), .B2(new_n247), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n278), .A2(KEYINPUT6), .A3(new_n205), .A4(new_n270), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G211gat), .B(G218gat), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G218gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT73), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G218gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT22), .B1(new_n287), .B2(G211gat), .ZN(new_n288));
  XOR2_X1   g087(.A(G197gat), .B(G204gat), .Z(new_n289));
  OAI21_X1  g088(.A(new_n282), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT22), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT73), .B(G218gat), .ZN(new_n292));
  INV_X1    g091(.A(G211gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n289), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(new_n295), .A3(new_n281), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G226gat), .A2(G233gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT74), .ZN(new_n299));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n301), .B1(new_n303), .B2(KEYINPUT26), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT68), .B(KEYINPUT26), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n305), .B1(new_n306), .B2(new_n302), .ZN(new_n307));
  AND2_X1   g106(.A1(KEYINPUT68), .A2(KEYINPUT26), .ZN(new_n308));
  NOR2_X1   g107(.A1(KEYINPUT68), .A2(KEYINPUT26), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n305), .B(new_n302), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n304), .B1(new_n307), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G183gat), .A2(G190gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G183gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT27), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT27), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G183gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT66), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT66), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n316), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT28), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(G190gat), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n320), .A2(KEYINPUT67), .A3(new_n322), .A4(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n323), .B1(new_n319), .B2(G190gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT67), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n314), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT65), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NOR3_X1   g133(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n300), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n337));
  AND2_X1   g136(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n313), .A2(new_n337), .B1(new_n338), .B2(G190gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n332), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n313), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(G190gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT23), .ZN(new_n344));
  INV_X1    g143(.A(G169gat), .ZN(new_n345));
  INV_X1    g144(.A(G176gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n301), .B1(new_n347), .B2(new_n333), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT64), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n340), .B(KEYINPUT25), .C1(new_n349), .C2(new_n332), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n336), .A2(new_n339), .ZN(new_n352));
  OAI211_X1 g151(.A(KEYINPUT65), .B(new_n351), .C1(new_n352), .C2(KEYINPUT64), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n299), .B1(new_n331), .B2(new_n354), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n350), .A2(new_n353), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n328), .A2(new_n329), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(new_n325), .A3(new_n326), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n302), .B1(new_n308), .B2(new_n309), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT69), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n310), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n361), .A2(new_n304), .B1(G183gat), .B2(G190gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n356), .A2(KEYINPUT74), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n298), .B1(new_n355), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n298), .ZN(new_n366));
  AOI211_X1 g165(.A(KEYINPUT29), .B(new_n366), .C1(new_n356), .C2(new_n363), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n297), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  XOR2_X1   g167(.A(KEYINPUT75), .B(KEYINPUT29), .Z(new_n369));
  NAND4_X1  g168(.A1(new_n355), .A2(new_n364), .A3(new_n369), .A4(new_n298), .ZN(new_n370));
  INV_X1    g169(.A(new_n297), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n363), .A3(new_n366), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  XOR2_X1   g173(.A(G8gat), .B(G36gat), .Z(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(KEYINPUT76), .ZN(new_n376));
  XNOR2_X1  g175(.A(G64gat), .B(G92gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n376), .B(new_n377), .Z(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT77), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n378), .B1(new_n368), .B2(new_n373), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n368), .A2(new_n373), .A3(KEYINPUT30), .A4(new_n378), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n373), .A3(new_n378), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT30), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n381), .A2(new_n384), .A3(new_n385), .A4(new_n388), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n280), .A2(new_n389), .A3(KEYINPUT35), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT86), .ZN(new_n391));
  XNOR2_X1  g190(.A(G78gat), .B(G106gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(KEYINPUT31), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(G50gat), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT29), .B1(new_n290), .B2(new_n296), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT84), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n256), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI211_X1 g196(.A(KEYINPUT84), .B(KEYINPUT29), .C1(new_n290), .C2(new_n296), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n234), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT85), .ZN(new_n400));
  INV_X1    g199(.A(new_n369), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(new_n251), .B2(new_n256), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n400), .B1(new_n402), .B2(new_n297), .ZN(new_n403));
  INV_X1    g202(.A(G228gat), .ZN(new_n404));
  INV_X1    g203(.A(G233gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI211_X1 g205(.A(KEYINPUT3), .B(new_n232), .C1(new_n224), .C2(new_n226), .ZN(new_n407));
  OAI211_X1 g206(.A(KEYINPUT85), .B(new_n371), .C1(new_n407), .C2(new_n401), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n399), .A2(new_n403), .A3(new_n406), .A4(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(G22gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n402), .A2(new_n297), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n297), .A2(new_n369), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n251), .B1(new_n412), .B2(new_n256), .ZN(new_n413));
  OAI22_X1  g212(.A1(new_n411), .A2(new_n413), .B1(new_n404), .B2(new_n405), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n409), .A2(new_n410), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n410), .B1(new_n409), .B2(new_n414), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n391), .B(new_n394), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n409), .A2(new_n414), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G22gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n409), .A2(new_n410), .A3(new_n414), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n394), .B1(new_n422), .B2(new_n391), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(KEYINPUT86), .A3(new_n421), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n418), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n241), .A2(KEYINPUT70), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT70), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n242), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n426), .B(new_n428), .C1(new_n331), .C2(new_n354), .ZN(new_n429));
  INV_X1    g228(.A(G227gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n430), .A2(new_n405), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n356), .A2(new_n427), .A3(new_n363), .A4(new_n242), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT71), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n429), .A2(new_n432), .A3(KEYINPUT71), .A4(new_n431), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT33), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n429), .A2(new_n432), .ZN(new_n440));
  INV_X1    g239(.A(new_n431), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT34), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT34), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n440), .A2(new_n444), .A3(new_n441), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  XOR2_X1   g245(.A(G15gat), .B(G43gat), .Z(new_n447));
  XNOR2_X1  g246(.A(G71gat), .B(G99gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n439), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n437), .A2(KEYINPUT32), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n444), .B1(new_n440), .B2(new_n441), .ZN(new_n453));
  AOI211_X1 g252(.A(KEYINPUT34), .B(new_n431), .C1(new_n429), .C2(new_n432), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT33), .B1(new_n435), .B2(new_n436), .ZN(new_n456));
  INV_X1    g255(.A(new_n449), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n450), .A2(new_n452), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n452), .B1(new_n450), .B2(new_n458), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n390), .A2(new_n425), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT78), .ZN(new_n463));
  INV_X1    g262(.A(new_n384), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n385), .B1(new_n382), .B2(new_n383), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n278), .A2(new_n205), .A3(new_n270), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(new_n266), .A3(new_n267), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n468), .A2(new_n279), .B1(new_n387), .B2(new_n386), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n381), .A2(KEYINPUT78), .A3(new_n384), .A4(new_n385), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n466), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n446), .B1(new_n439), .B2(new_n449), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n451), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n450), .A2(new_n452), .A3(new_n458), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n425), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT92), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n461), .A2(KEYINPUT92), .A3(new_n425), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n471), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT35), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n462), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n275), .A2(new_n279), .A3(new_n386), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT90), .B1(new_n374), .B2(KEYINPUT37), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n374), .A2(KEYINPUT37), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT90), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT37), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n368), .A2(new_n373), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n484), .A2(new_n485), .A3(new_n379), .A4(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n483), .B1(KEYINPUT38), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n484), .A2(new_n379), .A3(new_n488), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n371), .B1(new_n365), .B2(new_n367), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n370), .A2(new_n297), .A3(new_n372), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(KEYINPUT37), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT89), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT38), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n493), .A2(new_n494), .A3(new_n498), .A4(KEYINPUT37), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n492), .A2(new_n501), .A3(KEYINPUT91), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT91), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(new_n491), .B2(new_n500), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n490), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n423), .A2(new_n424), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n417), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT39), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n508), .B(new_n247), .C1(new_n264), .C2(new_n253), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n262), .A2(new_n246), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT39), .B1(new_n245), .B2(new_n247), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n271), .B(new_n509), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT40), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n274), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n277), .A2(new_n247), .ZN(new_n515));
  INV_X1    g314(.A(new_n511), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n272), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT40), .B1(new_n517), .B2(new_n509), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n389), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT88), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n507), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n389), .A2(new_n519), .A3(KEYINPUT88), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n525), .A2(KEYINPUT72), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(KEYINPUT72), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n474), .B(new_n475), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  OAI22_X1  g327(.A1(new_n459), .A2(new_n460), .B1(KEYINPUT72), .B2(new_n525), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n528), .A2(new_n529), .B1(new_n471), .B2(new_n507), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n482), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n533), .A2(KEYINPUT98), .ZN(new_n534));
  XOR2_X1   g333(.A(G57gat), .B(G64gat), .Z(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(KEYINPUT98), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G71gat), .B(G78gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n534), .A2(new_n535), .A3(new_n538), .A4(new_n536), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT21), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G231gat), .A2(G233gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G127gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(G183gat), .B(G211gat), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n546), .B(G127gat), .ZN(new_n551));
  INV_X1    g350(.A(new_n549), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G1gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT16), .ZN(new_n556));
  INV_X1    g355(.A(G15gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n410), .ZN(new_n558));
  NAND2_X1  g357(.A1(G15gat), .A2(G22gat), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n556), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT94), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(G8gat), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n562), .A2(G8gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n558), .A2(G1gat), .A3(new_n559), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n561), .A2(new_n563), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n565), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n562), .B(G8gat), .C1(new_n567), .C2(new_n560), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(new_n542), .B2(new_n543), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT99), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(new_n216), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n571), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n554), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(G29gat), .ZN(new_n576));
  INV_X1    g375(.A(G36gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n577), .A3(KEYINPUT14), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT14), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n579), .B1(G29gat), .B2(G36gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(G43gat), .ZN(new_n583));
  INV_X1    g382(.A(G50gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G43gat), .A2(G50gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT15), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT93), .B(G29gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(G36gat), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT15), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n585), .A2(new_n591), .A3(new_n586), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n582), .A2(new_n588), .A3(new_n590), .A4(new_n592), .ZN(new_n593));
  OR2_X1    g392(.A1(KEYINPUT93), .A2(G29gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(KEYINPUT93), .A2(G29gat), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n577), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g395(.A(KEYINPUT15), .B(new_n587), .C1(new_n596), .C2(new_n581), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT17), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n593), .A2(new_n597), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT17), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G99gat), .A2(G106gat), .ZN(new_n603));
  INV_X1    g402(.A(G85gat), .ZN(new_n604));
  INV_X1    g403(.A(G92gat), .ZN(new_n605));
  AOI22_X1  g404(.A1(KEYINPUT8), .A2(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT103), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT7), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n607), .B(new_n608), .C1(new_n604), .C2(new_n605), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  OAI211_X1 g409(.A(G85gat), .B(G92gat), .C1(KEYINPUT103), .C2(KEYINPUT7), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n606), .B(new_n609), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G99gat), .B(G106gat), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n610), .A2(new_n611), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n616), .A2(new_n613), .A3(new_n609), .A4(new_n606), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n599), .A2(new_n602), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT100), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT41), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n618), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n623), .B1(new_n624), .B2(new_n600), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n619), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(G190gat), .ZN(new_n627));
  INV_X1    g426(.A(G190gat), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n619), .A2(new_n628), .A3(new_n625), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(G218gat), .A3(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n630), .A2(KEYINPUT102), .ZN(new_n631));
  INV_X1    g430(.A(new_n629), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n628), .B1(new_n619), .B2(new_n625), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n283), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n631), .A2(new_n217), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n634), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n630), .A2(KEYINPUT102), .ZN(new_n637));
  OAI21_X1  g436(.A(G162gat), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n622), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(KEYINPUT101), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G134gat), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n635), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n217), .B1(new_n631), .B2(new_n634), .ZN(new_n644));
  AND4_X1   g443(.A1(KEYINPUT102), .A2(new_n634), .A3(new_n630), .A4(new_n217), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n575), .B1(new_n642), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G113gat), .B(G141gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G197gat), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT11), .B(G169gat), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT12), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT95), .B1(new_n598), .B2(new_n569), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT95), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n600), .A2(new_n656), .A3(new_n568), .A4(new_n566), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n598), .A2(new_n569), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G229gat), .A2(G233gat), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n661), .B(KEYINPUT13), .Z(new_n662));
  NAND3_X1  g461(.A1(new_n660), .A2(KEYINPUT96), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT96), .ZN(new_n664));
  AOI22_X1  g463(.A1(new_n655), .A2(new_n657), .B1(new_n569), .B2(new_n598), .ZN(new_n665));
  INV_X1    g464(.A(new_n662), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n599), .A2(new_n569), .A3(new_n602), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n658), .A2(new_n661), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT18), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n658), .A2(new_n669), .A3(KEYINPUT18), .A4(new_n661), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n654), .B1(new_n668), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n663), .A2(new_n667), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n676), .A2(new_n653), .A3(new_n672), .A4(new_n673), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n675), .A2(KEYINPUT97), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT97), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n679), .B(new_n654), .C1(new_n668), .C2(new_n674), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(G230gat), .A2(G233gat), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n540), .A2(new_n615), .A3(new_n541), .A4(new_n617), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT10), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n542), .A2(new_n618), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT104), .B(KEYINPUT10), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n686), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n687), .A2(KEYINPUT105), .A3(new_n684), .A4(new_n688), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n683), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n687), .A2(new_n684), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n683), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(G120gat), .B(G148gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(G176gat), .B(G204gat), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n696), .B(new_n697), .Z(new_n698));
  OR2_X1    g497(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n689), .A2(new_n690), .ZN(new_n700));
  INV_X1    g499(.A(new_n686), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(new_n692), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n682), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n694), .A2(new_n683), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n704), .A3(new_n698), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n648), .A2(new_n681), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n532), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n468), .A2(new_n279), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(new_n555), .ZN(G1324gat));
  INV_X1    g510(.A(new_n708), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n389), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT42), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT16), .B(G8gat), .ZN(new_n715));
  OR3_X1    g514(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(G8gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n714), .B1(new_n713), .B2(new_n715), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT106), .ZN(G1325gat));
  NAND2_X1  g519(.A1(new_n528), .A2(new_n529), .ZN(new_n721));
  OAI21_X1  g520(.A(G15gat), .B1(new_n708), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n461), .A2(new_n557), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n708), .B2(new_n723), .ZN(G1326gat));
  NAND2_X1  g523(.A1(new_n712), .A2(new_n507), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT107), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT43), .B(G22gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1327gat));
  NOR3_X1   g527(.A1(new_n644), .A2(new_n643), .A3(new_n645), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n641), .B1(new_n635), .B2(new_n638), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n462), .ZN(new_n732));
  INV_X1    g531(.A(new_n471), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT92), .B1(new_n461), .B2(new_n425), .ZN(new_n734));
  AND4_X1   g533(.A1(KEYINPUT92), .A2(new_n425), .A3(new_n475), .A4(new_n474), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n732), .B1(new_n736), .B2(KEYINPUT35), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n524), .A2(new_n530), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n731), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n575), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n741), .A2(new_n681), .A3(new_n706), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n743), .A2(new_n709), .A3(new_n589), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n744), .B(KEYINPUT45), .Z(new_n745));
  AOI21_X1  g544(.A(KEYINPUT44), .B1(new_n532), .B2(new_n731), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n646), .A2(new_n642), .ZN(new_n748));
  AOI211_X1 g547(.A(new_n747), .B(new_n748), .C1(new_n482), .C2(new_n531), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n742), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n589), .B1(new_n751), .B2(new_n709), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n745), .A2(new_n752), .ZN(G1328gat));
  INV_X1    g552(.A(new_n389), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n577), .B1(new_n755), .B2(KEYINPUT108), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n743), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(KEYINPUT108), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G36gat), .B1(new_n751), .B2(new_n754), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(G1329gat));
  INV_X1    g560(.A(new_n461), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n583), .B1(new_n743), .B2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n721), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G43gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n751), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g566(.A(G50gat), .B1(new_n751), .B2(new_n425), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n740), .A2(new_n584), .A3(new_n507), .A4(new_n742), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT48), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n770), .B(new_n772), .ZN(G1331gat));
  NAND3_X1  g572(.A1(new_n647), .A2(new_n681), .A3(new_n706), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT110), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n482), .B2(new_n531), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n709), .B(KEYINPUT111), .Z(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g578(.A(new_n754), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT112), .ZN(new_n782));
  NOR2_X1   g581(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1333gat));
  NAND2_X1  g583(.A1(new_n776), .A2(new_n764), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n762), .A2(G71gat), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n785), .A2(G71gat), .B1(new_n776), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g587(.A1(new_n776), .A2(new_n507), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g589(.A1(new_n678), .A2(new_n680), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n741), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n731), .B(new_n792), .C1(new_n737), .C2(new_n738), .ZN(new_n793));
  AND2_X1   g592(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n532), .A2(new_n731), .A3(new_n792), .A4(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n795), .A2(new_n706), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n604), .B1(new_n799), .B2(new_n709), .ZN(new_n800));
  INV_X1    g599(.A(new_n709), .ZN(new_n801));
  INV_X1    g600(.A(new_n706), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n741), .A2(new_n791), .A3(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n750), .A2(G85gat), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT114), .ZN(G1336gat));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n750), .A2(new_n389), .A3(new_n803), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G92gat), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n807), .B1(new_n809), .B2(KEYINPUT115), .ZN(new_n810));
  OR3_X1    g609(.A1(new_n799), .A2(G92gat), .A3(new_n754), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n809), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n811), .B(new_n809), .C1(KEYINPUT115), .C2(new_n807), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(G1337gat));
  NAND3_X1  g614(.A1(new_n750), .A2(new_n764), .A3(new_n803), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT116), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(G99gat), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n816), .A2(KEYINPUT116), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n762), .A2(G99gat), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n818), .A2(new_n819), .B1(new_n799), .B2(new_n820), .ZN(G1338gat));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n425), .A2(G106gat), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n795), .A2(new_n706), .A3(new_n798), .A4(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n750), .A2(KEYINPUT118), .A3(new_n507), .A4(new_n803), .ZN(new_n827));
  INV_X1    g626(.A(G106gat), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n739), .A2(new_n747), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n532), .A2(KEYINPUT44), .A3(new_n731), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n829), .A2(new_n507), .A3(new_n830), .A4(new_n803), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI211_X1 g632(.A(new_n822), .B(new_n826), .C1(new_n827), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n831), .A2(new_n832), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n827), .A2(new_n835), .A3(G106gat), .ZN(new_n836));
  INV_X1    g635(.A(new_n826), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT119), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n831), .A2(G106gat), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n824), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT117), .B1(new_n840), .B2(KEYINPUT53), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n842));
  AOI211_X1 g641(.A(new_n842), .B(new_n825), .C1(new_n839), .C2(new_n824), .ZN(new_n843));
  OAI22_X1  g642(.A1(new_n834), .A2(new_n838), .B1(new_n841), .B2(new_n843), .ZN(G1339gat));
  NAND3_X1  g643(.A1(new_n691), .A2(new_n683), .A3(new_n692), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n703), .A2(KEYINPUT54), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n698), .B1(new_n693), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n848), .A3(KEYINPUT55), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n705), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT121), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n846), .A2(new_n848), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n849), .A2(new_n855), .A3(new_n705), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n851), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n660), .A2(new_n662), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n661), .B1(new_n658), .B2(new_n669), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n652), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n677), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n857), .A2(new_n731), .A3(new_n861), .ZN(new_n862));
  AOI22_X1  g661(.A1(new_n857), .A2(new_n791), .B1(new_n706), .B2(new_n861), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(new_n731), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n741), .A2(new_n748), .A3(new_n681), .A4(new_n802), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT120), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n647), .A2(new_n867), .A3(new_n681), .A4(new_n802), .ZN(new_n868));
  AOI22_X1  g667(.A1(new_n864), .A2(new_n575), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n870), .A2(new_n777), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n734), .A2(new_n735), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n871), .A2(new_n873), .A3(new_n754), .ZN(new_n874));
  AOI21_X1  g673(.A(G113gat), .B1(new_n874), .B2(new_n791), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n869), .A2(new_n507), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n389), .A2(new_n709), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n876), .A2(new_n461), .A3(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n791), .A2(G113gat), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n875), .B1(new_n878), .B2(new_n879), .ZN(G1340gat));
  AOI21_X1  g679(.A(G120gat), .B1(new_n874), .B2(new_n706), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n706), .A2(G120gat), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n878), .B2(new_n882), .ZN(G1341gat));
  NAND3_X1  g682(.A1(new_n874), .A2(new_n547), .A3(new_n741), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n878), .A2(new_n741), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n547), .ZN(G1342gat));
  AND2_X1   g685(.A1(new_n878), .A2(new_n731), .ZN(new_n887));
  INV_X1    g686(.A(G134gat), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n888), .A3(new_n731), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(KEYINPUT56), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n891), .B1(KEYINPUT56), .B2(new_n890), .ZN(G1343gat));
  NAND2_X1  g691(.A1(new_n721), .A2(new_n877), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n849), .A2(new_n705), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n894), .A2(new_n678), .A3(new_n680), .A4(new_n854), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n706), .A2(new_n861), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n731), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n856), .A2(new_n854), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n851), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n646), .A2(new_n642), .A3(new_n861), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n575), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n866), .A2(new_n868), .ZN(new_n905));
  OAI211_X1 g704(.A(KEYINPUT122), .B(new_n575), .C1(new_n897), .C2(new_n901), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n507), .A2(KEYINPUT57), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n911), .B1(new_n869), .B2(new_n425), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n893), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(G141gat), .A3(new_n791), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n764), .A2(new_n425), .A3(new_n389), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n871), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n208), .B1(new_n916), .B2(new_n681), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  XOR2_X1   g717(.A(new_n918), .B(KEYINPUT58), .Z(G1344gat));
  NAND2_X1  g718(.A1(new_n228), .A2(new_n229), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n922), .B1(new_n913), .B2(new_n706), .ZN(new_n923));
  INV_X1    g722(.A(new_n893), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n791), .A2(new_n898), .A3(new_n851), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n731), .B1(new_n925), .B2(new_n896), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n575), .B1(new_n926), .B2(new_n901), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n908), .B1(new_n927), .B2(new_n905), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n425), .B1(new_n902), .B2(new_n865), .ZN(new_n930));
  OAI22_X1  g729(.A1(new_n928), .A2(new_n929), .B1(new_n930), .B2(KEYINPUT57), .ZN(new_n931));
  AOI211_X1 g730(.A(KEYINPUT123), .B(new_n908), .C1(new_n927), .C2(new_n905), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n706), .B(new_n924), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT124), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT123), .B1(new_n869), .B2(new_n908), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n902), .A2(new_n865), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n911), .B1(new_n936), .B2(new_n425), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n928), .A2(new_n929), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n939), .A2(new_n940), .A3(new_n706), .A4(new_n924), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n934), .A2(new_n941), .A3(G148gat), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n923), .B1(new_n942), .B2(KEYINPUT59), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n916), .A2(new_n920), .A3(new_n802), .ZN(new_n944));
  OAI21_X1  g743(.A(KEYINPUT125), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n946));
  INV_X1    g745(.A(new_n944), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n210), .B1(new_n933), .B2(KEYINPUT124), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n921), .B1(new_n948), .B2(new_n941), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n946), .B(new_n947), .C1(new_n949), .C2(new_n923), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n945), .A2(new_n950), .ZN(G1345gat));
  INV_X1    g750(.A(new_n916), .ZN(new_n952));
  AOI21_X1  g751(.A(G155gat), .B1(new_n952), .B2(new_n741), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n741), .A2(G155gat), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT126), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n953), .B1(new_n913), .B2(new_n955), .ZN(G1346gat));
  NOR3_X1   g755(.A1(new_n916), .A2(G162gat), .A3(new_n748), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n217), .B1(new_n913), .B2(new_n731), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n957), .A2(new_n958), .ZN(G1347gat));
  NOR2_X1   g758(.A1(new_n777), .A2(new_n754), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n876), .A2(new_n461), .A3(new_n960), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n961), .A2(new_n345), .A3(new_n681), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n869), .A2(new_n801), .A3(new_n754), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n963), .A2(new_n873), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(new_n791), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n962), .B1(new_n345), .B2(new_n965), .ZN(G1348gat));
  NAND3_X1  g765(.A1(new_n964), .A2(new_n346), .A3(new_n706), .ZN(new_n967));
  OAI21_X1  g766(.A(G176gat), .B1(new_n961), .B2(new_n802), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(G1349gat));
  NAND4_X1  g768(.A1(new_n964), .A2(new_n320), .A3(new_n322), .A4(new_n741), .ZN(new_n970));
  OAI21_X1  g769(.A(G183gat), .B1(new_n961), .B2(new_n575), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g772(.A(G190gat), .B1(new_n961), .B2(new_n748), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT61), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n964), .A2(new_n628), .A3(new_n731), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1351gat));
  AND3_X1   g776(.A1(new_n963), .A2(new_n507), .A3(new_n721), .ZN(new_n978));
  AOI21_X1  g777(.A(G197gat), .B1(new_n978), .B2(new_n791), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n764), .A2(new_n754), .A3(new_n777), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n939), .A2(new_n980), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n791), .A2(G197gat), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(G1352gat));
  INV_X1    g782(.A(G204gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n978), .A2(new_n984), .A3(new_n706), .ZN(new_n985));
  XOR2_X1   g784(.A(new_n985), .B(KEYINPUT62), .Z(new_n986));
  AND3_X1   g785(.A1(new_n939), .A2(new_n706), .A3(new_n980), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n986), .B1(new_n984), .B2(new_n987), .ZN(G1353gat));
  NAND3_X1  g787(.A1(new_n939), .A2(new_n741), .A3(new_n980), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n990));
  OAI211_X1 g789(.A(new_n989), .B(G211gat), .C1(new_n990), .C2(KEYINPUT63), .ZN(new_n991));
  AND2_X1   g790(.A1(new_n990), .A2(KEYINPUT63), .ZN(new_n992));
  OR2_X1    g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n293), .A3(new_n741), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n991), .A2(new_n992), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(G1354gat));
  AOI21_X1  g795(.A(G218gat), .B1(new_n978), .B2(new_n731), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n748), .A2(new_n292), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n997), .B1(new_n981), .B2(new_n998), .ZN(G1355gat));
endmodule


