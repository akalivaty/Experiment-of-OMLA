//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n565, new_n566, new_n567, new_n568, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n600, new_n601,
    new_n602, new_n603, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n649, new_n650, new_n651,
    new_n652, new_n655, new_n657, new_n658, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1221, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(new_n462), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n465), .B1(new_n469), .B2(G137), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI211_X1 g048(.A(G137), .B(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(KEYINPUT69), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n464), .B1(new_n470), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n477), .B1(new_n472), .B2(new_n473), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n467), .A2(KEYINPUT68), .A3(new_n468), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n478), .A2(new_n479), .A3(G125), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n471), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n476), .A2(new_n482), .ZN(G160));
  NAND2_X1  g058(.A1(new_n469), .A2(G136), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n471), .B1(new_n467), .B2(new_n468), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n471), .A2(G112), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n484), .B(new_n486), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT70), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n492), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n478), .A2(new_n479), .A3(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n471), .A2(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT71), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n501), .A2(new_n503), .A3(new_n504), .A4(G2104), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n500), .A2(new_n505), .B1(new_n485), .B2(G126), .ZN(new_n506));
  AND3_X1   g081(.A1(new_n497), .A2(new_n506), .A3(KEYINPUT72), .ZN(new_n507));
  AOI21_X1  g082(.A(KEYINPUT72), .B1(new_n497), .B2(new_n506), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(G164));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT73), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT73), .A2(G651), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT6), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT74), .B1(new_n518), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT74), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT5), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n519), .A2(new_n522), .B1(new_n518), .B2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n510), .A2(new_n517), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  OR2_X1    g102(.A1(KEYINPUT73), .A2(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(KEYINPUT73), .A2(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n526), .A2(new_n532), .ZN(G166));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n523), .A2(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G89), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n524), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n541), .B1(new_n516), .B2(G543), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n516), .A2(new_n541), .A3(G543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n540), .B1(new_n545), .B2(G51), .ZN(G168));
  AOI21_X1  g121(.A(new_n514), .B1(new_n530), .B2(KEYINPUT6), .ZN(new_n547));
  NOR3_X1   g122(.A1(new_n547), .A2(KEYINPUT75), .A3(new_n521), .ZN(new_n548));
  OAI21_X1  g123(.A(G52), .B1(new_n548), .B2(new_n542), .ZN(new_n549));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n518), .A2(G543), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n520), .B1(KEYINPUT5), .B2(new_n521), .ZN(new_n552));
  NOR3_X1   g127(.A1(new_n518), .A2(KEYINPUT74), .A3(G543), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(G64), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n550), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n556), .A2(KEYINPUT76), .A3(new_n530), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n547), .A2(new_n554), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G90), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n561), .B2(new_n531), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n549), .A2(new_n557), .A3(new_n559), .A4(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(G171));
  AOI22_X1  g139(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G81), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n565), .A2(new_n531), .B1(new_n524), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n545), .B2(G43), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  AOI22_X1  g148(.A1(new_n523), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G651), .ZN(new_n575));
  INV_X1    g150(.A(G91), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n574), .A2(new_n575), .B1(new_n524), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  NAND2_X1  g154(.A1(G53), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n516), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n582), .A2(KEYINPUT77), .A3(KEYINPUT9), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n580), .B1(new_n513), .B2(new_n515), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n585), .B1(new_n586), .B2(new_n579), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT9), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n586), .B2(new_n585), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n583), .B(new_n584), .C1(new_n587), .C2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n582), .A2(KEYINPUT77), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT6), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n528), .B2(new_n529), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n585), .B(new_n581), .C1(new_n594), .C2(new_n514), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(KEYINPUT9), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n584), .B1(new_n597), .B2(new_n583), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n578), .B1(new_n591), .B2(new_n598), .ZN(G299));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n563), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n563), .A2(new_n600), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n602), .A2(new_n603), .ZN(G301));
  INV_X1    g179(.A(G168), .ZN(G286));
  INV_X1    g180(.A(G166), .ZN(G303));
  NAND3_X1  g181(.A1(new_n516), .A2(new_n523), .A3(G87), .ZN(new_n607));
  OAI21_X1  g182(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n516), .A2(G49), .A3(G543), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(G288));
  NAND3_X1  g185(.A1(new_n516), .A2(new_n523), .A3(G86), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n516), .A2(G48), .A3(G543), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g188(.A1(new_n523), .A2(G61), .ZN(new_n614));
  AND2_X1   g189(.A1(G73), .A2(G543), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n530), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n613), .A2(new_n616), .ZN(G305));
  AOI22_X1  g192(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(new_n531), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(G85), .B2(new_n558), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n545), .A2(G47), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(G290));
  INV_X1    g197(.A(G868), .ZN(new_n623));
  NOR2_X1   g198(.A1(G301), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n558), .A2(G92), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT10), .Z(new_n626));
  NAND2_X1  g201(.A1(G79), .A2(G543), .ZN(new_n627));
  INV_X1    g202(.A(G66), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n554), .B2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT81), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g206(.A(KEYINPUT81), .B(new_n627), .C1(new_n554), .C2(new_n628), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(G651), .A3(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n634));
  OAI21_X1  g209(.A(G54), .B1(new_n548), .B2(new_n542), .ZN(new_n635));
  AND3_X1   g210(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n634), .B1(new_n633), .B2(new_n635), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n626), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT83), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n633), .A2(new_n635), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT82), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n644), .A2(KEYINPUT83), .A3(new_n626), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n624), .B1(new_n646), .B2(new_n623), .ZN(G284));
  AOI21_X1  g222(.A(new_n624), .B1(new_n646), .B2(new_n623), .ZN(G321));
  NAND2_X1  g223(.A1(G286), .A2(G868), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n583), .B1(new_n587), .B2(new_n589), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(KEYINPUT79), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n577), .B1(new_n651), .B2(new_n590), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n649), .B1(new_n652), .B2(G868), .ZN(G297));
  OAI21_X1  g228(.A(new_n649), .B1(new_n652), .B2(G868), .ZN(G280));
  INV_X1    g229(.A(G559), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n646), .B1(new_n655), .B2(G860), .ZN(G148));
  NAND2_X1  g231(.A1(new_n646), .A2(new_n655), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G868), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(G868), .B2(new_n568), .ZN(G323));
  XNOR2_X1  g234(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g235(.A1(new_n478), .A2(new_n479), .A3(new_n463), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT12), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT13), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n663), .A2(G2100), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(G2100), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n469), .A2(G135), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n485), .A2(G123), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n471), .A2(G111), .ZN(new_n668));
  OAI21_X1  g243(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n666), .B(new_n667), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT84), .B(G2096), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n664), .A2(new_n665), .A3(new_n672), .ZN(G156));
  XNOR2_X1  g248(.A(G2427), .B(G2438), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2430), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT15), .B(G2435), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n677), .A2(KEYINPUT14), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT85), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2451), .B(G2454), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT16), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2443), .B(G2446), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n680), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1341), .B(G1348), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n687), .A2(new_n688), .A3(G14), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G401));
  XNOR2_X1  g265(.A(G2072), .B(G2078), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT17), .ZN(new_n692));
  XNOR2_X1  g267(.A(G2067), .B(G2678), .ZN(new_n693));
  XOR2_X1   g268(.A(G2084), .B(G2090), .Z(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT86), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n692), .A2(new_n693), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n698), .B(new_n695), .C1(new_n691), .C2(new_n693), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n694), .A2(new_n691), .A3(new_n693), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT18), .Z(new_n701));
  NAND3_X1  g276(.A1(new_n697), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(G2096), .B(G2100), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(G227));
  XOR2_X1   g279(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n705));
  XNOR2_X1  g280(.A(G1971), .B(G1976), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1956), .B(G2474), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1961), .B(G1966), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT20), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n708), .A2(new_n709), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n713), .A2(new_n710), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n712), .B(new_n714), .C1(new_n707), .C2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1981), .B(G1986), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT88), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n718), .B(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(G1991), .B(G1996), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(G229));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n724));
  MUX2_X1   g299(.A(G23), .B(G288), .S(G16), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT92), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT33), .B(G1976), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  MUX2_X1   g303(.A(G6), .B(G305), .S(G16), .Z(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT32), .B(G1981), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G22), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G166), .B2(new_n732), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G1971), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n728), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n737), .A2(KEYINPUT34), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(KEYINPUT34), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  MUX2_X1   g315(.A(G24), .B(G290), .S(G16), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1986), .ZN(new_n742));
  OAI21_X1  g317(.A(KEYINPUT89), .B1(G95), .B2(G2105), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NOR3_X1   g319(.A1(KEYINPUT89), .A2(G95), .A3(G2105), .ZN(new_n745));
  OAI221_X1 g320(.A(G2104), .B1(G107), .B2(new_n471), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n469), .A2(G131), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n485), .A2(G119), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  MUX2_X1   g324(.A(G25), .B(new_n749), .S(G29), .Z(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT35), .B(G1991), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT90), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT91), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n750), .B(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n742), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n724), .B1(new_n740), .B2(new_n755), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n724), .B(new_n755), .C1(new_n738), .C2(new_n739), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G29), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G35), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G162), .B2(new_n760), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT29), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G2090), .ZN(new_n764));
  NOR2_X1   g339(.A1(G29), .A2(G33), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT25), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n469), .A2(G139), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n478), .A2(new_n479), .A3(G127), .ZN(new_n770));
  INV_X1    g345(.A(G115), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(new_n462), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n769), .B1(new_n772), .B2(G2105), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n765), .B1(new_n773), .B2(G29), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G2072), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT96), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n774), .A2(G2072), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT94), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n764), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n763), .A2(G2090), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G29), .B2(G32), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n469), .A2(G141), .B1(G105), .B2(new_n463), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n485), .A2(G129), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT26), .Z(new_n786));
  NAND3_X1  g361(.A1(new_n783), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(new_n760), .ZN(new_n788));
  MUX2_X1   g363(.A(new_n782), .B(new_n781), .S(new_n788), .Z(new_n789));
  XOR2_X1   g364(.A(KEYINPUT27), .B(G1996), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n760), .A2(G26), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT28), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n469), .A2(G140), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n485), .A2(G128), .ZN(new_n795));
  OR2_X1    g370(.A1(G104), .A2(G2105), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n796), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n793), .B1(new_n799), .B2(new_n760), .ZN(new_n800));
  INV_X1    g375(.A(G2067), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT30), .B(G28), .ZN(new_n803));
  OR2_X1    g378(.A1(KEYINPUT31), .A2(G11), .ZN(new_n804));
  NAND2_X1  g379(.A1(KEYINPUT31), .A2(G11), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n803), .A2(new_n760), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n670), .B2(new_n760), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT100), .Z(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT95), .B(KEYINPUT24), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G34), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(G29), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G160), .B2(G29), .ZN(new_n812));
  INV_X1    g387(.A(G2084), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n791), .A2(new_n802), .A3(new_n808), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n732), .A2(G19), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT93), .Z(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n568), .B2(new_n732), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(G1341), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n760), .A2(G27), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G164), .B2(new_n760), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT104), .B(G2078), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n821), .B(new_n822), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  NOR4_X1   g399(.A1(new_n779), .A2(new_n780), .A3(new_n815), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(G5), .A2(G16), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT102), .Z(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n563), .B2(new_n732), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT103), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n829), .A2(G1961), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n829), .A2(G1961), .ZN(new_n831));
  NAND2_X1  g406(.A1(G168), .A2(G16), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT98), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(G16), .B2(G21), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(KEYINPUT98), .B2(new_n832), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT99), .Z(new_n837));
  AOI211_X1 g412(.A(new_n830), .B(new_n831), .C1(new_n837), .C2(G1966), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n732), .A2(G20), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT23), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n652), .B2(new_n732), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G1956), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n825), .A2(new_n838), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n837), .A2(G1966), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT101), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n732), .A2(G4), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n646), .B2(new_n732), .ZN(new_n848));
  INV_X1    g423(.A(G1348), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n844), .A2(new_n846), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n759), .A2(new_n851), .ZN(G311));
  AND2_X1   g427(.A1(new_n844), .A2(new_n846), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n853), .B(new_n850), .C1(new_n756), .C2(new_n758), .ZN(G150));
  NAND2_X1  g429(.A1(new_n646), .A2(G559), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT38), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n858));
  INV_X1    g433(.A(G93), .ZN(new_n859));
  OAI22_X1  g434(.A1(new_n858), .A2(new_n531), .B1(new_n524), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(new_n545), .B2(G55), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n568), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n857), .B(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(G860), .B1(new_n863), .B2(KEYINPUT39), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n568), .B(new_n861), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n857), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n855), .B(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n862), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT105), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT105), .ZN(new_n872));
  AOI211_X1 g447(.A(new_n872), .B(KEYINPUT39), .C1(new_n866), .C2(new_n868), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n864), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(G860), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n861), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(G145));
  NAND2_X1  g453(.A1(new_n773), .A2(KEYINPUT106), .ZN(new_n879));
  INV_X1    g454(.A(new_n787), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n497), .A2(new_n506), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n773), .A2(KEYINPUT106), .A3(new_n787), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n882), .B1(new_n881), .B2(new_n883), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n798), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n885), .A2(new_n798), .A3(new_n886), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n469), .A2(G142), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n485), .A2(G130), .ZN(new_n892));
  OR2_X1    g467(.A1(G106), .A2(G2105), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n893), .B(G2104), .C1(G118), .C2(new_n471), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n749), .B(KEYINPUT107), .ZN(new_n897));
  INV_X1    g472(.A(new_n662), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n898), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n896), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n901), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n904), .A2(new_n899), .A3(new_n895), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n906), .A3(KEYINPUT108), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT108), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n902), .B2(new_n905), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n890), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n907), .B(new_n909), .C1(new_n888), .C2(new_n889), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n490), .B(new_n670), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n914), .B(G160), .Z(new_n915));
  AOI21_X1  g490(.A(G37), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(new_n890), .B2(new_n910), .ZN(new_n917));
  OAI22_X1  g492(.A1(new_n888), .A2(new_n889), .B1(new_n905), .B2(new_n902), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n917), .A2(KEYINPUT109), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT109), .B1(new_n917), .B2(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(KEYINPUT110), .B(KEYINPUT40), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n921), .B(new_n922), .ZN(G395));
  NAND2_X1  g498(.A1(new_n657), .A2(new_n865), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n638), .A2(G299), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n644), .A2(new_n652), .A3(new_n626), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n646), .A2(new_n655), .A3(new_n862), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n924), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT41), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n925), .A2(new_n926), .A3(KEYINPUT41), .ZN(new_n932));
  AOI22_X1  g507(.A1(new_n924), .A2(new_n928), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT42), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(G290), .B(G305), .ZN(new_n935));
  XOR2_X1   g510(.A(G166), .B(G288), .Z(new_n936));
  OR2_X1    g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n936), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n931), .A2(new_n932), .ZN(new_n941));
  INV_X1    g516(.A(new_n928), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n862), .B1(new_n646), .B2(new_n655), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT42), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n924), .A2(new_n927), .A3(new_n928), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n934), .A2(new_n940), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n940), .B1(new_n934), .B2(new_n947), .ZN(new_n949));
  OAI21_X1  g524(.A(G868), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n950), .B1(G868), .B2(new_n861), .ZN(G295));
  OAI21_X1  g526(.A(new_n950), .B1(G868), .B2(new_n861), .ZN(G331));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n939), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n937), .A2(KEYINPUT112), .A3(new_n938), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n557), .A2(new_n559), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n957), .A2(KEYINPUT80), .A3(new_n562), .A4(new_n549), .ZN(new_n958));
  AOI21_X1  g533(.A(G286), .B1(new_n601), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(G171), .A2(G168), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n862), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n862), .B1(new_n959), .B2(new_n960), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT111), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n862), .B(new_n964), .C1(new_n959), .C2(new_n960), .ZN(new_n965));
  AOI211_X1 g540(.A(new_n927), .B(new_n961), .C1(new_n963), .C2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n959), .ZN(new_n967));
  INV_X1    g542(.A(new_n960), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n865), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n962), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n970), .A2(new_n931), .A3(new_n932), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n956), .B1(new_n966), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G37), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n969), .A2(new_n962), .A3(new_n925), .A4(new_n926), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n961), .B1(new_n963), .B2(new_n965), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n939), .B(new_n974), .C1(new_n975), .C2(new_n941), .ZN(new_n976));
  AND4_X1   g551(.A1(KEYINPUT43), .A2(new_n972), .A3(new_n973), .A4(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n976), .A2(new_n973), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n974), .B1(new_n975), .B2(new_n941), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n956), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT43), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT44), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  AND4_X1   g559(.A1(new_n984), .A2(new_n972), .A3(new_n973), .A4(new_n976), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n984), .B1(new_n978), .B2(new_n980), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n982), .A2(new_n987), .ZN(G397));
  NAND2_X1  g563(.A1(new_n480), .A2(new_n481), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(G2105), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n469), .A2(new_n465), .A3(G137), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n474), .A2(KEYINPUT69), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n991), .A2(new_n992), .B1(G101), .B2(new_n463), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n990), .A2(G40), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(G1384), .B1(new_n497), .B2(new_n506), .ZN(new_n995));
  XOR2_X1   g570(.A(KEYINPUT113), .B(KEYINPUT45), .Z(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n994), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1996), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT46), .ZN(new_n1001));
  INV_X1    g576(.A(new_n998), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n798), .B(new_n801), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n1003), .A2(new_n880), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1001), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT47), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT127), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n787), .B(new_n999), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n749), .A2(new_n752), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1003), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n799), .A2(new_n801), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1002), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(G290), .A2(G1986), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n998), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n1017), .A2(KEYINPUT48), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1011), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n749), .A2(new_n752), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1010), .A2(new_n1003), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n1017), .A2(KEYINPUT48), .B1(new_n1021), .B2(new_n998), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1014), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1008), .A2(new_n1009), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT63), .ZN(new_n1025));
  INV_X1    g600(.A(G1384), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(new_n507), .B2(new_n508), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n996), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT45), .ZN(new_n1029));
  AOI211_X1 g604(.A(new_n1029), .B(G1384), .C1(new_n497), .C2(new_n506), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(new_n994), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT114), .B(G1971), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n994), .B1(new_n1027), .B2(KEYINPUT50), .ZN(new_n1036));
  INV_X1    g611(.A(G2090), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n882), .A2(new_n1026), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT115), .B1(new_n1038), .B2(KEYINPUT50), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n995), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1036), .A2(new_n1037), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1035), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G8), .ZN(new_n1046));
  NOR2_X1   g621(.A1(G166), .A2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1047), .B(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1045), .A2(G8), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1049), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1033), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1041), .B1(new_n882), .B2(new_n1026), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(new_n994), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1041), .B(new_n1026), .C1(new_n507), .C2(new_n508), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1054), .A2(new_n1055), .A3(new_n1037), .ZN(new_n1056));
  OAI21_X1  g631(.A(G8), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1051), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1981), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n613), .A2(new_n616), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n615), .B1(new_n523), .B2(G61), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(new_n531), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n611), .A2(new_n612), .ZN(new_n1063));
  OAI21_X1  g638(.A(G1981), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT49), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(G8), .B1(new_n994), .B2(new_n1038), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1060), .A2(new_n1064), .A3(KEYINPUT49), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n607), .A2(new_n608), .A3(new_n609), .A4(G1976), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1070), .B(KEYINPUT117), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT52), .B1(new_n1072), .B2(new_n1066), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1066), .ZN(new_n1074));
  INV_X1    g649(.A(G1976), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT52), .B1(G288), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1074), .A2(new_n1071), .A3(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1069), .A2(new_n1073), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1050), .A2(new_n1058), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G40), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n476), .A2(new_n482), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1081), .B(new_n1082), .C1(KEYINPUT45), .C2(new_n995), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT45), .B1(new_n882), .B2(new_n1026), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT120), .B1(new_n1084), .B2(new_n994), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1026), .B(new_n997), .C1(new_n507), .C2(new_n508), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1966), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1036), .A2(new_n813), .A3(new_n1043), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(G8), .A3(G168), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1025), .B1(new_n1079), .B2(new_n1092), .ZN(new_n1093));
  AND4_X1   g668(.A1(KEYINPUT63), .A2(new_n1091), .A3(G8), .A4(G168), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1045), .A2(G8), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1051), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1094), .A2(new_n1050), .A3(new_n1096), .A4(new_n1078), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1066), .B(KEYINPUT118), .ZN(new_n1098));
  OR2_X1    g673(.A1(G288), .A2(G1976), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1060), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1098), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1069), .A2(new_n1073), .A3(new_n1077), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1102), .B1(new_n1050), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1102), .B(KEYINPUT119), .C1(new_n1050), .C2(new_n1103), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1093), .A2(new_n1097), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n1032), .B2(G2078), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1109), .A2(G2078), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1083), .A2(new_n1085), .A3(new_n1086), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(G1961), .B1(new_n1036), .B2(new_n1043), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1112), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G1961), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT72), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n882), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n497), .A2(new_n506), .A3(KEYINPUT72), .ZN(new_n1121));
  AOI21_X1  g696(.A(G1384), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1081), .B1(new_n1122), .B2(new_n1041), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1042), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1040), .B1(new_n995), .B2(new_n1041), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1118), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(KEYINPUT124), .A3(new_n1114), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1111), .B1(new_n1117), .B2(new_n1128), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1079), .A2(new_n1129), .A3(G301), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1089), .A2(G168), .A3(new_n1090), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(new_n1132), .A3(G8), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(G168), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(G8), .A3(new_n1131), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1134), .B1(new_n1137), .B2(KEYINPUT51), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1130), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1131), .A2(G8), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT51), .B1(new_n1141), .B2(new_n1135), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1142), .A2(new_n1139), .A3(new_n1133), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1108), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1146));
  INV_X1    g721(.A(G1956), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT56), .B(G2072), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1028), .A2(new_n1031), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT57), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n578), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n650), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n652), .B2(new_n1152), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1151), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1158), .A2(new_n1155), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1159));
  OAI211_X1 g734(.A(KEYINPUT122), .B(KEYINPUT61), .C1(new_n1157), .C2(new_n1159), .ZN(new_n1160));
  AOI22_X1  g735(.A1(G299), .A2(KEYINPUT57), .B1(new_n650), .B2(new_n1154), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1161), .A2(KEYINPUT122), .A3(new_n1148), .A4(new_n1150), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1151), .A2(KEYINPUT122), .A3(new_n1156), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1160), .A2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1031), .B(new_n999), .C1(new_n1122), .C2(new_n997), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n1168));
  XOR2_X1   g743(.A(KEYINPUT58), .B(G1341), .Z(new_n1169));
  OAI21_X1  g744(.A(new_n1169), .B1(new_n994), .B2(new_n1038), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n1167), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1168), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n568), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(KEYINPUT59), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT59), .ZN(new_n1175));
  OAI211_X1 g750(.A(new_n1175), .B(new_n568), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1036), .A2(new_n1043), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n849), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n994), .A2(new_n1038), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n801), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1179), .A2(KEYINPUT60), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1182), .A2(new_n640), .A3(new_n645), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT60), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI22_X1  g761(.A1(new_n1178), .A2(new_n849), .B1(new_n801), .B2(new_n1180), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n646), .A2(KEYINPUT60), .A3(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1183), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1166), .A2(new_n1177), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1157), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1187), .B1(new_n640), .B2(new_n645), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1191), .B1(new_n1192), .B2(new_n1159), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1145), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(G2078), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1195), .A2(KEYINPUT126), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1195), .A2(KEYINPUT126), .ZN(new_n1197));
  NOR4_X1   g772(.A1(new_n1030), .A2(new_n1109), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n994), .B1(new_n1038), .B2(new_n996), .ZN(new_n1199));
  AND2_X1   g774(.A1(new_n1199), .A2(KEYINPUT125), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1199), .A2(KEYINPUT125), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1198), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1202), .A2(new_n1110), .A3(G301), .A4(new_n1127), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1203), .B1(new_n1129), .B2(G301), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT54), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1129), .A2(G301), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1202), .A2(new_n1110), .A3(new_n1127), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1205), .B1(new_n1208), .B2(G171), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1079), .B1(new_n1142), .B2(new_n1133), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1206), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1194), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1190), .A2(new_n1145), .A3(new_n1193), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1144), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n1015), .A2(new_n1021), .ZN(new_n1216));
  NAND2_X1  g791(.A1(G290), .A2(G1986), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1002), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1024), .B1(new_n1215), .B2(new_n1218), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g794(.A1(G227), .A2(new_n460), .ZN(new_n1221));
  NOR3_X1   g795(.A1(G229), .A2(G401), .A3(new_n1221), .ZN(new_n1222));
  OAI211_X1 g796(.A(new_n921), .B(new_n1222), .C1(new_n985), .C2(new_n986), .ZN(G225));
  INV_X1    g797(.A(G225), .ZN(G308));
endmodule


