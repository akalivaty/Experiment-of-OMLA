//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n537, new_n538, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n555, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n611, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XNOR2_X1  g029(.A(G325), .B(KEYINPUT65), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(G2105), .ZN(new_n457));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n462));
  AND3_X1   g037(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n462), .B1(new_n459), .B2(new_n461), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n457), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n458), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n470), .B1(new_n460), .B2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n458), .A2(KEYINPUT67), .A3(KEYINPUT3), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n471), .A2(new_n472), .A3(new_n457), .A4(new_n461), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n467), .A2(new_n475), .ZN(G160));
  NAND4_X1  g051(.A1(new_n471), .A2(new_n472), .A3(G2105), .A4(new_n461), .ZN(new_n477));
  INV_X1    g052(.A(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n457), .A2(G112), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  OAI22_X1  g055(.A1(new_n477), .A2(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n473), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(G136), .B2(new_n482), .ZN(G162));
  AND2_X1   g058(.A1(G126), .A2(G2105), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n471), .A2(new_n472), .A3(new_n461), .A4(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR3_X1   g065(.A1(new_n490), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n463), .B2(new_n464), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n490), .A2(G2105), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n471), .A2(new_n472), .A3(new_n493), .A4(new_n461), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n489), .B1(new_n492), .B2(new_n495), .ZN(G164));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  XNOR2_X1  g072(.A(KEYINPUT5), .B(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G62), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(KEYINPUT68), .B1(G75), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n498), .A2(new_n501), .A3(G62), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n497), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n503), .A2(new_n509), .ZN(G166));
  NAND3_X1  g085(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n511));
  XNOR2_X1  g086(.A(new_n511), .B(KEYINPUT7), .ZN(new_n512));
  INV_X1    g087(.A(G51), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n504), .A2(G89), .ZN(new_n518));
  NAND2_X1  g093(.A1(G63), .A2(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n514), .A2(new_n520), .ZN(G168));
  NAND3_X1  g096(.A1(new_n498), .A2(new_n504), .A3(G90), .ZN(new_n522));
  INV_X1    g097(.A(G52), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n523), .B2(new_n507), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n498), .A2(G64), .ZN(new_n525));
  NAND2_X1  g100(.A1(G77), .A2(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n497), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(G171));
  AOI22_X1  g103(.A1(new_n498), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n497), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n504), .A2(G43), .A3(G543), .ZN(new_n531));
  INV_X1    g106(.A(G81), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n505), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G860), .ZN(G153));
  NAND4_X1  g110(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g111(.A1(G1), .A2(G3), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT8), .ZN(new_n538));
  NAND4_X1  g113(.A1(G319), .A2(G483), .A3(G661), .A4(new_n538), .ZN(G188));
  AND2_X1   g114(.A1(new_n504), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G53), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n541), .B1(KEYINPUT69), .B2(KEYINPUT9), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n540), .B(new_n542), .C1(KEYINPUT69), .C2(KEYINPUT9), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT69), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT9), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n544), .B(new_n545), .C1(new_n507), .C2(new_n541), .ZN(new_n546));
  NAND2_X1  g121(.A1(G78), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G65), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n517), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n498), .A2(new_n504), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G91), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n543), .A2(new_n546), .A3(new_n550), .A4(new_n552), .ZN(G299));
  INV_X1    g128(.A(G171), .ZN(G301));
  AOI22_X1  g129(.A1(new_n504), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n555));
  OAI221_X1 g130(.A(new_n512), .B1(new_n507), .B2(new_n513), .C1(new_n555), .C2(new_n517), .ZN(G286));
  INV_X1    g131(.A(G166), .ZN(G303));
  OAI21_X1  g132(.A(G651), .B1(new_n498), .B2(G74), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n504), .A2(G49), .A3(G543), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT70), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n551), .A2(G87), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(G288));
  INV_X1    g139(.A(KEYINPUT72), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n498), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n566), .B2(new_n497), .ZN(new_n567));
  OAI21_X1  g142(.A(G61), .B1(new_n515), .B2(new_n516), .ZN(new_n568));
  NAND2_X1  g143(.A1(G73), .A2(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n570), .A2(KEYINPUT72), .A3(G651), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n551), .A2(G86), .ZN(new_n572));
  AND2_X1   g147(.A1(KEYINPUT6), .A2(G651), .ZN(new_n573));
  NOR2_X1   g148(.A1(KEYINPUT6), .A2(G651), .ZN(new_n574));
  OAI211_X1 g149(.A(G48), .B(G543), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT73), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n504), .A2(KEYINPUT73), .A3(G48), .A4(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n567), .A2(new_n571), .A3(new_n572), .A4(new_n579), .ZN(G305));
  INV_X1    g155(.A(G85), .ZN(new_n581));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n505), .A2(new_n581), .B1(new_n507), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n498), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n497), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n551), .A2(KEYINPUT10), .A3(G92), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  INV_X1    g165(.A(G92), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n505), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n517), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(G651), .A2(new_n596), .B1(new_n540), .B2(G54), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n588), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n588), .B1(new_n599), .B2(G868), .ZN(G321));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(G299), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n602), .B2(G168), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT74), .Z(G297));
  XOR2_X1   g180(.A(new_n604), .B(KEYINPUT75), .Z(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n599), .B1(new_n607), .B2(G860), .ZN(G148));
  OAI21_X1  g183(.A(KEYINPUT76), .B1(new_n534), .B2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n599), .A2(new_n607), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  MUX2_X1   g186(.A(KEYINPUT76), .B(new_n609), .S(new_n611), .Z(G323));
  XNOR2_X1  g187(.A(KEYINPUT77), .B(KEYINPUT11), .ZN(new_n613));
  XNOR2_X1  g188(.A(G323), .B(new_n613), .ZN(G282));
  NOR2_X1   g189(.A1(new_n460), .A2(G2104), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n616));
  OAI21_X1  g191(.A(KEYINPUT66), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n468), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT13), .Z(new_n623));
  INV_X1    g198(.A(G2100), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  OR2_X1    g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n627), .B(G2104), .C1(G111), .C2(new_n457), .ZN(new_n628));
  INV_X1    g203(.A(G123), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n477), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(G135), .B2(new_n482), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2096), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n625), .A2(new_n626), .A3(new_n632), .ZN(G156));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT80), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2427), .B(G2430), .Z(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT81), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G1341), .ZN(new_n643));
  INV_X1    g218(.A(G1348), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(G1341), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n642), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n645), .A2(new_n648), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(G14), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n653), .B1(new_n645), .B2(new_n648), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(G401));
  INV_X1    g232(.A(KEYINPUT18), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n658), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n624), .ZN(new_n665));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n661), .B2(KEYINPUT18), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(G2096), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1981), .B(G1986), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n675), .A2(new_n676), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n674), .A2(new_n679), .A3(new_n677), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n674), .A2(new_n679), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n682));
  AOI211_X1 g257(.A(new_n678), .B(new_n680), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1991), .B(G1996), .Z(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n683), .A2(new_n684), .A3(new_n686), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n690), .B1(new_n688), .B2(new_n691), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n671), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n694), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n696), .A2(new_n670), .A3(new_n692), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n695), .A2(new_n697), .ZN(G229));
  MUX2_X1   g273(.A(G23), .B(G288), .S(G16), .Z(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT33), .B(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(G6), .A2(G16), .ZN(new_n702));
  INV_X1    g277(.A(G305), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(G16), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT32), .B(G1981), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(G16), .A2(G22), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G166), .B2(G16), .ZN(new_n708));
  INV_X1    g283(.A(G1971), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  AND3_X1   g285(.A1(new_n701), .A2(new_n706), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT34), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G24), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n586), .B2(new_n715), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1986), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G25), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT83), .Z(new_n721));
  AND2_X1   g296(.A1(new_n482), .A2(G131), .ZN(new_n722));
  OR2_X1    g297(.A1(G95), .A2(G2105), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n723), .B(G2104), .C1(G107), .C2(new_n457), .ZN(new_n724));
  INV_X1    g299(.A(G119), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n477), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n721), .B1(new_n727), .B2(new_n719), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT35), .B(G1991), .Z(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n728), .A2(new_n730), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n718), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n713), .A2(new_n714), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT36), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n715), .A2(G5), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G171), .B2(new_n715), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(G1961), .ZN(new_n738));
  NOR2_X1   g313(.A1(G16), .A2(G19), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n534), .B2(G16), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT84), .B(G1341), .Z(new_n741));
  AOI21_X1  g316(.A(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n740), .B2(new_n741), .ZN(new_n743));
  NOR2_X1   g318(.A1(G4), .A2(G16), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n599), .B2(G16), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1348), .ZN(new_n746));
  INV_X1    g321(.A(G34), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n747), .A2(KEYINPUT24), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(KEYINPUT24), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n719), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G160), .B2(new_n719), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G2084), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n743), .A2(new_n746), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G29), .A2(G35), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G162), .B2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT29), .B(G2090), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n715), .A2(G20), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT23), .Z(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G299), .B2(G16), .ZN(new_n760));
  INV_X1    g335(.A(G1956), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n719), .A2(G32), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT26), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n766), .A2(new_n767), .B1(G105), .B2(new_n468), .ZN(new_n768));
  INV_X1    g343(.A(G129), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n477), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n482), .A2(G141), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n763), .B1(new_n772), .B2(new_n719), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT27), .Z(new_n774));
  AOI211_X1 g349(.A(new_n757), .B(new_n762), .C1(new_n774), .C2(G1996), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n719), .A2(G33), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n457), .A2(G103), .A3(G2104), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT25), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G139), .B2(new_n482), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n619), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(new_n457), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n776), .B1(new_n782), .B2(new_n719), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G2072), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n719), .A2(G27), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G164), .B2(new_n719), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2078), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n774), .A2(G1996), .ZN(new_n789));
  AND4_X1   g364(.A1(new_n753), .A2(new_n775), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n719), .A2(G26), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT28), .ZN(new_n792));
  INV_X1    g367(.A(G128), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n477), .A2(new_n793), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT85), .Z(new_n795));
  OAI21_X1  g370(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n796));
  INV_X1    g371(.A(G116), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G2105), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n482), .B2(G140), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n792), .B1(new_n801), .B2(new_n719), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT86), .ZN(new_n803));
  INV_X1    g378(.A(G2067), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n715), .A2(G21), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G168), .B2(new_n715), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT87), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(G1966), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT88), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n631), .A2(G29), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT31), .B(G11), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT89), .ZN(new_n813));
  INV_X1    g388(.A(G28), .ZN(new_n814));
  AOI21_X1  g389(.A(G29), .B1(new_n814), .B2(KEYINPUT30), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(KEYINPUT30), .B2(new_n814), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n811), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT90), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n737), .A2(G1961), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n808), .A2(G1966), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n810), .A2(new_n818), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT91), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n735), .A2(new_n790), .A3(new_n805), .A4(new_n822), .ZN(G150));
  INV_X1    g398(.A(G150), .ZN(G311));
  INV_X1    g399(.A(G67), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n517), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(G80), .A2(G543), .ZN(new_n827));
  OAI21_X1  g402(.A(G651), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n551), .A2(G93), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT93), .B(G55), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n540), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n828), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G860), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT97), .B(KEYINPUT37), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT94), .ZN(new_n836));
  INV_X1    g411(.A(G93), .ZN(new_n837));
  INV_X1    g412(.A(new_n830), .ZN(new_n838));
  OAI22_X1  g413(.A1(new_n505), .A2(new_n837), .B1(new_n507), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n827), .B1(new_n498), .B2(G67), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n840), .A2(new_n497), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n836), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n828), .A2(new_n829), .A3(new_n831), .A4(KEYINPUT94), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n842), .A2(new_n843), .A3(new_n534), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n832), .B(new_n836), .C1(new_n530), .C2(new_n533), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT95), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n599), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  XOR2_X1   g424(.A(KEYINPUT92), .B(KEYINPUT38), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT96), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(G860), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n851), .B2(KEYINPUT39), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n835), .B1(new_n854), .B2(new_n856), .ZN(G145));
  INV_X1    g432(.A(KEYINPUT100), .ZN(new_n858));
  INV_X1    g433(.A(G37), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n489), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n485), .A2(KEYINPUT98), .A3(new_n488), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n861), .A2(new_n862), .B1(new_n492), .B2(new_n495), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(new_n795), .B2(new_n799), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n772), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n795), .A2(new_n799), .A3(new_n863), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n866), .B1(new_n865), .B2(new_n867), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n781), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n872), .A2(new_n782), .A3(new_n868), .ZN(new_n873));
  INV_X1    g448(.A(new_n622), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n727), .ZN(new_n875));
  OR2_X1    g450(.A1(G106), .A2(G2105), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n876), .B(G2104), .C1(G118), .C2(new_n457), .ZN(new_n877));
  INV_X1    g452(.A(G130), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n477), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(G142), .B2(new_n482), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n622), .B1(new_n722), .B2(new_n726), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n875), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n880), .B1(new_n875), .B2(new_n881), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n871), .A2(new_n873), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(G160), .B(new_n631), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(G162), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT99), .ZN(new_n889));
  INV_X1    g464(.A(new_n882), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n889), .B1(new_n890), .B2(new_n883), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n884), .A2(KEYINPUT99), .A3(new_n882), .ZN(new_n892));
  AOI22_X1  g467(.A1(new_n871), .A2(new_n873), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n859), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n871), .A2(new_n873), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n891), .A2(new_n892), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n871), .A2(new_n873), .A3(new_n892), .A4(new_n891), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n887), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n858), .B1(new_n894), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n887), .ZN(new_n901));
  INV_X1    g476(.A(new_n898), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n901), .B1(new_n902), .B2(new_n893), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n897), .A2(new_n887), .A3(new_n885), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n903), .A2(new_n904), .A3(KEYINPUT100), .A4(new_n859), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n900), .A2(KEYINPUT40), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT40), .B1(new_n900), .B2(new_n905), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(G395));
  OR2_X1    g483(.A1(new_n703), .A2(G288), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n703), .A2(G288), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(G166), .B(G290), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(G166), .B(new_n586), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n909), .A3(new_n910), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n919), .A2(KEYINPUT103), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(KEYINPUT103), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n916), .A2(KEYINPUT42), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n610), .B(KEYINPUT101), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n844), .A2(new_n845), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n925), .B(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT41), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n598), .A2(G299), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n598), .A2(G299), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n598), .A2(G299), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n598), .A2(G299), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(KEYINPUT41), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n927), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n929), .A2(new_n930), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n927), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n924), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n924), .A3(new_n938), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n923), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n939), .B1(new_n923), .B2(new_n940), .ZN(new_n942));
  OAI21_X1  g517(.A(G868), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n832), .A2(new_n602), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(G295));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n944), .ZN(G331));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n525), .A2(new_n526), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(G651), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n540), .A2(G52), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT105), .A4(new_n522), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(new_n524), .B2(new_n527), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(new_n954), .A3(G286), .ZN(new_n955));
  NAND3_X1  g530(.A1(G171), .A2(G168), .A3(KEYINPUT105), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n846), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n844), .A2(new_n955), .A3(new_n845), .A4(new_n956), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n958), .A2(new_n937), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n955), .A2(new_n956), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(new_n926), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n959), .A2(KEYINPUT106), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n958), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n931), .A2(new_n934), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n960), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(G37), .B1(new_n967), .B2(new_n916), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n926), .A2(new_n962), .A3(new_n961), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n959), .A2(KEYINPUT106), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n958), .A2(new_n937), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n958), .A2(new_n959), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n971), .A2(new_n972), .B1(new_n966), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT107), .B1(new_n974), .B2(new_n916), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT107), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n971), .A2(new_n972), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n935), .B1(new_n958), .B2(new_n959), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n976), .B(new_n917), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n968), .A2(KEYINPUT43), .A3(new_n975), .A4(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n981));
  INV_X1    g556(.A(new_n960), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n846), .A2(new_n957), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n983), .B1(new_n969), .B2(new_n970), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n982), .B(new_n916), .C1(new_n984), .C2(new_n935), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n859), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n965), .A2(new_n966), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n916), .B1(new_n987), .B2(new_n982), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n981), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n948), .B1(new_n980), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n968), .A2(new_n981), .A3(new_n975), .A4(new_n979), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT43), .B1(new_n986), .B2(new_n988), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n948), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n947), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT44), .B1(new_n992), .B2(new_n993), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n990), .A2(new_n997), .A3(KEYINPUT108), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n996), .A2(new_n998), .ZN(G397));
  INV_X1    g574(.A(KEYINPUT63), .ZN(new_n1000));
  XNOR2_X1  g575(.A(KEYINPUT109), .B(G1384), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n485), .A2(KEYINPUT98), .A3(new_n488), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT98), .B1(new_n485), .B2(new_n488), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n619), .A2(new_n491), .B1(KEYINPUT4), .B2(new_n494), .ZN(new_n1005));
  OAI211_X1 g580(.A(KEYINPUT45), .B(new_n1001), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G40), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n467), .A2(new_n1007), .A3(new_n475), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(G164), .B2(G1384), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1006), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n709), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT112), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(new_n1014), .A3(new_n709), .ZN(new_n1015));
  INV_X1    g590(.A(G2090), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n1017));
  INV_X1    g592(.A(new_n491), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1018), .B1(new_n617), .B2(new_n618), .ZN(new_n1019));
  OAI22_X1  g594(.A1(new_n1002), .A2(new_n1003), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1384), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT50), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  NOR3_X1   g598(.A1(G164), .A2(new_n1023), .A3(G1384), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1016), .B(new_n1008), .C1(new_n1022), .C2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1013), .A2(new_n1015), .A3(new_n1025), .ZN(new_n1026));
  OAI211_X1 g601(.A(KEYINPUT55), .B(G8), .C1(new_n503), .C2(new_n509), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1027), .A2(KEYINPUT113), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(KEYINPUT113), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n1030));
  INV_X1    g605(.A(G8), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1030), .B1(G166), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1026), .A2(G8), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1033), .ZN(new_n1035));
  INV_X1    g610(.A(new_n489), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(new_n1023), .A3(new_n1021), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1008), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1023), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1041), .A2(new_n1016), .B1(new_n709), .B2(new_n1011), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1035), .B1(new_n1042), .B2(new_n1031), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n567), .A2(new_n1044), .A3(new_n571), .ZN(new_n1045));
  NAND3_X1  g620(.A1(G305), .A2(G1981), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT72), .B1(new_n570), .B2(G651), .ZN(new_n1047));
  AOI211_X1 g622(.A(new_n565), .B(new_n497), .C1(new_n568), .C2(new_n569), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n577), .A2(new_n578), .B1(new_n551), .B2(G86), .ZN(new_n1050));
  INV_X1    g625(.A(G1981), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1049), .B(new_n1050), .C1(new_n1044), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1046), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT49), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n863), .A2(G1384), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1031), .B1(new_n1056), .B2(new_n1008), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1046), .A2(new_n1052), .A3(KEYINPUT49), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1060));
  INV_X1    g635(.A(new_n475), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n619), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n1062));
  OAI211_X1 g637(.A(G40), .B(new_n1061), .C1(new_n1062), .C2(new_n457), .ZN(new_n1063));
  OAI21_X1  g638(.A(G8), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1976), .ZN(new_n1065));
  NOR2_X1   g640(.A1(G288), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT52), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n560), .A2(new_n562), .A3(G1976), .A4(new_n563), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT52), .B1(G288), .B2(new_n1065), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1057), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1059), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1034), .A2(new_n1043), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G2084), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(new_n1008), .C1(new_n1022), .C2(new_n1024), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT45), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1075));
  NOR3_X1   g650(.A1(G164), .A2(new_n1009), .A3(G1384), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n1075), .A2(new_n1076), .A3(new_n1063), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1074), .B1(new_n1077), .B2(G1966), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1078), .A2(G8), .A3(G168), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1000), .B1(new_n1072), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1000), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1081), .A2(new_n1034), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1059), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1059), .A2(new_n1067), .A3(new_n1070), .A4(KEYINPUT115), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1026), .A2(G8), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1085), .A2(new_n1086), .B1(new_n1087), .B2(new_n1035), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1082), .B1(new_n1088), .B2(KEYINPUT118), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n1035), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1090), .A2(KEYINPUT118), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1080), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1034), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n560), .A2(new_n562), .A3(new_n1065), .A4(new_n563), .ZN(new_n1097));
  XOR2_X1   g672(.A(new_n1097), .B(KEYINPUT116), .Z(new_n1098));
  AOI21_X1  g673(.A(new_n1064), .B1(new_n1054), .B2(new_n1053), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1099), .B2(new_n1058), .ZN(new_n1100));
  NOR2_X1   g675(.A1(G305), .A2(G1981), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1096), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1101), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1059), .ZN(new_n1104));
  OAI211_X1 g679(.A(KEYINPUT117), .B(new_n1103), .C1(new_n1104), .C2(new_n1098), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(new_n1105), .A3(new_n1057), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1095), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1008), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1961), .ZN(new_n1111));
  OAI211_X1 g686(.A(KEYINPUT121), .B(new_n1008), .C1(new_n1022), .C2(new_n1024), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1114), .A2(G2078), .ZN(new_n1115));
  INV_X1    g690(.A(G2078), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1006), .A2(new_n1008), .A3(new_n1116), .A4(new_n1010), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1077), .A2(new_n1115), .B1(new_n1117), .B2(new_n1114), .ZN(new_n1118));
  AOI21_X1  g693(.A(G301), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1034), .A2(new_n1119), .A3(new_n1043), .A4(new_n1071), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1074), .B(G168), .C1(new_n1077), .C2(G1966), .ZN(new_n1121));
  AND2_X1   g696(.A1(KEYINPUT124), .A2(G8), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT51), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1078), .A2(G8), .A3(G286), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT51), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1121), .A2(new_n1126), .A3(new_n1122), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1120), .B1(KEYINPUT62), .B2(new_n1128), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n1128), .A2(KEYINPUT62), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1107), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT57), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1132), .A2(KEYINPUT119), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(KEYINPUT119), .ZN(new_n1134));
  XOR2_X1   g709(.A(new_n1134), .B(KEYINPUT120), .Z(new_n1135));
  AND3_X1   g710(.A1(G299), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1135), .B1(G299), .B2(new_n1133), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n761), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT56), .B(G2072), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1006), .A2(new_n1008), .A3(new_n1010), .A4(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1138), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1110), .A2(new_n644), .A3(new_n1112), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1056), .A2(new_n804), .A3(new_n1008), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n599), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1139), .A2(new_n1138), .A3(new_n1141), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1143), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT45), .B1(new_n1037), .B2(new_n1021), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1150), .A2(new_n1063), .ZN(new_n1151));
  INV_X1    g726(.A(G1996), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1151), .A2(KEYINPUT122), .A3(new_n1152), .A4(new_n1006), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1006), .A2(new_n1008), .A3(new_n1152), .A4(new_n1010), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT122), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1056), .A2(new_n1008), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT58), .B(G1341), .Z(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1153), .A2(new_n1156), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n534), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT59), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT59), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1160), .A2(new_n1163), .A3(new_n534), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n598), .A2(KEYINPUT60), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1144), .A2(new_n1145), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n1168), .A2(KEYINPUT123), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1169), .B1(new_n1148), .B2(new_n1142), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1168), .A2(KEYINPUT123), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g747(.A(KEYINPUT123), .B(new_n1168), .C1(new_n1148), .C2(new_n1142), .ZN(new_n1173));
  AND4_X1   g748(.A1(new_n1165), .A2(new_n1167), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1147), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1146), .A2(new_n599), .ZN(new_n1176));
  OAI21_X1  g751(.A(KEYINPUT60), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1149), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1127), .A2(new_n1125), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1126), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1181), .A2(new_n1072), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1113), .A2(G301), .A3(new_n1118), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1117), .A2(new_n1114), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1020), .A2(new_n1001), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(new_n1009), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1186), .A2(new_n1008), .A3(new_n1006), .A4(new_n1115), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1113), .A2(new_n1189), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1110), .A2(new_n1112), .A3(KEYINPUT125), .A4(new_n1111), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1188), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g767(.A(KEYINPUT54), .B(new_n1183), .C1(new_n1192), .C2(G301), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1119), .B1(new_n1192), .B2(G301), .ZN(new_n1194));
  OAI211_X1 g769(.A(new_n1182), .B(new_n1193), .C1(KEYINPUT54), .C2(new_n1194), .ZN(new_n1195));
  OAI211_X1 g770(.A(new_n1093), .B(new_n1131), .C1(new_n1178), .C2(new_n1195), .ZN(new_n1196));
  OR3_X1    g771(.A1(new_n1186), .A2(KEYINPUT110), .A3(new_n1063), .ZN(new_n1197));
  OAI21_X1  g772(.A(KEYINPUT110), .B1(new_n1186), .B2(new_n1063), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1197), .A2(new_n1152), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(KEYINPUT111), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT111), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1197), .A2(new_n1201), .A3(new_n1152), .A4(new_n1198), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n866), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n800), .B(G2067), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n772), .A2(new_n1152), .ZN(new_n1205));
  OR2_X1    g780(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  AND2_X1   g781(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1207));
  AND2_X1   g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1203), .A2(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n727), .B(new_n729), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1207), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g787(.A(G1986), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n586), .B(new_n1213), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1212), .B1(new_n1207), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1196), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n727), .A2(new_n729), .ZN(new_n1217));
  XOR2_X1   g792(.A(new_n1217), .B(KEYINPUT126), .Z(new_n1218));
  NOR3_X1   g793(.A1(new_n1203), .A2(new_n1208), .A3(new_n1218), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n800), .A2(G2067), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1207), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1207), .A2(new_n1213), .A3(new_n586), .ZN(new_n1222));
  XNOR2_X1  g797(.A(new_n1222), .B(KEYINPUT48), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1223), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1224));
  INV_X1    g799(.A(KEYINPUT47), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1226));
  INV_X1    g801(.A(KEYINPUT46), .ZN(new_n1227));
  XNOR2_X1  g802(.A(new_n1226), .B(new_n1227), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1207), .B1(new_n866), .B2(new_n1204), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n1225), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g805(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1231));
  AOI21_X1  g806(.A(KEYINPUT46), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1232));
  OAI211_X1 g807(.A(new_n1225), .B(new_n1229), .C1(new_n1231), .C2(new_n1232), .ZN(new_n1233));
  INV_X1    g808(.A(new_n1233), .ZN(new_n1234));
  OAI211_X1 g809(.A(new_n1221), .B(new_n1224), .C1(new_n1230), .C2(new_n1234), .ZN(new_n1235));
  INV_X1    g810(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1216), .A2(new_n1236), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g812(.A(G319), .ZN(new_n1239));
  OR2_X1    g813(.A1(G227), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g814(.A(new_n1240), .B1(new_n695), .B2(new_n697), .ZN(new_n1241));
  OAI21_X1  g815(.A(new_n1241), .B1(new_n655), .B2(new_n656), .ZN(new_n1242));
  NAND2_X1  g816(.A1(new_n1242), .A2(KEYINPUT127), .ZN(new_n1243));
  INV_X1    g817(.A(KEYINPUT127), .ZN(new_n1244));
  OAI211_X1 g818(.A(new_n1241), .B(new_n1244), .C1(new_n655), .C2(new_n656), .ZN(new_n1245));
  NAND2_X1  g819(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g820(.A1(new_n900), .A2(new_n905), .ZN(new_n1247));
  NAND3_X1  g821(.A1(new_n1246), .A2(new_n1247), .A3(new_n994), .ZN(G225));
  INV_X1    g822(.A(G225), .ZN(G308));
endmodule


