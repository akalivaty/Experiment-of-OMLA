//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n543, new_n544,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1185, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT67), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(KEYINPUT68), .A2(G113), .A3(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n461), .B1(new_n471), .B2(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n462), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n473), .A2(new_n465), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n475), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n474), .A2(G137), .A3(new_n459), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND3_X1  g054(.A1(new_n474), .A2(G2105), .A3(new_n476), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n459), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  OAI22_X1  g058(.A1(new_n480), .A2(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n476), .A2(new_n473), .A3(new_n459), .A4(new_n465), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n484), .B1(G136), .B2(new_n486), .ZN(G162));
  NAND4_X1  g062(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n459), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT4), .A2(G138), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n485), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n476), .A2(new_n473), .A3(new_n465), .A4(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n492), .A2(new_n498), .ZN(G164));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G62), .ZN(new_n506));
  NAND2_X1  g081(.A1(G75), .A2(G543), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n500), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT71), .B(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n508), .A2(new_n509), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  INV_X1    g095(.A(new_n512), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n521), .A2(G89), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n523), .B(new_n525), .C1(new_n526), .C2(new_n514), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n522), .A2(new_n527), .ZN(G168));
  AOI22_X1  g103(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n500), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n512), .A2(new_n531), .B1(new_n514), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(G171));
  AOI22_X1  g109(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n500), .ZN(new_n536));
  INV_X1    g111(.A(G81), .ZN(new_n537));
  XOR2_X1   g112(.A(KEYINPUT73), .B(G43), .Z(new_n538));
  OAI22_X1  g113(.A1(new_n537), .A2(new_n512), .B1(new_n514), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n505), .B(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G65), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g124(.A1(G78), .A2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(G651), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OR3_X1    g127(.A1(new_n514), .A2(KEYINPUT9), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT9), .B1(new_n514), .B2(new_n552), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n553), .A2(new_n554), .B1(G91), .B2(new_n521), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(G299));
  INV_X1    g131(.A(G171), .ZN(G301));
  OR2_X1    g132(.A1(new_n522), .A2(new_n527), .ZN(G286));
  INV_X1    g133(.A(new_n514), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n521), .A2(G87), .B1(new_n559), .B2(G49), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(KEYINPUT75), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(KEYINPUT75), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(G288));
  INV_X1    g139(.A(G61), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(new_n503), .B2(new_n504), .ZN(new_n566));
  NAND2_X1  g141(.A1(G73), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n505), .A2(G86), .A3(new_n511), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n511), .A2(G48), .A3(G543), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  XOR2_X1   g147(.A(new_n572), .B(KEYINPUT76), .Z(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G305));
  AOI22_X1  g149(.A1(new_n521), .A2(G85), .B1(new_n559), .B2(G47), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n500), .B2(new_n576), .ZN(G290));
  INV_X1    g152(.A(G66), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n547), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g154(.A1(G79), .A2(G543), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n521), .A2(KEYINPUT10), .A3(G92), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT10), .ZN(new_n583));
  INV_X1    g158(.A(G92), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n512), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n582), .A2(new_n585), .B1(G54), .B2(new_n559), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n587), .A2(KEYINPUT77), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n587), .A2(KEYINPUT77), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(G868), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(G868), .B2(G171), .ZN(G284));
  XNOR2_X1  g168(.A(G284), .B(KEYINPUT78), .ZN(G321));
  NAND2_X1  g169(.A1(G286), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(G299), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G297));
  OAI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n590), .B1(new_n599), .B2(G860), .ZN(G148));
  NAND2_X1  g175(.A1(new_n590), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G868), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G868), .B2(new_n540), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g179(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n605));
  NOR3_X1   g180(.A1(new_n462), .A2(new_n464), .A3(G2105), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n605), .B(new_n606), .Z(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT13), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(G2100), .Z(new_n609));
  INV_X1    g184(.A(G123), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT80), .ZN(new_n611));
  NOR3_X1   g186(.A1(new_n611), .A2(new_n459), .A3(G111), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n459), .B2(G111), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n613), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n614));
  OAI22_X1  g189(.A1(new_n480), .A2(new_n610), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(G135), .B2(new_n486), .ZN(new_n616));
  XOR2_X1   g191(.A(KEYINPUT81), .B(G2096), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n609), .A2(new_n618), .ZN(G156));
  XNOR2_X1  g194(.A(G2427), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT15), .B(G2435), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n623), .A2(KEYINPUT14), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2451), .B(G2454), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT16), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n625), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(G2443), .B(G2446), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G1341), .B(G1348), .Z(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT82), .ZN(new_n633));
  OAI21_X1  g208(.A(G14), .B1(new_n630), .B2(new_n631), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n633), .A2(new_n634), .ZN(G401));
  INV_X1    g210(.A(KEYINPUT18), .ZN(new_n636));
  XOR2_X1   g211(.A(G2084), .B(G2090), .Z(new_n637));
  XNOR2_X1  g212(.A(G2067), .B(G2678), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT17), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n636), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2096), .B(G2100), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(new_n639), .B2(KEYINPUT18), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT83), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(G227));
  XOR2_X1   g223(.A(G1971), .B(G1976), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT19), .ZN(new_n650));
  XOR2_X1   g225(.A(G1956), .B(G2474), .Z(new_n651));
  XOR2_X1   g226(.A(G1961), .B(G1966), .Z(new_n652));
  AND2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n651), .A2(new_n652), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  MUX2_X1   g233(.A(new_n658), .B(new_n657), .S(new_n650), .Z(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1981), .B(G1986), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT85), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n662), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1991), .B(G1996), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G229));
  INV_X1    g242(.A(G16), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n668), .A2(G23), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(G288), .B2(G16), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT89), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT33), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(G6), .A2(G16), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n573), .B2(G16), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT32), .B(G1981), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(G16), .A2(G22), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(G166), .B2(G16), .ZN(new_n679));
  INV_X1    g254(.A(G1971), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n673), .A2(new_n677), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT88), .B(KEYINPUT34), .Z(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n486), .A2(G131), .ZN(new_n686));
  INV_X1    g261(.A(G119), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n459), .A2(G107), .ZN(new_n688));
  OAI21_X1  g263(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n689));
  OAI221_X1 g264(.A(new_n686), .B1(new_n480), .B2(new_n687), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT86), .B(G29), .Z(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G25), .B2(new_n696), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT35), .B(G1991), .Z(new_n699));
  AND2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  MUX2_X1   g276(.A(G24), .B(G290), .S(G16), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1986), .ZN(new_n703));
  NOR3_X1   g278(.A1(new_n700), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n682), .A2(new_n684), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n685), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G4), .A2(G16), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n590), .B2(G16), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G1348), .ZN(new_n711));
  INV_X1    g286(.A(new_n696), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(G35), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G162), .B2(new_n712), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT29), .ZN(new_n715));
  INV_X1    g290(.A(G2090), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n668), .A2(G20), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G299), .B2(G16), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1956), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT24), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(G34), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(G34), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n696), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n478), .B2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G2084), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT97), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n727), .A2(G32), .ZN(new_n732));
  NAND3_X1  g307(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT94), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT93), .B(KEYINPUT26), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G129), .ZN(new_n739));
  INV_X1    g314(.A(G141), .ZN(new_n740));
  OAI22_X1  g315(.A1(new_n480), .A2(new_n739), .B1(new_n740), .B2(new_n485), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n732), .B1(new_n742), .B2(new_n727), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT27), .B(G1996), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT95), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n743), .B(new_n745), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n717), .A2(new_n722), .A3(new_n731), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n727), .A2(G33), .ZN(new_n748));
  INV_X1    g323(.A(G139), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n485), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT91), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT25), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n463), .A2(new_n465), .A3(G127), .ZN(new_n755));
  INV_X1    g330(.A(G115), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(new_n464), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n754), .B1(G2105), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n752), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT92), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n748), .B1(new_n761), .B2(new_n727), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(G2072), .ZN(new_n763));
  NOR2_X1   g338(.A1(G171), .A2(new_n668), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G5), .B2(new_n668), .ZN(new_n765));
  INV_X1    g340(.A(G1961), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n668), .A2(G21), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G168), .B2(new_n668), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(G1966), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n540), .A2(G16), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G16), .B2(G19), .ZN(new_n772));
  INV_X1    g347(.A(G1341), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n769), .A2(G1966), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n767), .A2(new_n770), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT31), .B(G11), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT96), .ZN(new_n778));
  INV_X1    g353(.A(G28), .ZN(new_n779));
  AOI21_X1  g354(.A(G29), .B1(new_n779), .B2(KEYINPUT30), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(KEYINPUT30), .B2(new_n779), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n616), .B2(new_n712), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n728), .B2(new_n729), .ZN(new_n784));
  OAI22_X1  g359(.A1(new_n765), .A2(new_n766), .B1(new_n772), .B2(new_n773), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n776), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n762), .A2(G2072), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n696), .A2(G26), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT28), .ZN(new_n789));
  OR2_X1    g364(.A1(G104), .A2(G2105), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n790), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n791));
  INV_X1    g366(.A(G140), .ZN(new_n792));
  INV_X1    g367(.A(G128), .ZN(new_n793));
  OAI221_X1 g368(.A(new_n791), .B1(new_n792), .B2(new_n485), .C1(new_n480), .C2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n789), .B1(new_n795), .B2(new_n727), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G2067), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n712), .A2(G27), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G164), .B2(new_n712), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G2078), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n763), .A2(new_n786), .A3(new_n787), .A4(new_n801), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n711), .A2(new_n747), .A3(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n708), .A2(new_n804), .ZN(G311));
  INV_X1    g380(.A(G311), .ZN(G150));
  NAND2_X1  g381(.A1(new_n590), .A2(G559), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT38), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n505), .A2(G67), .ZN(new_n809));
  AND2_X1   g384(.A1(G80), .A2(G543), .ZN(new_n810));
  OAI21_X1  g385(.A(G651), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT99), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT100), .B(G93), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n521), .A2(new_n814), .B1(new_n559), .B2(G55), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n811), .A2(new_n812), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(new_n540), .ZN(new_n819));
  INV_X1    g394(.A(new_n540), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n816), .B2(new_n817), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n808), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n824));
  AOI21_X1  g399(.A(G860), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n824), .B2(new_n823), .ZN(new_n826));
  OAI21_X1  g401(.A(G860), .B1(new_n816), .B2(new_n817), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(G145));
  INV_X1    g404(.A(new_n607), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT101), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n498), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n491), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n474), .A2(new_n459), .A3(new_n476), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n494), .A2(KEYINPUT101), .A3(new_n497), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n832), .A2(new_n490), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n795), .A2(new_n836), .ZN(new_n837));
  AND3_X1   g412(.A1(new_n494), .A2(KEYINPUT101), .A3(new_n497), .ZN(new_n838));
  AOI21_X1  g413(.A(KEYINPUT101), .B1(new_n494), .B2(new_n497), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n492), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(new_n794), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n837), .A2(new_n742), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n742), .B1(new_n837), .B2(new_n841), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n761), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT102), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT102), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n761), .B(new_n847), .C1(new_n843), .C2(new_n844), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n759), .B(KEYINPUT92), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n837), .A2(new_n841), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n738), .A2(new_n741), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n850), .A2(new_n853), .A3(new_n842), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT103), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n850), .A2(new_n853), .A3(KEYINPUT103), .A4(new_n842), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n486), .A2(G142), .ZN(new_n859));
  INV_X1    g434(.A(G130), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT104), .ZN(new_n861));
  NOR3_X1   g436(.A1(new_n861), .A2(new_n459), .A3(G118), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n459), .B2(G118), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n863), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n864));
  OAI221_X1 g439(.A(new_n859), .B1(new_n480), .B2(new_n860), .C1(new_n862), .C2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n694), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n849), .A2(new_n858), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n867), .B1(new_n849), .B2(new_n858), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n830), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n849), .A2(new_n858), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n866), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n849), .A2(new_n858), .A3(new_n867), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n607), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n616), .B(new_n478), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(G162), .ZN(new_n877));
  AOI21_X1  g452(.A(G37), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n870), .A2(new_n874), .A3(new_n879), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n878), .A2(KEYINPUT40), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT40), .B1(new_n878), .B2(new_n880), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(G395));
  AND2_X1   g458(.A1(new_n819), .A2(new_n821), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n601), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(G299), .A2(new_n587), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n551), .A2(new_n581), .A3(new_n555), .A4(new_n586), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n886), .A2(KEYINPUT105), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n885), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n888), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n886), .A2(KEYINPUT41), .A3(new_n887), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n885), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n573), .B(G290), .ZN(new_n900));
  INV_X1    g475(.A(G288), .ZN(new_n901));
  XNOR2_X1  g476(.A(G303), .B(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n900), .B(new_n902), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n903), .B(KEYINPUT42), .Z(new_n904));
  AND3_X1   g479(.A1(new_n894), .A2(new_n899), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n894), .B2(new_n899), .ZN(new_n906));
  OAI21_X1  g481(.A(G868), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(G868), .B2(new_n818), .ZN(G295));
  OAI21_X1  g483(.A(new_n907), .B1(G868), .B2(new_n818), .ZN(G331));
  INV_X1    g484(.A(new_n903), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n911));
  NAND2_X1  g486(.A1(G286), .A2(G301), .ZN(new_n912));
  NAND2_X1  g487(.A1(G168), .A2(G171), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n884), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n913), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n822), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n911), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n822), .A2(new_n916), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(KEYINPUT106), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n918), .A2(new_n892), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n914), .B1(new_n821), .B2(new_n819), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n923), .A2(new_n898), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n910), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n926));
  INV_X1    g501(.A(G37), .ZN(new_n927));
  INV_X1    g502(.A(new_n898), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n918), .B2(new_n920), .ZN(new_n929));
  INV_X1    g504(.A(new_n888), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n923), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n931), .A3(new_n903), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n925), .A2(new_n926), .A3(new_n927), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT107), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n927), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT106), .B1(new_n919), .B2(new_n922), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n915), .A2(new_n911), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n938), .A2(new_n928), .B1(new_n930), .B2(new_n923), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n939), .A2(new_n903), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT43), .B1(new_n935), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(G37), .B1(new_n939), .B2(new_n903), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n942), .A2(new_n943), .A3(new_n926), .A4(new_n925), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n934), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n935), .A2(new_n940), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n942), .A2(KEYINPUT43), .A3(new_n925), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT44), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n947), .A2(new_n951), .ZN(G397));
  XNOR2_X1  g527(.A(new_n742), .B(G1996), .ZN(new_n953));
  INV_X1    g528(.A(G2067), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n794), .B(new_n954), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n695), .A2(new_n699), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n695), .A2(new_n699), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n469), .A2(new_n470), .ZN(new_n961));
  OAI21_X1  g536(.A(G2105), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n962), .A2(new_n477), .A3(G40), .A4(new_n460), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n472), .A2(KEYINPUT109), .A3(G40), .A4(new_n477), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n836), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n959), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(G290), .A2(G1986), .ZN(new_n974));
  AND2_X1   g549(.A1(G290), .A2(G1986), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n977), .B(KEYINPUT110), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT45), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n836), .A2(new_n980), .A3(new_n970), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n980), .B1(new_n836), .B2(new_n970), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G2078), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n970), .B(new_n969), .C1(new_n492), .C2(new_n498), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n965), .A2(new_n966), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n983), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT123), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT123), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n983), .A2(new_n989), .A3(new_n984), .A4(new_n986), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(KEYINPUT53), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT111), .B1(new_n840), .B2(G1384), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n836), .A2(new_n980), .A3(new_n970), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT50), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n970), .B1(new_n492), .B2(new_n498), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT50), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n967), .B1(new_n994), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n836), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n995), .A2(new_n968), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n967), .A2(new_n984), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n999), .A2(new_n766), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n991), .A2(G301), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1003), .A2(new_n1000), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n984), .A2(KEYINPUT124), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n984), .A2(KEYINPUT124), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1000), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1001), .A2(G40), .A3(G160), .A4(new_n1010), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n1011), .A2(new_n971), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n965), .A2(new_n966), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1014), .B1(new_n981), .B2(new_n982), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1013), .B1(new_n1015), .B2(new_n997), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1007), .B(new_n1012), .C1(new_n1016), .C2(G1961), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1006), .B1(new_n1017), .B2(G171), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1005), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT125), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1005), .A2(new_n1018), .A3(KEYINPUT125), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G8), .ZN(new_n1024));
  NOR2_X1   g599(.A1(G168), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n729), .B(new_n967), .C1(new_n994), .C2(new_n998), .ZN(new_n1027));
  INV_X1    g602(.A(G1966), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT45), .B1(new_n992), .B2(new_n993), .ZN(new_n1029));
  INV_X1    g604(.A(new_n986), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1026), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT51), .B1(new_n1025), .B2(KEYINPUT121), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n983), .A2(new_n986), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1016), .A2(new_n729), .B1(new_n1034), .B2(new_n1028), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1026), .B(new_n1033), .C1(new_n1035), .C2(new_n1024), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1033), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1038));
  OAI211_X1 g613(.A(G8), .B(new_n1037), .C1(new_n1038), .C2(G286), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1032), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n716), .B(new_n967), .C1(new_n994), .C2(new_n998), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1015), .A2(new_n997), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1044), .A2(KEYINPUT112), .A3(new_n716), .A4(new_n967), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n967), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n680), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G303), .A2(G8), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1049), .B(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1048), .A2(G8), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT50), .B1(new_n981), .B2(new_n982), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1013), .B1(new_n1014), .B2(new_n996), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n716), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1047), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1051), .B1(new_n1056), .B2(G8), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n967), .A2(new_n992), .A3(new_n993), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n901), .A2(G1976), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(G8), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT52), .ZN(new_n1061));
  INV_X1    g636(.A(G1976), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT52), .B1(G288), .B2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1058), .A2(new_n1059), .A3(new_n1063), .A4(G8), .ZN(new_n1064));
  INV_X1    g639(.A(G1981), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n569), .A2(new_n570), .A3(new_n1065), .A4(new_n571), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT49), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(KEYINPUT113), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(new_n1066), .B2(KEYINPUT113), .ZN(new_n1070));
  OAI211_X1 g645(.A(G1981), .B(new_n572), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1070), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n572), .A2(G1981), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(new_n1073), .A3(new_n1068), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1058), .A2(new_n1071), .A3(G8), .A4(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1061), .A2(new_n1064), .A3(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1057), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1052), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1040), .A2(new_n1078), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1080));
  AOI21_X1  g655(.A(G301), .B1(new_n991), .B2(new_n1004), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1017), .A2(G171), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1023), .A2(new_n1079), .A3(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT56), .B(G2072), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(KEYINPUT117), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1046), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT116), .B(G1956), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n967), .B1(KEYINPUT50), .B2(new_n995), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1014), .B1(new_n992), .B2(new_n993), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n551), .A2(new_n555), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1088), .A2(new_n1092), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1348), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n999), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1058), .A2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n981), .A2(new_n982), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(KEYINPUT118), .A3(new_n967), .ZN(new_n1104));
  AOI21_X1  g679(.A(G2067), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1100), .B1(new_n1105), .B2(KEYINPUT119), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT118), .B1(new_n1103), .B2(new_n967), .ZN(new_n1107));
  AND4_X1   g682(.A1(KEYINPUT118), .A2(new_n967), .A3(new_n992), .A4(new_n993), .ZN(new_n1108));
  OAI211_X1 g683(.A(KEYINPUT119), .B(new_n954), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n590), .B(new_n1098), .C1(new_n1106), .C2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1089), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1096), .B1(new_n1113), .B2(new_n1087), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n954), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1118), .A2(KEYINPUT60), .A3(new_n1109), .A4(new_n1100), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n591), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1116), .A2(new_n1117), .B1(new_n1099), .B2(new_n999), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1121), .A2(KEYINPUT60), .A3(new_n590), .A4(new_n1109), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT60), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1120), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT58), .B(G1341), .Z(new_n1126));
  NAND3_X1  g701(.A1(new_n1102), .A2(new_n1104), .A3(new_n1126), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1046), .A2(G1996), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1129), .A2(KEYINPUT120), .A3(new_n540), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT59), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1129), .A2(KEYINPUT120), .A3(new_n1132), .A4(new_n540), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1098), .A2(new_n1114), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT61), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1098), .A2(new_n1114), .A3(new_n1136), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1131), .A2(new_n1133), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1115), .B1(new_n1125), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1084), .A2(new_n1139), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1052), .A2(new_n1081), .A3(new_n1077), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1032), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT62), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n1145));
  AOI211_X1 g720(.A(new_n1145), .B(new_n1032), .C1(new_n1036), .C2(new_n1039), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1141), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1058), .A2(G8), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT114), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1075), .A2(new_n1062), .A3(new_n901), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1066), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(new_n1052), .B2(new_n1076), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT115), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g730(.A(KEYINPUT115), .B(new_n1152), .C1(new_n1052), .C2(new_n1076), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n1035), .A2(new_n1024), .A3(G286), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1052), .A2(new_n1077), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1051), .B1(new_n1048), .B2(G8), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT63), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1076), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1052), .A2(new_n1158), .A3(new_n1162), .ZN(new_n1163));
  OAI22_X1  g738(.A1(new_n1159), .A2(KEYINPUT63), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1147), .A2(new_n1157), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n978), .B1(new_n1140), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n972), .A2(new_n974), .ZN(new_n1167));
  XNOR2_X1  g742(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1170));
  AOI211_X1 g745(.A(new_n1169), .B(new_n1170), .C1(new_n959), .C2(new_n972), .ZN(new_n1171));
  INV_X1    g746(.A(G1996), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n972), .A2(new_n1172), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1173), .B(KEYINPUT46), .Z(new_n1174));
  NAND2_X1  g749(.A1(new_n955), .A2(new_n742), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n972), .A2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT126), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1174), .A2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT47), .ZN(new_n1179));
  INV_X1    g754(.A(new_n956), .ZN(new_n1180));
  OAI22_X1  g755(.A1(new_n1180), .A2(new_n958), .B1(G2067), .B2(new_n794), .ZN(new_n1181));
  AOI211_X1 g756(.A(new_n1171), .B(new_n1179), .C1(new_n972), .C2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1166), .A2(new_n1182), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g758(.A1(new_n878), .A2(new_n880), .ZN(new_n1185));
  INV_X1    g759(.A(G319), .ZN(new_n1186));
  NOR4_X1   g760(.A1(G229), .A2(G401), .A3(new_n1186), .A4(G227), .ZN(new_n1187));
  AND3_X1   g761(.A1(new_n1185), .A2(new_n945), .A3(new_n1187), .ZN(G308));
  NAND3_X1  g762(.A1(new_n1185), .A2(new_n945), .A3(new_n1187), .ZN(G225));
endmodule


