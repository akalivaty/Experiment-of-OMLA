//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  NAND3_X1  g001(.A1(new_n202), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT14), .B(G29gat), .Z(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(G36gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(G43gat), .B(G50gat), .ZN(new_n206));
  OR2_X1    g005(.A1(new_n206), .A2(KEYINPUT15), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT88), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n209), .B1(new_n206), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(new_n210), .B2(new_n206), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n205), .B(new_n211), .C1(new_n210), .C2(new_n206), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT17), .ZN(new_n216));
  XNOR2_X1  g015(.A(G15gat), .B(G22gat), .ZN(new_n217));
  INV_X1    g016(.A(G1gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT16), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G1gat), .B2(new_n217), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(G8gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n213), .A2(new_n224), .A3(new_n214), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n216), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G229gat), .A2(G233gat), .ZN(new_n227));
  INV_X1    g026(.A(new_n215), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(new_n222), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n226), .A2(KEYINPUT18), .A3(new_n227), .A4(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n227), .B(KEYINPUT13), .Z(new_n231));
  NOR2_X1   g030(.A1(new_n228), .A2(new_n222), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n223), .A2(new_n215), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G113gat), .B(G141gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G197gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT11), .B(G169gat), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT12), .Z(new_n240));
  NOR2_X1   g039(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT18), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT89), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT89), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n242), .A2(new_n246), .A3(new_n243), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n241), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n244), .A2(new_n234), .A3(new_n230), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n240), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT35), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT25), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT23), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(G169gat), .B2(G176gat), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n256), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n254), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G169gat), .ZN(new_n264));
  INV_X1    g063(.A(G176gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n266), .B1(KEYINPUT23), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n261), .A2(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n263), .B(new_n269), .Z(new_n270));
  INV_X1    g069(.A(KEYINPUT26), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n266), .B1(new_n271), .B2(new_n267), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n272), .B1(new_n271), .B2(new_n267), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n258), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(KEYINPUT66), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(KEYINPUT66), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT27), .B(G183gat), .ZN(new_n277));
  INV_X1    g076(.A(G190gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n280), .A2(KEYINPUT28), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n279), .B(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n270), .B1(new_n275), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT76), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G226gat), .A2(G233gat), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G211gat), .ZN(new_n291));
  INV_X1    g090(.A(G218gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(G197gat), .A2(G204gat), .ZN(new_n294));
  AND2_X1   g093(.A1(G197gat), .A2(G204gat), .ZN(new_n295));
  OAI22_X1  g094(.A1(new_n293), .A2(KEYINPUT22), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(KEYINPUT75), .ZN(new_n298));
  XOR2_X1   g097(.A(G211gat), .B(G218gat), .Z(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n290), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G8gat), .B(G36gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(G64gat), .B(G92gat), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n302), .B(new_n303), .Z(new_n304));
  OR2_X1    g103(.A1(new_n284), .A2(KEYINPUT76), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n284), .A2(KEYINPUT76), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n305), .A2(G226gat), .A3(G233gat), .A4(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n300), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n284), .A2(new_n286), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n301), .A2(new_n304), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n311), .B(KEYINPUT30), .ZN(new_n312));
  INV_X1    g111(.A(new_n304), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n301), .A2(new_n314), .A3(new_n310), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n314), .B1(new_n301), .B2(new_n310), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n313), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT82), .ZN(new_n319));
  INV_X1    g118(.A(G148gat), .ZN(new_n320));
  OR3_X1    g119(.A1(new_n320), .A2(KEYINPUT78), .A3(G141gat), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT78), .B1(new_n320), .B2(G141gat), .ZN(new_n322));
  INV_X1    g121(.A(G141gat), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n321), .B(new_n322), .C1(new_n323), .C2(G148gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(G155gat), .B(G162gat), .ZN(new_n325));
  INV_X1    g124(.A(G155gat), .ZN(new_n326));
  INV_X1    g125(.A(G162gat), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT2), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n329));
  OR2_X1    g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n329), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n324), .A2(new_n325), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G141gat), .B(G148gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(KEYINPUT2), .ZN(new_n334));
  OR2_X1    g133(.A1(new_n334), .A2(new_n325), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G127gat), .B(G134gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT67), .ZN(new_n339));
  INV_X1    g138(.A(G120gat), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n340), .A2(G113gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(G113gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n339), .B1(KEYINPUT1), .B2(new_n343), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n341), .A2(KEYINPUT68), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n341), .A2(KEYINPUT68), .ZN(new_n346));
  XOR2_X1   g145(.A(KEYINPUT69), .B(G113gat), .Z(new_n347));
  OAI211_X1 g146(.A(new_n345), .B(new_n346), .C1(new_n340), .C2(new_n347), .ZN(new_n348));
  OR2_X1    g147(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n349));
  NAND2_X1  g148(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n348), .A2(new_n338), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n337), .A2(new_n344), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n344), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT71), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n337), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n354), .B1(new_n357), .B2(new_n353), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT5), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n337), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n336), .A2(KEYINPUT3), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n362), .A3(new_n355), .ZN(new_n363));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n358), .A2(new_n359), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n352), .A2(new_n353), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n365), .B(new_n367), .C1(new_n357), .C2(new_n353), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n355), .A2(new_n336), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n352), .ZN(new_n370));
  INV_X1    g169(.A(new_n364), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n359), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n366), .A2(new_n373), .ZN(new_n374));
  XOR2_X1   g173(.A(G1gat), .B(G29gat), .Z(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(KEYINPUT81), .ZN(new_n376));
  XOR2_X1   g175(.A(G57gat), .B(G85gat), .Z(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  OAI21_X1  g179(.A(new_n319), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n380), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n382), .B1(new_n366), .B2(new_n373), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT6), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n366), .A2(new_n373), .A3(KEYINPUT82), .A4(new_n382), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n381), .A2(new_n384), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n383), .A2(KEYINPUT6), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n312), .A2(new_n318), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT83), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n312), .A2(new_n318), .A3(new_n389), .A4(KEYINPUT83), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT29), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n300), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n337), .B1(new_n396), .B2(new_n360), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n300), .B1(new_n361), .B2(new_n395), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G228gat), .A2(G233gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n297), .A2(new_n299), .ZN(new_n401));
  INV_X1    g200(.A(new_n299), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT29), .B1(new_n402), .B2(new_n296), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT3), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n400), .B1(new_n337), .B2(new_n404), .ZN(new_n405));
  OAI22_X1  g204(.A1(new_n399), .A2(new_n400), .B1(new_n398), .B2(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(KEYINPUT31), .B(G50gat), .Z(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(G22gat), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n408), .B(new_n410), .Z(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT71), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n355), .B(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(new_n284), .ZN(new_n415));
  AND2_X1   g214(.A1(G227gat), .A2(G233gat), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT34), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT73), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n416), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n420), .A2(KEYINPUT32), .ZN(new_n421));
  XNOR2_X1  g220(.A(G15gat), .B(G43gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(G71gat), .B(G99gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT33), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n419), .B1(new_n421), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n420), .A2(KEYINPUT32), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n429), .A2(KEYINPUT73), .A3(new_n426), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(KEYINPUT72), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT72), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n420), .A2(new_n433), .A3(KEYINPUT32), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n424), .B1(new_n420), .B2(new_n425), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n418), .B1(new_n431), .B2(new_n437), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n417), .B(KEYINPUT34), .Z(new_n439));
  OAI211_X1 g238(.A(new_n439), .B(new_n436), .C1(new_n428), .C2(new_n430), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT74), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(KEYINPUT74), .B(new_n418), .C1(new_n431), .C2(new_n437), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n412), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n253), .B1(new_n394), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n438), .A2(new_n440), .ZN(new_n446));
  NOR4_X1   g245(.A1(new_n390), .A2(new_n446), .A3(KEYINPUT35), .A4(new_n412), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n446), .A2(KEYINPUT36), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n442), .A2(KEYINPUT36), .A3(new_n443), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n392), .A2(new_n412), .A3(new_n393), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT37), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n301), .A2(new_n454), .A3(new_n310), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n304), .A2(KEYINPUT38), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT86), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n287), .A2(new_n308), .A3(new_n289), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n308), .B1(new_n307), .B2(new_n309), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n458), .B2(new_n459), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n457), .B1(new_n463), .B2(KEYINPUT37), .ZN(new_n464));
  AOI211_X1 g263(.A(KEYINPUT86), .B(new_n454), .C1(new_n460), .C2(new_n462), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n455), .B(new_n456), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n389), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n467), .A3(new_n311), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n301), .A2(new_n310), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT77), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n454), .B1(new_n470), .B2(new_n315), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT87), .B1(new_n471), .B2(new_n304), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT37), .B1(new_n316), .B2(new_n317), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT87), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n313), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n475), .A3(new_n455), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n468), .B1(KEYINPUT38), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT40), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n364), .B1(new_n358), .B2(new_n363), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT39), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT39), .B1(new_n370), .B2(new_n371), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n481), .B(new_n382), .C1(new_n479), .C2(new_n482), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n483), .A2(KEYINPUT84), .A3(new_n478), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT84), .B1(new_n483), .B2(new_n478), .ZN(new_n485));
  OAI221_X1 g284(.A(new_n384), .B1(new_n478), .B2(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n312), .A2(new_n318), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n411), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n452), .B(new_n453), .C1(new_n477), .C2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n252), .B1(new_n448), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g289(.A1(G232gat), .A2(G233gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(KEYINPUT41), .ZN(new_n492));
  XNOR2_X1  g291(.A(G134gat), .B(G162gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(G85gat), .A2(G92gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT7), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT97), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT8), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(G99gat), .B2(G106gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT8), .ZN(new_n505));
  OR2_X1    g304(.A1(G85gat), .A2(G92gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT97), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n498), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(G99gat), .B(G106gat), .Z(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT99), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT7), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n505), .A2(KEYINPUT97), .A3(new_n506), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT97), .B1(new_n505), .B2(new_n506), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT99), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(new_n509), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT100), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n510), .B(new_n512), .C1(new_n513), .C2(new_n514), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT98), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n507), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT98), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n522), .A2(new_n523), .A3(new_n510), .A4(new_n512), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n518), .A2(new_n519), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n519), .B1(new_n518), .B2(new_n525), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n528), .A2(new_n228), .B1(KEYINPUT41), .B2(new_n491), .ZN(new_n529));
  XOR2_X1   g328(.A(G190gat), .B(G218gat), .Z(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT101), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n518), .A2(new_n525), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT100), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n511), .A2(new_n517), .B1(new_n521), .B2(new_n524), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n519), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n213), .A2(new_n224), .A3(new_n214), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n224), .B1(new_n213), .B2(new_n214), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n532), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n532), .B(new_n540), .C1(new_n526), .C2(new_n527), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n529), .B(new_n531), .C1(new_n541), .C2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n540), .B1(new_n526), .B2(new_n527), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT101), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n542), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n531), .B1(new_n548), .B2(new_n529), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n495), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n529), .B1(new_n541), .B2(new_n543), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n530), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(new_n494), .A3(new_n544), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G71gat), .A2(G78gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT90), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n555), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT90), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT91), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT91), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n558), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT92), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n565), .B1(new_n559), .B2(KEYINPUT9), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n555), .A2(KEYINPUT92), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G64gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(G57gat), .ZN(new_n570));
  INV_X1    g369(.A(G57gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(G64gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n566), .A2(new_n568), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n562), .A2(new_n564), .A3(new_n574), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n571), .A2(KEYINPUT93), .A3(KEYINPUT94), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT93), .ZN(new_n577));
  OAI21_X1  g376(.A(G64gat), .B1(new_n577), .B2(G57gat), .ZN(new_n578));
  OAI22_X1  g377(.A1(new_n576), .A2(new_n578), .B1(KEYINPUT94), .B2(new_n570), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n559), .A2(new_n556), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n579), .A2(new_n580), .A3(new_n568), .A4(new_n566), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n586));
  OR2_X1    g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G183gat), .B(G211gat), .Z(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n587), .A2(new_n592), .A3(new_n588), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT96), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n595), .B1(new_n575), .B2(new_n581), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n575), .A2(new_n581), .A3(new_n595), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(KEYINPUT21), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n223), .ZN(new_n600));
  XNOR2_X1  g399(.A(G127gat), .B(G155gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n601), .B(new_n602), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n599), .A2(new_n223), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n594), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n591), .A2(new_n604), .A3(new_n606), .A4(new_n593), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT102), .B1(new_n554), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT102), .ZN(new_n612));
  INV_X1    g411(.A(new_n610), .ZN(new_n613));
  AOI211_X1 g412(.A(new_n612), .B(new_n613), .C1(new_n550), .C2(new_n553), .ZN(new_n614));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT103), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n598), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n618), .A2(new_n596), .A3(new_n619), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n534), .A2(new_n620), .A3(new_n536), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n575), .A2(new_n581), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n515), .A2(new_n509), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(new_n525), .A3(new_n623), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n624), .B(new_n619), .C1(new_n622), .C2(new_n535), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n617), .B1(new_n621), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n624), .B1(new_n535), .B2(new_n622), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n616), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n627), .A2(new_n629), .A3(new_n633), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n611), .A2(new_n614), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n490), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n639), .A2(new_n389), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(new_n218), .ZN(G1324gat));
  INV_X1    g440(.A(new_n487), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n490), .A2(new_n642), .A3(new_n638), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT16), .B(G8gat), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT42), .ZN(new_n645));
  OR3_X1    g444(.A1(new_n643), .A2(KEYINPUT105), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT105), .B1(new_n643), .B2(new_n645), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n643), .A2(KEYINPUT104), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n643), .A2(KEYINPUT104), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n649), .A2(G8gat), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n644), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n649), .B2(new_n650), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n648), .B(new_n651), .C1(new_n653), .C2(KEYINPUT42), .ZN(G1325gat));
  OAI21_X1  g453(.A(G15gat), .B1(new_n639), .B2(new_n452), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n446), .A2(G15gat), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n655), .B1(new_n639), .B2(new_n656), .ZN(G1326gat));
  OR3_X1    g456(.A1(new_n639), .A2(KEYINPUT106), .A3(new_n411), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT106), .B1(new_n639), .B2(new_n411), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT43), .B(G22gat), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n660), .B1(new_n658), .B2(new_n659), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(G1327gat));
  AND3_X1   g462(.A1(new_n466), .A2(new_n467), .A3(new_n311), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n476), .A2(KEYINPUT38), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n488), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n453), .A2(new_n450), .A3(new_n449), .ZN(new_n667));
  OAI22_X1  g466(.A1(new_n666), .A2(new_n667), .B1(new_n445), .B2(new_n447), .ZN(new_n668));
  INV_X1    g467(.A(new_n554), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n668), .A2(KEYINPUT44), .A3(new_n669), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n252), .A2(new_n637), .A3(new_n610), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n672), .A2(new_n467), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(G29gat), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n554), .A2(new_n610), .A3(new_n637), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n389), .A2(G29gat), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n668), .A2(new_n251), .A3(new_n677), .A4(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n676), .A2(KEYINPUT108), .A3(new_n681), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(G1328gat));
  NOR2_X1   g485(.A1(new_n487), .A2(G36gat), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n668), .A2(new_n251), .A3(new_n677), .A4(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT46), .Z(new_n689));
  NAND4_X1  g488(.A1(new_n672), .A2(new_n642), .A3(new_n673), .A4(new_n674), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G36gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT109), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n689), .A2(new_n691), .A3(KEYINPUT109), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(G1329gat));
  AND2_X1   g495(.A1(new_n490), .A2(new_n677), .ZN(new_n697));
  INV_X1    g496(.A(new_n446), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(G43gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n672), .A2(new_n673), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n452), .A2(new_n700), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(new_n674), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT47), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n701), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(G1330gat));
  NAND4_X1  g508(.A1(new_n672), .A2(new_n412), .A3(new_n673), .A4(new_n674), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G50gat), .ZN(new_n711));
  INV_X1    g510(.A(G50gat), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n712), .A3(new_n412), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT48), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n711), .A2(new_n713), .A3(KEYINPUT48), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(G1331gat));
  NOR2_X1   g517(.A1(new_n611), .A2(new_n614), .ZN(new_n719));
  AND4_X1   g518(.A1(new_n668), .A2(new_n252), .A3(new_n719), .A4(new_n637), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n467), .ZN(new_n721));
  XOR2_X1   g520(.A(KEYINPUT93), .B(G57gat), .Z(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1332gat));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n642), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(KEYINPUT49), .B(G64gat), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n720), .A2(new_n642), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1333gat));
  NAND2_X1  g529(.A1(new_n720), .A2(new_n451), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n446), .A2(G71gat), .ZN(new_n732));
  AOI22_X1  g531(.A1(new_n731), .A2(G71gat), .B1(new_n720), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g533(.A1(new_n720), .A2(new_n412), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g535(.A1(new_n251), .A2(new_n610), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n637), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n702), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(G85gat), .B1(new_n741), .B2(new_n389), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n554), .B1(new_n448), .B2(new_n489), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT51), .B1(new_n743), .B2(new_n737), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n670), .A2(new_n745), .A3(new_n738), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n389), .A2(G85gat), .A3(new_n739), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n748), .B(KEYINPUT111), .Z(new_n749));
  OAI21_X1  g548(.A(new_n742), .B1(new_n747), .B2(new_n749), .ZN(G1336gat));
  NAND4_X1  g549(.A1(new_n672), .A2(new_n642), .A3(new_n673), .A4(new_n740), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G92gat), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n487), .A2(G92gat), .A3(new_n739), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n747), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT52), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n752), .B(new_n757), .C1(new_n747), .C2(new_n754), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(G1337gat));
  OAI21_X1  g558(.A(G99gat), .B1(new_n741), .B2(new_n452), .ZN(new_n760));
  OR3_X1    g559(.A1(new_n446), .A2(G99gat), .A3(new_n739), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n747), .B2(new_n761), .ZN(G1338gat));
  NAND4_X1  g561(.A1(new_n672), .A2(new_n412), .A3(new_n673), .A4(new_n740), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G106gat), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n411), .A2(G106gat), .A3(new_n739), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n744), .B2(new_n746), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n764), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT53), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n764), .A2(new_n766), .A3(new_n767), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(G1339gat));
  INV_X1    g571(.A(new_n239), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n226), .A2(new_n229), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(G229gat), .A3(G233gat), .ZN(new_n775));
  OR3_X1    g574(.A1(new_n232), .A2(new_n233), .A3(new_n231), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n773), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n245), .A2(new_n247), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n241), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n637), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT113), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n534), .A2(new_n620), .A3(new_n536), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n783), .A2(new_n625), .A3(new_n616), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n616), .B1(new_n783), .B2(new_n625), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n786), .B(new_n617), .C1(new_n621), .C2(new_n626), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n634), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n782), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n783), .A2(new_n625), .A3(new_n616), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n627), .A2(KEYINPUT54), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n633), .B1(new_n785), .B2(new_n786), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(KEYINPUT55), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n790), .A2(new_n251), .A3(new_n636), .A4(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n669), .B1(new_n781), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n636), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT55), .B1(new_n792), .B2(new_n793), .ZN(new_n798));
  INV_X1    g597(.A(new_n777), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n248), .A2(new_n799), .ZN(new_n800));
  OR4_X1    g599(.A1(new_n554), .A2(new_n797), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n613), .B1(new_n796), .B2(new_n802), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n545), .A2(new_n549), .A3(new_n495), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n494), .B1(new_n552), .B2(new_n544), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n610), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n612), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n554), .A2(KEYINPUT102), .A3(new_n610), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n807), .A2(new_n252), .A3(new_n808), .A4(new_n739), .ZN(new_n809));
  AOI211_X1 g608(.A(new_n412), .B(new_n446), .C1(new_n803), .C2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n810), .A2(new_n467), .A3(new_n487), .ZN(new_n811));
  OAI21_X1  g610(.A(G113gat), .B1(new_n811), .B2(new_n252), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n389), .B1(new_n803), .B2(new_n809), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n813), .A2(new_n444), .A3(new_n487), .ZN(new_n814));
  INV_X1    g613(.A(new_n347), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n815), .A3(new_n251), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n812), .A2(new_n816), .ZN(G1340gat));
  NOR3_X1   g616(.A1(new_n811), .A2(new_n340), .A3(new_n739), .ZN(new_n818));
  AOI21_X1  g617(.A(G120gat), .B1(new_n814), .B2(new_n637), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(G1341gat));
  OAI21_X1  g619(.A(G127gat), .B1(new_n811), .B2(new_n613), .ZN(new_n821));
  INV_X1    g620(.A(G127gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n814), .A2(new_n822), .A3(new_n610), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(G1342gat));
  INV_X1    g623(.A(G134gat), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n814), .A2(new_n825), .A3(new_n669), .ZN(new_n826));
  XNOR2_X1  g625(.A(KEYINPUT114), .B(KEYINPUT56), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  OAI21_X1  g628(.A(G134gat), .B1(new_n811), .B2(new_n554), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(G1343gat));
  NOR3_X1   g630(.A1(new_n451), .A2(new_n411), .A3(new_n642), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n813), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n323), .B1(new_n833), .B2(new_n252), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n803), .A2(new_n809), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n412), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n836), .A2(KEYINPUT115), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n795), .A2(new_n780), .A3(KEYINPUT116), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n554), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT116), .B1(new_n795), .B2(new_n780), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n801), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n613), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n809), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n411), .A2(new_n837), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n411), .B1(new_n803), .B2(new_n809), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n848), .B2(KEYINPUT57), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n838), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n451), .A2(new_n389), .A3(new_n642), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n251), .A2(G141gat), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n834), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT58), .Z(G1344gat));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n850), .A2(new_n637), .A3(new_n851), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n320), .A2(KEYINPUT59), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n719), .A2(new_n862), .A3(new_n252), .A4(new_n739), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n809), .A2(KEYINPUT117), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n795), .A2(new_n780), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n554), .A3(new_n839), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n610), .B1(new_n869), .B2(new_n801), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n861), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n843), .A2(KEYINPUT118), .A3(new_n864), .A4(new_n863), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n412), .A3(new_n872), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n873), .A2(KEYINPUT119), .A3(new_n837), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT119), .B1(new_n873), .B2(new_n837), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n835), .A2(new_n845), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n851), .A2(new_n637), .ZN(new_n879));
  OAI21_X1  g678(.A(G148gat), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n860), .B1(new_n880), .B2(KEYINPUT59), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n833), .A2(G148gat), .A3(new_n739), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n857), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n882), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n873), .A2(new_n837), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n873), .A2(KEYINPUT119), .A3(new_n837), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n889), .A3(new_n876), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n637), .A3(new_n851), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n885), .B1(new_n891), .B2(G148gat), .ZN(new_n892));
  OAI211_X1 g691(.A(KEYINPUT120), .B(new_n884), .C1(new_n892), .C2(new_n860), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n883), .A2(new_n893), .ZN(G1345gat));
  OAI21_X1  g693(.A(G155gat), .B1(new_n853), .B2(new_n613), .ZN(new_n895));
  INV_X1    g694(.A(new_n833), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n326), .A3(new_n610), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(G1346gat));
  AOI21_X1  g697(.A(G162gat), .B1(new_n896), .B2(new_n669), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n554), .A2(new_n327), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n852), .B2(new_n900), .ZN(G1347gat));
  NOR2_X1   g700(.A1(new_n487), .A2(new_n467), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n810), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(G169gat), .B1(new_n903), .B2(new_n252), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT122), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n835), .A2(new_n389), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT121), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n444), .A2(new_n642), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n264), .A3(new_n251), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n905), .A2(new_n910), .ZN(G1348gat));
  NAND3_X1  g710(.A1(new_n909), .A2(new_n265), .A3(new_n637), .ZN(new_n912));
  OAI21_X1  g711(.A(G176gat), .B1(new_n903), .B2(new_n739), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1349gat));
  NOR2_X1   g713(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n909), .A2(new_n277), .A3(new_n610), .ZN(new_n916));
  OAI21_X1  g715(.A(G183gat), .B1(new_n903), .B2(new_n613), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g717(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n918), .B(new_n919), .ZN(G1350gat));
  OAI21_X1  g719(.A(G190gat), .B1(new_n903), .B2(new_n554), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT61), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n909), .A2(new_n278), .A3(new_n669), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1351gat));
  NOR3_X1   g723(.A1(new_n451), .A2(new_n411), .A3(new_n487), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT124), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n926), .A2(new_n907), .ZN(new_n927));
  AOI21_X1  g726(.A(G197gat), .B1(new_n927), .B2(new_n251), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n890), .A2(KEYINPUT125), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n888), .A2(new_n930), .A3(new_n889), .A4(new_n876), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n452), .A2(new_n902), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n934), .A2(G197gat), .A3(new_n251), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n928), .B1(new_n932), .B2(new_n935), .ZN(G1352gat));
  NOR2_X1   g735(.A1(new_n739), .A2(G204gat), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n927), .A2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n938), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n934), .A2(new_n637), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n941), .B1(new_n929), .B2(new_n931), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(G204gat), .B1(new_n942), .B2(new_n943), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n940), .B1(new_n944), .B2(new_n945), .ZN(G1353gat));
  NOR3_X1   g745(.A1(new_n878), .A2(new_n613), .A3(new_n933), .ZN(new_n947));
  OR3_X1    g746(.A1(new_n947), .A2(KEYINPUT63), .A3(new_n291), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n613), .A2(G211gat), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n927), .A2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n927), .A2(KEYINPUT127), .A3(new_n949), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(KEYINPUT63), .B1(new_n947), .B2(new_n291), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n948), .A2(new_n954), .A3(new_n955), .ZN(G1354gat));
  AOI21_X1  g755(.A(G218gat), .B1(new_n927), .B2(new_n669), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n933), .A2(new_n292), .A3(new_n554), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n932), .B2(new_n958), .ZN(G1355gat));
endmodule


