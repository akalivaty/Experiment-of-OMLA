

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770;

  XNOR2_X1 U377 ( .A(n555), .B(n374), .ZN(n586) );
  BUF_X1 U378 ( .A(n608), .Z(n570) );
  XNOR2_X1 U379 ( .A(n428), .B(n393), .ZN(n757) );
  NAND2_X1 U380 ( .A1(n354), .A2(n591), .ZN(n593) );
  NAND2_X1 U381 ( .A1(n587), .A2(n588), .ZN(n354) );
  XNOR2_X1 U382 ( .A(G119), .B(G128), .ZN(n462) );
  INV_X1 U383 ( .A(G953), .ZN(n762) );
  XOR2_X1 U384 ( .A(KEYINPUT103), .B(n528), .Z(n355) );
  INV_X1 U385 ( .A(n561), .ZN(n515) );
  OR2_X1 U386 ( .A1(n770), .A2(n629), .ZN(n630) );
  INV_X1 U387 ( .A(KEYINPUT46), .ZN(n373) );
  XNOR2_X1 U388 ( .A(n378), .B(KEYINPUT64), .ZN(n643) );
  XNOR2_X1 U389 ( .A(n371), .B(n370), .ZN(n640) );
  NAND2_X1 U390 ( .A1(n631), .A2(n372), .ZN(n371) );
  AND2_X1 U391 ( .A1(n584), .A2(n583), .ZN(n594) );
  XNOR2_X1 U392 ( .A(n630), .B(n373), .ZN(n372) );
  XNOR2_X1 U393 ( .A(n400), .B(n362), .ZN(n629) );
  NAND2_X1 U394 ( .A1(n571), .A2(n515), .ZN(n548) );
  AND2_X1 U395 ( .A1(n547), .A2(n702), .ZN(n571) );
  XNOR2_X1 U396 ( .A(n509), .B(G469), .ZN(n513) );
  OR2_X1 U397 ( .A1(n696), .A2(n610), .ZN(n514) );
  OR2_X1 U398 ( .A1(n738), .A2(G902), .ZN(n472) );
  XNOR2_X1 U399 ( .A(n442), .B(n416), .ZN(n758) );
  INV_X1 U400 ( .A(KEYINPUT4), .ZN(n393) );
  XNOR2_X1 U401 ( .A(n757), .B(G101), .ZN(n487) );
  XNOR2_X1 U402 ( .A(n491), .B(n490), .ZN(n503) );
  XNOR2_X1 U403 ( .A(G137), .B(G134), .ZN(n490) );
  NAND2_X1 U404 ( .A1(n586), .A2(n589), .ZN(n556) );
  AND2_X1 U405 ( .A1(n664), .A2(n672), .ZN(n568) );
  XOR2_X1 U406 ( .A(G146), .B(KEYINPUT5), .Z(n486) );
  INV_X1 U407 ( .A(n503), .ZN(n364) );
  XNOR2_X1 U408 ( .A(G146), .B(G125), .ZN(n442) );
  INV_X1 U409 ( .A(KEYINPUT70), .ZN(n624) );
  NAND2_X1 U410 ( .A1(G234), .A2(G237), .ZN(n477) );
  INV_X1 U411 ( .A(n610), .ZN(n367) );
  XNOR2_X1 U412 ( .A(n609), .B(n369), .ZN(n368) );
  INV_X1 U413 ( .A(KEYINPUT30), .ZN(n369) );
  XNOR2_X1 U414 ( .A(n408), .B(G478), .ZN(n551) );
  OR2_X1 U415 ( .A1(n732), .A2(G902), .ZN(n408) );
  AND2_X1 U416 ( .A1(n380), .A2(n360), .ZN(n379) );
  NAND2_X1 U417 ( .A1(n635), .A2(n395), .ZN(n380) );
  NAND2_X1 U418 ( .A1(n398), .A2(KEYINPUT2), .ZN(n395) );
  INV_X1 U419 ( .A(KEYINPUT9), .ZN(n394) );
  XNOR2_X1 U420 ( .A(n744), .B(n376), .ZN(n375) );
  XNOR2_X1 U421 ( .A(KEYINPUT73), .B(KEYINPUT72), .ZN(n376) );
  XNOR2_X1 U422 ( .A(n539), .B(n538), .ZN(n725) );
  XNOR2_X1 U423 ( .A(n628), .B(n627), .ZN(n632) );
  BUF_X1 U424 ( .A(n547), .Z(n703) );
  XNOR2_X1 U425 ( .A(n533), .B(n386), .ZN(n385) );
  INV_X1 U426 ( .A(KEYINPUT22), .ZN(n386) );
  BUF_X1 U427 ( .A(n513), .Z(n611) );
  XOR2_X1 U428 ( .A(G146), .B(G104), .Z(n498) );
  XNOR2_X1 U429 ( .A(n405), .B(n404), .ZN(n598) );
  INV_X1 U430 ( .A(KEYINPUT89), .ZN(n404) );
  INV_X1 U431 ( .A(n634), .ZN(n398) );
  NAND2_X1 U432 ( .A1(n397), .A2(n398), .ZN(n396) );
  INV_X1 U433 ( .A(n633), .ZN(n397) );
  XNOR2_X1 U434 ( .A(n407), .B(G122), .ZN(n430) );
  INV_X1 U435 ( .A(G107), .ZN(n407) );
  XNOR2_X1 U436 ( .A(G116), .B(G134), .ZN(n429) );
  XOR2_X1 U437 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n425) );
  XNOR2_X1 U438 ( .A(G140), .B(KEYINPUT12), .ZN(n410) );
  NAND2_X1 U439 ( .A1(n579), .A2(n681), .ZN(n405) );
  XNOR2_X1 U440 ( .A(n365), .B(n363), .ZN(n666) );
  XNOR2_X1 U441 ( .A(n364), .B(n488), .ZN(n363) );
  XNOR2_X1 U442 ( .A(n377), .B(G107), .ZN(n744) );
  INV_X1 U443 ( .A(G110), .ZN(n377) );
  XNOR2_X1 U444 ( .A(KEYINPUT69), .B(G140), .ZN(n502) );
  XNOR2_X1 U445 ( .A(G122), .B(G104), .ZN(n439) );
  XNOR2_X1 U446 ( .A(G113), .B(G143), .ZN(n418) );
  XOR2_X1 U447 ( .A(G131), .B(KEYINPUT68), .Z(n491) );
  INV_X1 U448 ( .A(KEYINPUT48), .ZN(n370) );
  OR2_X1 U449 ( .A1(n635), .A2(n633), .ZN(n761) );
  NOR2_X1 U450 ( .A1(n612), .A2(n366), .ZN(n626) );
  NAND2_X1 U451 ( .A1(n389), .A2(n388), .ZN(n387) );
  NOR2_X1 U452 ( .A1(n454), .A2(n455), .ZN(n388) );
  INV_X1 U453 ( .A(n540), .ZN(n599) );
  XNOR2_X1 U454 ( .A(n570), .B(KEYINPUT6), .ZN(n561) );
  INV_X1 U455 ( .A(n703), .ZN(n384) );
  NAND2_X1 U456 ( .A1(n381), .A2(n379), .ZN(n378) );
  NAND2_X1 U457 ( .A1(n688), .A2(n399), .ZN(n381) );
  XNOR2_X1 U458 ( .A(n409), .B(n435), .ZN(n732) );
  XNOR2_X1 U459 ( .A(n433), .B(n434), .ZN(n409) );
  XNOR2_X1 U460 ( .A(n743), .B(n446), .ZN(n447) );
  AND2_X1 U461 ( .A1(n648), .A2(G953), .ZN(n742) );
  NOR2_X1 U462 ( .A1(n719), .A2(n383), .ZN(n720) );
  INV_X1 U463 ( .A(n725), .ZN(n382) );
  NOR2_X1 U464 ( .A1(n725), .A2(n540), .ZN(n400) );
  XNOR2_X1 U465 ( .A(n401), .B(n361), .ZN(n770) );
  NOR2_X1 U466 ( .A1(n632), .A2(n681), .ZN(n401) );
  INV_X1 U467 ( .A(KEYINPUT35), .ZN(n374) );
  XNOR2_X1 U468 ( .A(n567), .B(n566), .ZN(n672) );
  AND2_X1 U469 ( .A1(n712), .A2(n405), .ZN(n356) );
  XNOR2_X1 U470 ( .A(n513), .B(KEYINPUT1), .ZN(n547) );
  AND2_X1 U471 ( .A1(n391), .A2(n390), .ZN(n357) );
  XNOR2_X1 U472 ( .A(n487), .B(n375), .ZN(n501) );
  XOR2_X1 U473 ( .A(n565), .B(n564), .Z(n358) );
  NAND2_X1 U474 ( .A1(n385), .A2(n384), .ZN(n558) );
  AND2_X1 U475 ( .A1(n696), .A2(n367), .ZN(n359) );
  NAND2_X1 U476 ( .A1(n396), .A2(n395), .ZN(n360) );
  AND2_X1 U477 ( .A1(n715), .A2(n714), .ZN(n712) );
  XOR2_X1 U478 ( .A(KEYINPUT109), .B(KEYINPUT40), .Z(n361) );
  XOR2_X1 U479 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n362) );
  XNOR2_X1 U480 ( .A(n447), .B(n501), .ZN(n658) );
  XNOR2_X1 U481 ( .A(n489), .B(n440), .ZN(n743) );
  INV_X1 U482 ( .A(KEYINPUT2), .ZN(n399) );
  NAND2_X1 U483 ( .A1(n672), .A2(n664), .ZN(n585) );
  XNOR2_X1 U484 ( .A(n487), .B(n489), .ZN(n365) );
  XNOR2_X2 U485 ( .A(n406), .B(n437), .ZN(n489) );
  NAND2_X1 U486 ( .A1(n368), .A2(n359), .ZN(n366) );
  INV_X1 U487 ( .A(n640), .ZN(n635) );
  XNOR2_X1 U488 ( .A(n586), .B(G122), .ZN(G24) );
  XNOR2_X2 U489 ( .A(G143), .B(G128), .ZN(n428) );
  XNOR2_X2 U490 ( .A(n596), .B(n595), .ZN(n688) );
  NAND2_X1 U491 ( .A1(n382), .A2(n403), .ZN(n726) );
  INV_X1 U492 ( .A(n403), .ZN(n383) );
  XNOR2_X2 U493 ( .A(n548), .B(KEYINPUT33), .ZN(n403) );
  NAND2_X1 U494 ( .A1(n385), .A2(n358), .ZN(n567) );
  NAND2_X1 U495 ( .A1(n389), .A2(n714), .ZN(n392) );
  NAND2_X2 U496 ( .A1(n357), .A2(n387), .ZN(n597) );
  INV_X1 U497 ( .A(n536), .ZN(n389) );
  NAND2_X1 U498 ( .A1(n454), .A2(n455), .ZN(n390) );
  NAND2_X1 U499 ( .A1(n536), .A2(n455), .ZN(n391) );
  NOR2_X1 U500 ( .A1(n619), .A2(n392), .ZN(n620) );
  OR2_X2 U501 ( .A1(n688), .A2(n641), .ZN(n642) );
  XNOR2_X1 U502 ( .A(n625), .B(n624), .ZN(n631) );
  NAND2_X1 U503 ( .A1(n594), .A2(n593), .ZN(n596) );
  XNOR2_X2 U504 ( .A(n642), .B(KEYINPUT77), .ZN(n693) );
  XNOR2_X1 U505 ( .A(n428), .B(n394), .ZN(n432) );
  INV_X1 U506 ( .A(n532), .ZN(n577) );
  NAND2_X1 U507 ( .A1(n403), .A2(n532), .ZN(n550) );
  XNOR2_X2 U508 ( .A(n527), .B(n402), .ZN(n532) );
  INV_X1 U509 ( .A(KEYINPUT0), .ZN(n402) );
  XNOR2_X2 U510 ( .A(n436), .B(n438), .ZN(n406) );
  XNOR2_X1 U511 ( .A(n542), .B(KEYINPUT105), .ZN(n579) );
  XOR2_X1 U512 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n411) );
  XNOR2_X1 U513 ( .A(n411), .B(n410), .ZN(n414) );
  NOR2_X2 U514 ( .A1(G953), .A2(G237), .ZN(n484) );
  NAND2_X1 U515 ( .A1(G214), .A2(n484), .ZN(n412) );
  XNOR2_X1 U516 ( .A(n412), .B(KEYINPUT11), .ZN(n413) );
  XNOR2_X1 U517 ( .A(n414), .B(n413), .ZN(n417) );
  INV_X1 U518 ( .A(KEYINPUT67), .ZN(n415) );
  XNOR2_X1 U519 ( .A(n415), .B(KEYINPUT10), .ZN(n416) );
  XNOR2_X1 U520 ( .A(n417), .B(n758), .ZN(n421) );
  XNOR2_X1 U521 ( .A(n418), .B(n439), .ZN(n419) );
  XNOR2_X1 U522 ( .A(n491), .B(n419), .ZN(n420) );
  XNOR2_X1 U523 ( .A(n421), .B(n420), .ZN(n644) );
  NOR2_X2 U524 ( .A1(n644), .A2(G902), .ZN(n423) );
  XNOR2_X1 U525 ( .A(KEYINPUT13), .B(G475), .ZN(n422) );
  XNOR2_X2 U526 ( .A(n423), .B(n422), .ZN(n528) );
  NAND2_X1 U527 ( .A1(G234), .A2(n762), .ZN(n424) );
  XNOR2_X1 U528 ( .A(n425), .B(n424), .ZN(n427) );
  INV_X1 U529 ( .A(KEYINPUT91), .ZN(n426) );
  XNOR2_X1 U530 ( .A(n427), .B(n426), .ZN(n457) );
  NAND2_X1 U531 ( .A1(n457), .A2(G217), .ZN(n435) );
  XNOR2_X1 U532 ( .A(KEYINPUT104), .B(KEYINPUT7), .ZN(n434) );
  XNOR2_X1 U533 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U534 ( .A(n432), .B(n431), .ZN(n433) );
  INV_X1 U535 ( .A(n551), .ZN(n541) );
  NAND2_X1 U536 ( .A1(n355), .A2(n541), .ZN(n681) );
  INV_X1 U537 ( .A(n681), .ZN(n456) );
  XNOR2_X1 U538 ( .A(G119), .B(G116), .ZN(n437) );
  XNOR2_X2 U539 ( .A(G113), .B(KEYINPUT71), .ZN(n436) );
  XNOR2_X2 U540 ( .A(KEYINPUT94), .B(KEYINPUT3), .ZN(n438) );
  XNOR2_X1 U541 ( .A(n439), .B(KEYINPUT16), .ZN(n440) );
  XNOR2_X1 U542 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n441) );
  XNOR2_X1 U543 ( .A(n442), .B(n441), .ZN(n445) );
  NAND2_X1 U544 ( .A1(n762), .A2(G224), .ZN(n443) );
  XNOR2_X1 U545 ( .A(n443), .B(KEYINPUT95), .ZN(n444) );
  XNOR2_X1 U546 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U547 ( .A(G902), .B(KEYINPUT15), .ZN(n634) );
  NAND2_X1 U548 ( .A1(n658), .A2(n634), .ZN(n451) );
  NOR2_X1 U549 ( .A1(G237), .A2(G902), .ZN(n448) );
  XNOR2_X1 U550 ( .A(n448), .B(KEYINPUT76), .ZN(n453) );
  INV_X1 U551 ( .A(G210), .ZN(n449) );
  OR2_X1 U552 ( .A1(n453), .A2(n449), .ZN(n450) );
  XNOR2_X2 U553 ( .A(n451), .B(n450), .ZN(n536) );
  INV_X1 U554 ( .A(G214), .ZN(n452) );
  OR2_X1 U555 ( .A1(n453), .A2(n452), .ZN(n714) );
  INV_X1 U556 ( .A(n714), .ZN(n454) );
  XNOR2_X1 U557 ( .A(KEYINPUT78), .B(KEYINPUT19), .ZN(n455) );
  AND2_X1 U558 ( .A1(n456), .A2(n597), .ZN(n511) );
  NAND2_X1 U559 ( .A1(n457), .A2(G221), .ZN(n467) );
  XNOR2_X1 U560 ( .A(G110), .B(KEYINPUT79), .ZN(n459) );
  XNOR2_X1 U561 ( .A(KEYINPUT98), .B(KEYINPUT23), .ZN(n458) );
  XNOR2_X1 U562 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U563 ( .A(n758), .B(n460), .ZN(n465) );
  XNOR2_X1 U564 ( .A(KEYINPUT24), .B(G137), .ZN(n461) );
  XNOR2_X1 U565 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U566 ( .A(n463), .B(n502), .ZN(n464) );
  XNOR2_X1 U567 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U568 ( .A(n467), .B(n466), .ZN(n738) );
  XOR2_X1 U569 ( .A(KEYINPUT20), .B(KEYINPUT99), .Z(n469) );
  NAND2_X1 U570 ( .A1(n634), .A2(G234), .ZN(n468) );
  XNOR2_X1 U571 ( .A(n469), .B(n468), .ZN(n473) );
  AND2_X1 U572 ( .A1(n473), .A2(G217), .ZN(n470) );
  XNOR2_X1 U573 ( .A(n470), .B(KEYINPUT25), .ZN(n471) );
  XNOR2_X2 U574 ( .A(n472), .B(n471), .ZN(n696) );
  NAND2_X1 U575 ( .A1(n473), .A2(G221), .ZN(n474) );
  XNOR2_X1 U576 ( .A(n474), .B(KEYINPUT100), .ZN(n476) );
  INV_X1 U577 ( .A(KEYINPUT21), .ZN(n475) );
  XNOR2_X1 U578 ( .A(n476), .B(n475), .ZN(n695) );
  XNOR2_X1 U579 ( .A(n477), .B(KEYINPUT14), .ZN(n480) );
  NAND2_X1 U580 ( .A1(n480), .A2(G902), .ZN(n478) );
  XOR2_X1 U581 ( .A(n478), .B(KEYINPUT97), .Z(n520) );
  OR2_X1 U582 ( .A1(n520), .A2(n762), .ZN(n479) );
  NOR2_X1 U583 ( .A1(G900), .A2(n479), .ZN(n482) );
  NAND2_X1 U584 ( .A1(G952), .A2(n480), .ZN(n724) );
  OR2_X1 U585 ( .A1(n724), .A2(G953), .ZN(n524) );
  INV_X1 U586 ( .A(n524), .ZN(n481) );
  OR2_X1 U587 ( .A1(n482), .A2(n481), .ZN(n483) );
  NAND2_X1 U588 ( .A1(n695), .A2(n483), .ZN(n610) );
  INV_X1 U589 ( .A(n514), .ZN(n494) );
  NAND2_X1 U590 ( .A1(n484), .A2(G210), .ZN(n485) );
  XNOR2_X1 U591 ( .A(n486), .B(n485), .ZN(n488) );
  INV_X1 U592 ( .A(G902), .ZN(n508) );
  NAND2_X1 U593 ( .A1(n666), .A2(n508), .ZN(n493) );
  XNOR2_X1 U594 ( .A(G472), .B(KEYINPUT74), .ZN(n492) );
  XNOR2_X1 U595 ( .A(n493), .B(n492), .ZN(n608) );
  NAND2_X1 U596 ( .A1(n494), .A2(n570), .ZN(n496) );
  INV_X1 U597 ( .A(KEYINPUT28), .ZN(n495) );
  XNOR2_X1 U598 ( .A(n496), .B(n495), .ZN(n510) );
  NAND2_X1 U599 ( .A1(G227), .A2(n762), .ZN(n497) );
  XNOR2_X1 U600 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U601 ( .A(n499), .B(KEYINPUT81), .Z(n500) );
  XNOR2_X1 U602 ( .A(n501), .B(n500), .ZN(n504) );
  XNOR2_X1 U603 ( .A(n503), .B(n502), .ZN(n760) );
  XNOR2_X1 U604 ( .A(n760), .B(KEYINPUT80), .ZN(n505) );
  OR2_X1 U605 ( .A1(n504), .A2(n505), .ZN(n507) );
  NAND2_X1 U606 ( .A1(n505), .A2(n504), .ZN(n506) );
  NAND2_X1 U607 ( .A1(n507), .A2(n506), .ZN(n652) );
  NAND2_X1 U608 ( .A1(n652), .A2(n508), .ZN(n509) );
  NAND2_X1 U609 ( .A1(n510), .A2(n611), .ZN(n540) );
  NAND2_X1 U610 ( .A1(n511), .A2(n599), .ZN(n603) );
  XNOR2_X1 U611 ( .A(n603), .B(G146), .ZN(G48) );
  BUF_X1 U612 ( .A(n536), .Z(n512) );
  NOR2_X1 U613 ( .A1(n681), .A2(n514), .ZN(n516) );
  NAND2_X1 U614 ( .A1(n516), .A2(n515), .ZN(n619) );
  NOR2_X1 U615 ( .A1(n703), .A2(n619), .ZN(n517) );
  NAND2_X1 U616 ( .A1(n714), .A2(n517), .ZN(n518) );
  XNOR2_X1 U617 ( .A(n518), .B(KEYINPUT43), .ZN(n519) );
  NAND2_X1 U618 ( .A1(n512), .A2(n519), .ZN(n637) );
  XNOR2_X1 U619 ( .A(n637), .B(G140), .ZN(G42) );
  INV_X1 U620 ( .A(n520), .ZN(n523) );
  NOR2_X1 U621 ( .A1(G898), .A2(n762), .ZN(n521) );
  XOR2_X1 U622 ( .A(KEYINPUT96), .B(n521), .Z(n746) );
  INV_X1 U623 ( .A(n746), .ZN(n522) );
  NAND2_X1 U624 ( .A1(n523), .A2(n522), .ZN(n525) );
  NAND2_X1 U625 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U626 ( .A1(n597), .A2(n526), .ZN(n527) );
  NOR2_X1 U627 ( .A1(n551), .A2(n528), .ZN(n529) );
  XNOR2_X1 U628 ( .A(n529), .B(KEYINPUT106), .ZN(n713) );
  NAND2_X1 U629 ( .A1(n713), .A2(n695), .ZN(n530) );
  XNOR2_X1 U630 ( .A(n530), .B(KEYINPUT107), .ZN(n531) );
  NAND2_X1 U631 ( .A1(n532), .A2(n531), .ZN(n533) );
  INV_X1 U632 ( .A(n558), .ZN(n535) );
  AND2_X1 U633 ( .A1(n561), .A2(n696), .ZN(n534) );
  NAND2_X1 U634 ( .A1(n535), .A2(n534), .ZN(n582) );
  XNOR2_X1 U635 ( .A(n582), .B(G101), .ZN(G3) );
  XNOR2_X1 U636 ( .A(n536), .B(KEYINPUT38), .ZN(n715) );
  NAND2_X1 U637 ( .A1(n713), .A2(n712), .ZN(n539) );
  INV_X1 U638 ( .A(KEYINPUT110), .ZN(n537) );
  XNOR2_X1 U639 ( .A(n537), .B(KEYINPUT41), .ZN(n538) );
  XOR2_X1 U640 ( .A(G137), .B(n629), .Z(G39) );
  NOR2_X2 U641 ( .A1(n355), .A2(n541), .ZN(n542) );
  BUF_X1 U642 ( .A(n579), .Z(n543) );
  INV_X1 U643 ( .A(n597), .ZN(n544) );
  NOR2_X1 U644 ( .A1(n543), .A2(n544), .ZN(n545) );
  NAND2_X1 U645 ( .A1(n545), .A2(n599), .ZN(n604) );
  XOR2_X1 U646 ( .A(G128), .B(KEYINPUT29), .Z(n546) );
  XNOR2_X1 U647 ( .A(n604), .B(n546), .ZN(G30) );
  AND2_X1 U648 ( .A1(n696), .A2(n695), .ZN(n702) );
  XNOR2_X1 U649 ( .A(KEYINPUT83), .B(KEYINPUT34), .ZN(n549) );
  XNOR2_X1 U650 ( .A(n550), .B(n549), .ZN(n554) );
  NAND2_X1 U651 ( .A1(n551), .A2(n528), .ZN(n613) );
  INV_X1 U652 ( .A(KEYINPUT82), .ZN(n552) );
  XNOR2_X1 U653 ( .A(n613), .B(n552), .ZN(n553) );
  NAND2_X1 U654 ( .A1(n554), .A2(n553), .ZN(n555) );
  INV_X1 U655 ( .A(KEYINPUT65), .ZN(n590) );
  NAND2_X1 U656 ( .A1(n556), .A2(n590), .ZN(n569) );
  INV_X1 U657 ( .A(KEYINPUT108), .ZN(n557) );
  XNOR2_X1 U658 ( .A(n558), .B(n557), .ZN(n560) );
  NOR2_X1 U659 ( .A1(n570), .A2(n696), .ZN(n559) );
  NAND2_X1 U660 ( .A1(n560), .A2(n559), .ZN(n664) );
  XNOR2_X1 U661 ( .A(n561), .B(KEYINPUT86), .ZN(n562) );
  INV_X1 U662 ( .A(n696), .ZN(n574) );
  AND2_X1 U663 ( .A1(n562), .A2(n574), .ZN(n563) );
  NAND2_X1 U664 ( .A1(n563), .A2(n703), .ZN(n565) );
  INV_X1 U665 ( .A(KEYINPUT85), .ZN(n564) );
  XNOR2_X1 U666 ( .A(KEYINPUT84), .B(KEYINPUT32), .ZN(n566) );
  NAND2_X1 U667 ( .A1(n569), .A2(n568), .ZN(n584) );
  NAND2_X1 U668 ( .A1(n571), .A2(n570), .ZN(n709) );
  OR2_X1 U669 ( .A1(n577), .A2(n709), .ZN(n573) );
  INV_X1 U670 ( .A(KEYINPUT31), .ZN(n572) );
  XNOR2_X1 U671 ( .A(n573), .B(n572), .ZN(n683) );
  NOR2_X1 U672 ( .A1(n574), .A2(n570), .ZN(n575) );
  NAND2_X1 U673 ( .A1(n611), .A2(n575), .ZN(n576) );
  NOR2_X1 U674 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U675 ( .A1(n695), .A2(n578), .ZN(n675) );
  NAND2_X1 U676 ( .A1(n683), .A2(n675), .ZN(n580) );
  NAND2_X1 U677 ( .A1(n580), .A2(n598), .ZN(n581) );
  AND2_X1 U678 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U679 ( .A1(n585), .A2(n590), .ZN(n588) );
  AND2_X1 U680 ( .A1(n586), .A2(KEYINPUT44), .ZN(n587) );
  INV_X1 U681 ( .A(KEYINPUT44), .ZN(n589) );
  NAND2_X1 U682 ( .A1(n590), .A2(n589), .ZN(n591) );
  INV_X1 U683 ( .A(KEYINPUT45), .ZN(n595) );
  AND2_X1 U684 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U685 ( .A1(n600), .A2(n599), .ZN(n602) );
  INV_X1 U686 ( .A(KEYINPUT47), .ZN(n601) );
  NAND2_X1 U687 ( .A1(n602), .A2(n601), .ZN(n607) );
  NAND2_X1 U688 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U689 ( .A1(n605), .A2(KEYINPUT47), .ZN(n606) );
  NAND2_X1 U690 ( .A1(n607), .A2(n606), .ZN(n617) );
  NAND2_X1 U691 ( .A1(n714), .A2(n608), .ZN(n609) );
  INV_X1 U692 ( .A(n611), .ZN(n612) );
  NOR2_X1 U693 ( .A1(n613), .A2(n512), .ZN(n614) );
  AND2_X1 U694 ( .A1(n626), .A2(n614), .ZN(n679) );
  INV_X1 U695 ( .A(KEYINPUT90), .ZN(n615) );
  XNOR2_X1 U696 ( .A(n679), .B(n615), .ZN(n616) );
  NAND2_X1 U697 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U698 ( .A(n618), .B(KEYINPUT75), .ZN(n623) );
  XNOR2_X1 U699 ( .A(n620), .B(KEYINPUT36), .ZN(n621) );
  AND2_X1 U700 ( .A1(n621), .A2(n703), .ZN(n685) );
  INV_X1 U701 ( .A(n685), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n715), .ZN(n628) );
  INV_X1 U704 ( .A(KEYINPUT39), .ZN(n627) );
  OR2_X1 U705 ( .A1(n632), .A2(n543), .ZN(n687) );
  NAND2_X1 U706 ( .A1(n687), .A2(n637), .ZN(n633) );
  NAND2_X1 U707 ( .A1(n687), .A2(KEYINPUT2), .ZN(n636) );
  XNOR2_X1 U708 ( .A(n636), .B(KEYINPUT87), .ZN(n638) );
  AND2_X1 U709 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X4 U711 ( .A1(n643), .A2(n693), .ZN(n737) );
  NAND2_X1 U712 ( .A1(n737), .A2(G475), .ZN(n647) );
  XOR2_X1 U713 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n645) );
  XNOR2_X1 U714 ( .A(n644), .B(n645), .ZN(n646) );
  XNOR2_X1 U715 ( .A(n647), .B(n646), .ZN(n649) );
  INV_X1 U716 ( .A(G952), .ZN(n648) );
  NOR2_X2 U717 ( .A1(n649), .A2(n742), .ZN(n650) );
  XNOR2_X1 U718 ( .A(n650), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U719 ( .A1(n737), .A2(G469), .ZN(n654) );
  XNOR2_X1 U720 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n651) );
  XNOR2_X1 U721 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X2 U723 ( .A1(n655), .A2(n742), .ZN(n657) );
  INV_X1 U724 ( .A(KEYINPUT119), .ZN(n656) );
  XNOR2_X1 U725 ( .A(n657), .B(n656), .ZN(G54) );
  NAND2_X1 U726 ( .A1(n737), .A2(G210), .ZN(n661) );
  XNOR2_X1 U727 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n659) );
  XNOR2_X1 U728 ( .A(n658), .B(n659), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n661), .B(n660), .ZN(n662) );
  NOR2_X2 U730 ( .A1(n662), .A2(n742), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n663), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U732 ( .A(n664), .B(G110), .ZN(G12) );
  NAND2_X1 U733 ( .A1(n737), .A2(G472), .ZN(n668) );
  XOR2_X1 U734 ( .A(KEYINPUT112), .B(KEYINPUT62), .Z(n665) );
  XNOR2_X1 U735 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U736 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X2 U737 ( .A1(n669), .A2(n742), .ZN(n671) );
  XNOR2_X1 U738 ( .A(KEYINPUT93), .B(KEYINPUT63), .ZN(n670) );
  XNOR2_X1 U739 ( .A(n671), .B(n670), .ZN(G57) );
  XNOR2_X1 U740 ( .A(n672), .B(G119), .ZN(G21) );
  NOR2_X1 U741 ( .A1(n681), .A2(n675), .ZN(n674) );
  XNOR2_X1 U742 ( .A(G104), .B(KEYINPUT113), .ZN(n673) );
  XNOR2_X1 U743 ( .A(n674), .B(n673), .ZN(G6) );
  NOR2_X1 U744 ( .A1(n543), .A2(n675), .ZN(n677) );
  XNOR2_X1 U745 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n676) );
  XNOR2_X1 U746 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U747 ( .A(G107), .B(n678), .ZN(G9) );
  XOR2_X1 U748 ( .A(G143), .B(n679), .Z(n680) );
  XNOR2_X1 U749 ( .A(KEYINPUT114), .B(n680), .ZN(G45) );
  NOR2_X1 U750 ( .A1(n681), .A2(n683), .ZN(n682) );
  XOR2_X1 U751 ( .A(G113), .B(n682), .Z(G15) );
  NOR2_X1 U752 ( .A1(n543), .A2(n683), .ZN(n684) );
  XOR2_X1 U753 ( .A(G116), .B(n684), .Z(G18) );
  XNOR2_X1 U754 ( .A(G125), .B(n685), .ZN(n686) );
  XNOR2_X1 U755 ( .A(n686), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U756 ( .A(G134), .B(n687), .ZN(G36) );
  NAND2_X1 U757 ( .A1(n688), .A2(n399), .ZN(n689) );
  XNOR2_X1 U758 ( .A(n689), .B(KEYINPUT92), .ZN(n691) );
  NAND2_X1 U759 ( .A1(n761), .A2(n399), .ZN(n690) );
  NAND2_X1 U760 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U761 ( .A(n692), .B(KEYINPUT88), .ZN(n694) );
  NOR2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n730) );
  XOR2_X1 U763 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n698) );
  NOR2_X1 U764 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U765 ( .A(n698), .B(n697), .Z(n699) );
  XNOR2_X1 U766 ( .A(n699), .B(KEYINPUT115), .ZN(n700) );
  NOR2_X1 U767 ( .A1(n570), .A2(n700), .ZN(n701) );
  XOR2_X1 U768 ( .A(KEYINPUT117), .B(n701), .Z(n707) );
  OR2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U770 ( .A(n704), .B(KEYINPUT118), .ZN(n705) );
  XNOR2_X1 U771 ( .A(KEYINPUT50), .B(n705), .ZN(n706) );
  NAND2_X1 U772 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U774 ( .A(KEYINPUT51), .B(n710), .ZN(n711) );
  NOR2_X1 U775 ( .A1(n711), .A2(n725), .ZN(n721) );
  INV_X1 U776 ( .A(n713), .ZN(n717) );
  NOR2_X1 U777 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U778 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U779 ( .A1(n356), .A2(n718), .ZN(n719) );
  NOR2_X1 U780 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U781 ( .A(n722), .B(KEYINPUT52), .ZN(n723) );
  NOR2_X1 U782 ( .A1(n724), .A2(n723), .ZN(n728) );
  NAND2_X1 U783 ( .A1(n726), .A2(n762), .ZN(n727) );
  OR2_X1 U784 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U785 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U786 ( .A(n731), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U787 ( .A1(n737), .A2(G478), .ZN(n734) );
  XOR2_X1 U788 ( .A(n732), .B(KEYINPUT121), .Z(n733) );
  XNOR2_X1 U789 ( .A(n734), .B(n733), .ZN(n735) );
  NOR2_X2 U790 ( .A1(n735), .A2(n742), .ZN(n736) );
  XNOR2_X1 U791 ( .A(n736), .B(KEYINPUT122), .ZN(G63) );
  NAND2_X1 U792 ( .A1(n737), .A2(G217), .ZN(n740) );
  XOR2_X1 U793 ( .A(KEYINPUT123), .B(n738), .Z(n739) );
  XNOR2_X1 U794 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U795 ( .A1(n742), .A2(n741), .ZN(G66) );
  XOR2_X1 U796 ( .A(n744), .B(G101), .Z(n745) );
  XNOR2_X1 U797 ( .A(n743), .B(n745), .ZN(n747) );
  NAND2_X1 U798 ( .A1(n747), .A2(n746), .ZN(n755) );
  INV_X1 U799 ( .A(n688), .ZN(n748) );
  NAND2_X1 U800 ( .A1(n748), .A2(n762), .ZN(n753) );
  NAND2_X1 U801 ( .A1(G953), .A2(G224), .ZN(n749) );
  XNOR2_X1 U802 ( .A(KEYINPUT61), .B(n749), .ZN(n750) );
  NAND2_X1 U803 ( .A1(n750), .A2(G898), .ZN(n751) );
  XNOR2_X1 U804 ( .A(n751), .B(KEYINPUT124), .ZN(n752) );
  NAND2_X1 U805 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U806 ( .A(n755), .B(n754), .ZN(n756) );
  XNOR2_X1 U807 ( .A(KEYINPUT125), .B(n756), .ZN(G69) );
  XNOR2_X1 U808 ( .A(n757), .B(n758), .ZN(n759) );
  XNOR2_X1 U809 ( .A(n760), .B(n759), .ZN(n765) );
  XNOR2_X1 U810 ( .A(n761), .B(n765), .ZN(n763) );
  NAND2_X1 U811 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U812 ( .A(n764), .B(KEYINPUT126), .ZN(n769) );
  XNOR2_X1 U813 ( .A(G227), .B(n765), .ZN(n766) );
  NAND2_X1 U814 ( .A1(n766), .A2(G900), .ZN(n767) );
  NAND2_X1 U815 ( .A1(G953), .A2(n767), .ZN(n768) );
  NAND2_X1 U816 ( .A1(n769), .A2(n768), .ZN(G72) );
  XOR2_X1 U817 ( .A(G131), .B(n770), .Z(G33) );
endmodule

