

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775;

  NOR2_X1 U375 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U376 ( .A(n547), .B(KEYINPUT85), .ZN(n565) );
  XNOR2_X2 U377 ( .A(n388), .B(n534), .ZN(n578) );
  NOR2_X2 U378 ( .A1(n774), .A2(n603), .ZN(n604) );
  NOR2_X2 U379 ( .A1(n555), .A2(KEYINPUT44), .ZN(n556) );
  XNOR2_X2 U380 ( .A(n550), .B(n357), .ZN(n725) );
  XNOR2_X2 U381 ( .A(n427), .B(n426), .ZN(n570) );
  XNOR2_X1 U382 ( .A(G113), .B(G101), .ZN(n378) );
  AND2_X1 U383 ( .A1(n692), .A2(G217), .ZN(n650) );
  AND2_X1 U384 ( .A1(n354), .A2(n390), .ZN(n371) );
  AND2_X1 U385 ( .A1(n417), .A2(n415), .ZN(n414) );
  AND2_X1 U386 ( .A1(n360), .A2(n400), .ZN(n398) );
  XNOR2_X1 U387 ( .A(n546), .B(KEYINPUT73), .ZN(n569) );
  XNOR2_X1 U388 ( .A(n379), .B(n378), .ZN(n377) );
  XNOR2_X1 U389 ( .A(n376), .B(KEYINPUT3), .ZN(n375) );
  XNOR2_X1 U390 ( .A(n381), .B(n421), .ZN(n505) );
  XNOR2_X1 U391 ( .A(G110), .B(G107), .ZN(n381) );
  XNOR2_X1 U392 ( .A(KEYINPUT78), .B(KEYINPUT98), .ZN(n379) );
  XNOR2_X1 U393 ( .A(G119), .B(G116), .ZN(n376) );
  BUF_X1 U394 ( .A(n609), .Z(n353) );
  XNOR2_X1 U395 ( .A(n377), .B(n375), .ZN(n506) );
  XNOR2_X1 U396 ( .A(n511), .B(n510), .ZN(n609) );
  OR2_X1 U397 ( .A1(n609), .A2(n521), .ZN(n606) );
  AND2_X1 U398 ( .A1(n736), .A2(n373), .ZN(n518) );
  NOR2_X1 U399 ( .A1(n735), .A2(n374), .ZN(n373) );
  INV_X1 U400 ( .A(n596), .ZN(n374) );
  XNOR2_X1 U401 ( .A(n425), .B(G469), .ZN(n426) );
  NOR2_X1 U402 ( .A1(G902), .A2(n693), .ZN(n427) );
  XNOR2_X1 U403 ( .A(n573), .B(n362), .ZN(n361) );
  INV_X1 U404 ( .A(KEYINPUT105), .ZN(n362) );
  XNOR2_X1 U405 ( .A(n367), .B(n453), .ZN(n474) );
  XNOR2_X1 U406 ( .A(n452), .B(n451), .ZN(n367) );
  XOR2_X1 U407 ( .A(G104), .B(G113), .Z(n435) );
  XNOR2_X1 U408 ( .A(n428), .B(G125), .ZN(n496) );
  INV_X1 U409 ( .A(G146), .ZN(n428) );
  XNOR2_X1 U410 ( .A(n407), .B(KEYINPUT96), .ZN(n390) );
  AND2_X1 U411 ( .A1(n575), .A2(n518), .ZN(n488) );
  NAND2_X1 U412 ( .A1(n408), .A2(n574), .ZN(n547) );
  NAND2_X1 U413 ( .A1(n385), .A2(n382), .ZN(n566) );
  AND2_X1 U414 ( .A1(n387), .A2(n386), .ZN(n385) );
  NAND2_X1 U415 ( .A1(n384), .A2(n383), .ZN(n382) );
  NAND2_X1 U416 ( .A1(n530), .A2(n531), .ZN(n386) );
  XNOR2_X1 U417 ( .A(n487), .B(n486), .ZN(n545) );
  XNOR2_X1 U418 ( .A(n506), .B(n380), .ZN(n676) );
  XNOR2_X1 U419 ( .A(n505), .B(n504), .ZN(n380) );
  XNOR2_X1 U420 ( .A(KEYINPUT83), .B(KEYINPUT16), .ZN(n503) );
  XNOR2_X1 U421 ( .A(n496), .B(n365), .ZN(n764) );
  XNOR2_X1 U422 ( .A(G140), .B(KEYINPUT10), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n476), .B(n363), .ZN(n478) );
  XNOR2_X1 U424 ( .A(n475), .B(n364), .ZN(n363) );
  INV_X1 U425 ( .A(G110), .ZN(n364) );
  INV_X1 U426 ( .A(n409), .ZN(n410) );
  XNOR2_X1 U427 ( .A(n606), .B(n523), .ZN(n621) );
  XNOR2_X1 U428 ( .A(n372), .B(n358), .ZN(n519) );
  NAND2_X1 U429 ( .A1(n518), .A2(n593), .ZN(n372) );
  INV_X1 U430 ( .A(n578), .ZN(n540) );
  NAND2_X1 U431 ( .A1(G953), .A2(G902), .ZN(n524) );
  AND2_X1 U432 ( .A1(n389), .A2(KEYINPUT0), .ZN(n383) );
  NOR2_X1 U433 ( .A1(G953), .A2(G237), .ZN(n434) );
  XNOR2_X1 U434 ( .A(G119), .B(KEYINPUT23), .ZN(n475) );
  XNOR2_X1 U435 ( .A(n500), .B(n392), .ZN(n391) );
  XNOR2_X1 U436 ( .A(G131), .B(G137), .ZN(n392) );
  XNOR2_X1 U437 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n500) );
  NAND2_X1 U438 ( .A1(n488), .A2(n405), .ZN(n404) );
  NOR2_X1 U439 ( .A1(n403), .A2(n606), .ZN(n402) );
  AND2_X1 U440 ( .A1(n416), .A2(n553), .ZN(n415) );
  NAND2_X1 U441 ( .A1(n571), .A2(KEYINPUT34), .ZN(n416) );
  XNOR2_X1 U442 ( .A(n570), .B(n411), .ZN(n574) );
  XNOR2_X1 U443 ( .A(G116), .B(G107), .ZN(n444) );
  XNOR2_X1 U444 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U445 ( .A(G101), .B(G140), .Z(n419) );
  XNOR2_X1 U446 ( .A(n763), .B(G146), .ZN(n464) );
  AND2_X1 U447 ( .A1(n368), .A2(n356), .ZN(n646) );
  INV_X1 U448 ( .A(KEYINPUT48), .ZN(n369) );
  BUF_X1 U449 ( .A(n679), .Z(n720) );
  INV_X1 U450 ( .A(KEYINPUT41), .ZN(n516) );
  NOR2_X1 U451 ( .A1(n731), .A2(n726), .ZN(n517) );
  OR2_X1 U452 ( .A1(n488), .A2(n393), .ZN(n400) );
  NAND2_X1 U453 ( .A1(KEYINPUT36), .A2(n406), .ZN(n393) );
  OR2_X1 U454 ( .A1(n488), .A2(KEYINPUT119), .ZN(n401) );
  NAND2_X1 U455 ( .A1(n508), .A2(n636), .ZN(n511) );
  OR2_X1 U456 ( .A1(n563), .A2(n562), .ZN(n601) );
  NAND2_X1 U457 ( .A1(n566), .A2(n532), .ZN(n388) );
  BUF_X1 U458 ( .A(n574), .Z(n409) );
  INV_X2 U459 ( .A(G953), .ZN(n766) );
  XNOR2_X1 U460 ( .A(n366), .B(n764), .ZN(n480) );
  BUF_X1 U461 ( .A(n555), .Z(n582) );
  NOR2_X1 U462 ( .A1(n745), .A2(n571), .ZN(n568) );
  NOR2_X1 U463 ( .A1(n622), .A2(n621), .ZN(n707) );
  INV_X1 U464 ( .A(n407), .ZN(n715) );
  XNOR2_X1 U465 ( .A(n466), .B(n465), .ZN(n738) );
  XNOR2_X1 U466 ( .A(n495), .B(G134), .ZN(n450) );
  AND2_X1 U467 ( .A1(n631), .A2(n630), .ZN(n354) );
  INV_X1 U468 ( .A(n530), .ZN(n389) );
  AND2_X1 U469 ( .A1(n566), .A2(n551), .ZN(n355) );
  AND2_X1 U470 ( .A1(n635), .A2(n717), .ZN(n356) );
  BUF_X1 U471 ( .A(n545), .Z(n736) );
  XOR2_X1 U472 ( .A(KEYINPUT79), .B(KEYINPUT33), .Z(n357) );
  XOR2_X1 U473 ( .A(KEYINPUT117), .B(KEYINPUT28), .Z(n358) );
  INV_X1 U474 ( .A(KEYINPUT119), .ZN(n406) );
  XOR2_X1 U475 ( .A(KEYINPUT95), .B(KEYINPUT45), .Z(n359) );
  XNOR2_X1 U476 ( .A(n450), .B(n391), .ZN(n763) );
  XNOR2_X1 U477 ( .A(n464), .B(n424), .ZN(n693) );
  NAND2_X1 U478 ( .A1(n399), .A2(KEYINPUT36), .ZN(n360) );
  XNOR2_X1 U479 ( .A(n370), .B(n369), .ZN(n368) );
  XNOR2_X1 U480 ( .A(n480), .B(n479), .ZN(n651) );
  NOR2_X1 U481 ( .A1(n361), .A2(n727), .ZN(n580) );
  NOR2_X1 U482 ( .A1(n588), .A2(n589), .ZN(n590) );
  NAND2_X1 U483 ( .A1(n557), .A2(n558), .ZN(n559) );
  NAND2_X1 U484 ( .A1(n537), .A2(n736), .ZN(n557) );
  NAND2_X1 U485 ( .A1(n632), .A2(n371), .ZN(n370) );
  NAND2_X1 U486 ( .A1(n474), .A2(G221), .ZN(n366) );
  NAND2_X1 U487 ( .A1(n621), .A2(n531), .ZN(n387) );
  INV_X1 U488 ( .A(n621), .ZN(n384) );
  NAND2_X1 U489 ( .A1(n394), .A2(n401), .ZN(n397) );
  NOR2_X1 U490 ( .A1(n396), .A2(n395), .ZN(n394) );
  INV_X1 U491 ( .A(n404), .ZN(n395) );
  NAND2_X1 U492 ( .A1(n402), .A2(n607), .ZN(n396) );
  NAND2_X1 U493 ( .A1(n398), .A2(n397), .ZN(n608) );
  NAND2_X1 U494 ( .A1(n404), .A2(n402), .ZN(n399) );
  NAND2_X1 U495 ( .A1(n488), .A2(n489), .ZN(n605) );
  NOR2_X1 U496 ( .A1(n489), .A2(KEYINPUT119), .ZN(n403) );
  AND2_X1 U497 ( .A1(n489), .A2(KEYINPUT119), .ZN(n405) );
  OR2_X2 U498 ( .A1(n608), .A2(n410), .ZN(n407) );
  INV_X1 U499 ( .A(n569), .ZN(n408) );
  NAND2_X1 U500 ( .A1(n409), .A2(n736), .ZN(n538) );
  NOR2_X1 U501 ( .A1(n409), .A2(n593), .ZN(n535) );
  NAND2_X1 U502 ( .A1(n569), .A2(n410), .ZN(n741) );
  INV_X1 U503 ( .A(KEYINPUT1), .ZN(n411) );
  XNOR2_X2 U504 ( .A(G143), .B(G128), .ZN(n495) );
  NAND2_X1 U505 ( .A1(n725), .A2(n355), .ZN(n417) );
  NAND2_X1 U506 ( .A1(n414), .A2(n412), .ZN(n554) );
  NAND2_X1 U507 ( .A1(n413), .A2(KEYINPUT34), .ZN(n412) );
  INV_X1 U508 ( .A(n725), .ZN(n413) );
  AND2_X2 U509 ( .A1(n649), .A2(n723), .ZN(n667) );
  NOR2_X1 U510 ( .A1(n519), .A2(n570), .ZN(n620) );
  INV_X1 U511 ( .A(KEYINPUT76), .ZN(n451) );
  XNOR2_X1 U512 ( .A(n764), .B(n433), .ZN(n440) );
  INV_X1 U513 ( .A(KEYINPUT36), .ZN(n607) );
  BUF_X1 U514 ( .A(n719), .Z(n765) );
  INV_X1 U515 ( .A(KEYINPUT31), .ZN(n567) );
  NAND2_X1 U516 ( .A1(G227), .A2(n766), .ZN(n418) );
  XNOR2_X1 U517 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U518 ( .A(n420), .B(KEYINPUT90), .Z(n423) );
  INV_X1 U519 ( .A(G104), .ZN(n421) );
  XOR2_X1 U520 ( .A(KEYINPUT101), .B(n505), .Z(n422) );
  XNOR2_X1 U521 ( .A(n423), .B(n422), .ZN(n424) );
  INV_X1 U522 ( .A(KEYINPUT77), .ZN(n425) );
  XOR2_X1 U523 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n430) );
  XNOR2_X1 U524 ( .A(G122), .B(KEYINPUT108), .ZN(n429) );
  XNOR2_X1 U525 ( .A(n430), .B(n429), .ZN(n432) );
  XOR2_X1 U526 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n431) );
  XNOR2_X1 U527 ( .A(G143), .B(G131), .ZN(n438) );
  XOR2_X1 U528 ( .A(KEYINPUT87), .B(n434), .Z(n459) );
  NAND2_X1 U529 ( .A1(G214), .A2(n459), .ZN(n436) );
  XNOR2_X1 U530 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U531 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U532 ( .A(n439), .B(n440), .ZN(n655) );
  NOR2_X1 U533 ( .A1(G902), .A2(n655), .ZN(n442) );
  XNOR2_X1 U534 ( .A(KEYINPUT109), .B(KEYINPUT13), .ZN(n441) );
  XNOR2_X1 U535 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U536 ( .A(n443), .B(G475), .ZN(n563) );
  XOR2_X1 U537 ( .A(KEYINPUT9), .B(G122), .Z(n445) );
  XNOR2_X1 U538 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U539 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n447) );
  XNOR2_X1 U540 ( .A(KEYINPUT7), .B(KEYINPUT110), .ZN(n446) );
  XNOR2_X1 U541 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U542 ( .A(n449), .B(n448), .Z(n456) );
  NAND2_X1 U543 ( .A1(G234), .A2(n766), .ZN(n452) );
  XOR2_X1 U544 ( .A(KEYINPUT8), .B(KEYINPUT75), .Z(n453) );
  AND2_X1 U545 ( .A1(G217), .A2(n474), .ZN(n454) );
  XNOR2_X1 U546 ( .A(n450), .B(n454), .ZN(n455) );
  XNOR2_X1 U547 ( .A(n456), .B(n455), .ZN(n688) );
  INV_X1 U548 ( .A(G902), .ZN(n491) );
  NAND2_X1 U549 ( .A1(n688), .A2(n491), .ZN(n458) );
  INV_X1 U550 ( .A(G478), .ZN(n457) );
  XNOR2_X1 U551 ( .A(n458), .B(n457), .ZN(n513) );
  INV_X1 U552 ( .A(n513), .ZN(n562) );
  INV_X1 U553 ( .A(n601), .ZN(n489) );
  NAND2_X1 U554 ( .A1(n459), .A2(G210), .ZN(n461) );
  XOR2_X1 U555 ( .A(KEYINPUT5), .B(KEYINPUT86), .Z(n460) );
  XNOR2_X1 U556 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U557 ( .A(n462), .B(n506), .ZN(n463) );
  XNOR2_X1 U558 ( .A(n464), .B(n463), .ZN(n662) );
  NAND2_X1 U559 ( .A1(n662), .A2(n491), .ZN(n466) );
  INV_X1 U560 ( .A(G472), .ZN(n465) );
  XNOR2_X1 U561 ( .A(n738), .B(KEYINPUT6), .ZN(n575) );
  XNOR2_X1 U562 ( .A(G902), .B(KEYINPUT15), .ZN(n636) );
  NAND2_X1 U563 ( .A1(n636), .A2(G234), .ZN(n467) );
  XNOR2_X1 U564 ( .A(n467), .B(KEYINPUT20), .ZN(n481) );
  NAND2_X1 U565 ( .A1(G221), .A2(n481), .ZN(n468) );
  XNOR2_X1 U566 ( .A(n468), .B(KEYINPUT21), .ZN(n735) );
  NAND2_X1 U567 ( .A1(n766), .A2(G952), .ZN(n526) );
  INV_X1 U568 ( .A(n526), .ZN(n470) );
  NOR2_X1 U569 ( .A1(G900), .A2(n524), .ZN(n469) );
  NOR2_X1 U570 ( .A1(n470), .A2(n469), .ZN(n473) );
  NAND2_X1 U571 ( .A1(G237), .A2(G234), .ZN(n472) );
  INV_X1 U572 ( .A(KEYINPUT14), .ZN(n471) );
  XNOR2_X1 U573 ( .A(n472), .B(n471), .ZN(n754) );
  NOR2_X1 U574 ( .A1(n473), .A2(n754), .ZN(n596) );
  XOR2_X1 U575 ( .A(KEYINPUT24), .B(KEYINPUT102), .Z(n476) );
  XNOR2_X1 U576 ( .A(G137), .B(G128), .ZN(n477) );
  XNOR2_X1 U577 ( .A(n478), .B(n477), .ZN(n479) );
  NAND2_X1 U578 ( .A1(n651), .A2(n491), .ZN(n487) );
  XOR2_X1 U579 ( .A(KEYINPUT25), .B(KEYINPUT103), .Z(n483) );
  NAND2_X1 U580 ( .A1(n481), .A2(G217), .ZN(n482) );
  XNOR2_X1 U581 ( .A(n483), .B(n482), .ZN(n485) );
  INV_X1 U582 ( .A(KEYINPUT89), .ZN(n484) );
  XNOR2_X1 U583 ( .A(n485), .B(n484), .ZN(n486) );
  NOR2_X1 U584 ( .A1(n409), .A2(n605), .ZN(n492) );
  INV_X1 U585 ( .A(G237), .ZN(n490) );
  NAND2_X1 U586 ( .A1(n491), .A2(n490), .ZN(n509) );
  NAND2_X1 U587 ( .A1(n509), .A2(G214), .ZN(n728) );
  NAND2_X1 U588 ( .A1(n492), .A2(n728), .ZN(n493) );
  XNOR2_X1 U589 ( .A(n493), .B(KEYINPUT43), .ZN(n512) );
  XNOR2_X1 U590 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n494) );
  XNOR2_X1 U591 ( .A(n495), .B(n494), .ZN(n497) );
  XNOR2_X1 U592 ( .A(n497), .B(n496), .ZN(n502) );
  NAND2_X1 U593 ( .A1(n766), .A2(G224), .ZN(n498) );
  XNOR2_X1 U594 ( .A(n498), .B(KEYINPUT99), .ZN(n499) );
  XNOR2_X1 U595 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U596 ( .A(n502), .B(n501), .ZN(n507) );
  XNOR2_X1 U597 ( .A(n503), .B(G122), .ZN(n504) );
  XNOR2_X1 U598 ( .A(n507), .B(n676), .ZN(n669) );
  INV_X1 U599 ( .A(n669), .ZN(n508) );
  NAND2_X1 U600 ( .A1(n509), .A2(G210), .ZN(n510) );
  NAND2_X1 U601 ( .A1(n512), .A2(n353), .ZN(n635) );
  XNOR2_X1 U602 ( .A(n635), .B(G140), .ZN(G42) );
  NAND2_X1 U603 ( .A1(n563), .A2(n513), .ZN(n731) );
  XNOR2_X1 U604 ( .A(KEYINPUT84), .B(KEYINPUT38), .ZN(n514) );
  XNOR2_X1 U605 ( .A(n609), .B(n514), .ZN(n729) );
  NAND2_X1 U606 ( .A1(n729), .A2(n728), .ZN(n515) );
  XNOR2_X1 U607 ( .A(n515), .B(KEYINPUT118), .ZN(n726) );
  XNOR2_X1 U608 ( .A(n517), .B(n516), .ZN(n756) );
  INV_X1 U609 ( .A(n738), .ZN(n593) );
  NAND2_X1 U610 ( .A1(n756), .A2(n620), .ZN(n520) );
  XOR2_X1 U611 ( .A(KEYINPUT42), .B(n520), .Z(n603) );
  XOR2_X1 U612 ( .A(n603), .B(G137), .Z(G39) );
  XNOR2_X1 U613 ( .A(n735), .B(KEYINPUT104), .ZN(n544) );
  NOR2_X1 U614 ( .A1(n731), .A2(n544), .ZN(n532) );
  INV_X1 U615 ( .A(n728), .ZN(n521) );
  XNOR2_X1 U616 ( .A(KEYINPUT88), .B(KEYINPUT19), .ZN(n522) );
  XNOR2_X1 U617 ( .A(n522), .B(KEYINPUT71), .ZN(n523) );
  XOR2_X1 U618 ( .A(KEYINPUT100), .B(G898), .Z(n682) );
  INV_X1 U619 ( .A(n524), .ZN(n525) );
  NAND2_X1 U620 ( .A1(n682), .A2(n525), .ZN(n527) );
  NAND2_X1 U621 ( .A1(n527), .A2(n526), .ZN(n529) );
  INV_X1 U622 ( .A(n754), .ZN(n528) );
  NAND2_X1 U623 ( .A1(n529), .A2(n528), .ZN(n530) );
  INV_X1 U624 ( .A(KEYINPUT0), .ZN(n531) );
  XNOR2_X1 U625 ( .A(KEYINPUT82), .B(KEYINPUT22), .ZN(n533) );
  XNOR2_X1 U626 ( .A(n533), .B(KEYINPUT68), .ZN(n534) );
  NAND2_X1 U627 ( .A1(n540), .A2(n535), .ZN(n536) );
  XNOR2_X1 U628 ( .A(n536), .B(KEYINPUT67), .ZN(n537) );
  XNOR2_X1 U629 ( .A(n557), .B(G110), .ZN(G12) );
  NOR2_X1 U630 ( .A1(n538), .A2(n575), .ZN(n539) );
  XNOR2_X1 U631 ( .A(n539), .B(KEYINPUT92), .ZN(n541) );
  NAND2_X1 U632 ( .A1(n541), .A2(n540), .ZN(n543) );
  XNOR2_X1 U633 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n542) );
  XNOR2_X1 U634 ( .A(n543), .B(n542), .ZN(n558) );
  XNOR2_X1 U635 ( .A(n558), .B(G119), .ZN(G21) );
  INV_X1 U636 ( .A(KEYINPUT115), .ZN(n548) );
  XNOR2_X1 U637 ( .A(n565), .B(n548), .ZN(n549) );
  NAND2_X1 U638 ( .A1(n549), .A2(n575), .ZN(n550) );
  INV_X1 U639 ( .A(KEYINPUT34), .ZN(n551) );
  INV_X1 U640 ( .A(n563), .ZN(n552) );
  NAND2_X1 U641 ( .A1(n552), .A2(n562), .ZN(n610) );
  XNOR2_X1 U642 ( .A(n610), .B(KEYINPUT91), .ZN(n553) );
  XNOR2_X1 U643 ( .A(n554), .B(KEYINPUT35), .ZN(n555) );
  XOR2_X1 U644 ( .A(n582), .B(G122), .Z(G24) );
  XNOR2_X1 U645 ( .A(n556), .B(KEYINPUT72), .ZN(n560) );
  XNOR2_X1 U646 ( .A(n559), .B(KEYINPUT97), .ZN(n585) );
  NAND2_X1 U647 ( .A1(n560), .A2(n585), .ZN(n561) );
  XNOR2_X1 U648 ( .A(n561), .B(KEYINPUT80), .ZN(n591) );
  NAND2_X1 U649 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U650 ( .A(n564), .B(KEYINPUT113), .ZN(n710) );
  OR2_X1 U651 ( .A1(n710), .A2(n489), .ZN(n619) );
  INV_X1 U652 ( .A(n619), .ZN(n727) );
  NAND2_X1 U653 ( .A1(n565), .A2(n593), .ZN(n745) );
  INV_X1 U654 ( .A(n566), .ZN(n571) );
  XNOR2_X1 U655 ( .A(n568), .B(n567), .ZN(n711) );
  NOR2_X1 U656 ( .A1(n569), .A2(n570), .ZN(n595) );
  NAND2_X1 U657 ( .A1(n595), .A2(n738), .ZN(n572) );
  NOR2_X1 U658 ( .A1(n572), .A2(n571), .ZN(n701) );
  NOR2_X1 U659 ( .A1(n711), .A2(n701), .ZN(n573) );
  NOR2_X1 U660 ( .A1(n409), .A2(n736), .ZN(n577) );
  INV_X1 U661 ( .A(n575), .ZN(n576) );
  NAND2_X1 U662 ( .A1(n577), .A2(n576), .ZN(n579) );
  NOR2_X1 U663 ( .A1(n579), .A2(n578), .ZN(n699) );
  NOR2_X1 U664 ( .A1(n580), .A2(n699), .ZN(n581) );
  XNOR2_X1 U665 ( .A(n581), .B(KEYINPUT114), .ZN(n584) );
  NAND2_X1 U666 ( .A1(n582), .A2(KEYINPUT44), .ZN(n583) );
  NAND2_X1 U667 ( .A1(n584), .A2(n583), .ZN(n589) );
  INV_X1 U668 ( .A(n585), .ZN(n586) );
  NAND2_X1 U669 ( .A1(n586), .A2(KEYINPUT44), .ZN(n587) );
  XNOR2_X1 U670 ( .A(n587), .B(KEYINPUT65), .ZN(n588) );
  NAND2_X1 U671 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X2 U672 ( .A(n592), .B(n359), .ZN(n679) );
  NAND2_X1 U673 ( .A1(n593), .A2(n728), .ZN(n594) );
  XNOR2_X1 U674 ( .A(KEYINPUT30), .B(n594), .ZN(n598) );
  NAND2_X1 U675 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n612) );
  NAND2_X1 U677 ( .A1(n612), .A2(n729), .ZN(n600) );
  XNOR2_X1 U678 ( .A(KEYINPUT81), .B(KEYINPUT39), .ZN(n599) );
  XNOR2_X1 U679 ( .A(n600), .B(n599), .ZN(n634) );
  NOR2_X1 U680 ( .A1(n634), .A2(n601), .ZN(n602) );
  XNOR2_X1 U681 ( .A(n602), .B(KEYINPUT40), .ZN(n774) );
  XNOR2_X1 U682 ( .A(n604), .B(KEYINPUT46), .ZN(n632) );
  NOR2_X1 U683 ( .A1(n610), .A2(n353), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U685 ( .A(n613), .B(KEYINPUT116), .ZN(n775) );
  INV_X1 U686 ( .A(n775), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n614), .A2(KEYINPUT93), .ZN(n618) );
  NAND2_X1 U688 ( .A1(n727), .A2(KEYINPUT47), .ZN(n615) );
  NAND2_X1 U689 ( .A1(KEYINPUT93), .A2(n615), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n775), .A2(n616), .ZN(n617) );
  NAND2_X1 U691 ( .A1(n618), .A2(n617), .ZN(n631) );
  NAND2_X1 U692 ( .A1(KEYINPUT74), .A2(n619), .ZN(n625) );
  NOR2_X1 U693 ( .A1(KEYINPUT47), .A2(n625), .ZN(n623) );
  INV_X1 U694 ( .A(n620), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n623), .A2(n707), .ZN(n629) );
  NAND2_X1 U696 ( .A1(KEYINPUT93), .A2(n727), .ZN(n624) );
  NAND2_X1 U697 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U698 ( .A1(n707), .A2(n626), .ZN(n627) );
  NAND2_X1 U699 ( .A1(n627), .A2(KEYINPUT47), .ZN(n628) );
  AND2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n630) );
  INV_X1 U701 ( .A(n710), .ZN(n633) );
  OR2_X1 U702 ( .A1(n634), .A2(n633), .ZN(n717) );
  XNOR2_X1 U703 ( .A(n646), .B(KEYINPUT94), .ZN(n719) );
  INV_X1 U704 ( .A(n636), .ZN(n639) );
  AND2_X1 U705 ( .A1(n719), .A2(n639), .ZN(n637) );
  NAND2_X1 U706 ( .A1(n679), .A2(n637), .ZN(n645) );
  NAND2_X1 U707 ( .A1(KEYINPUT2), .A2(KEYINPUT70), .ZN(n638) );
  OR2_X1 U708 ( .A1(n636), .A2(n638), .ZN(n643) );
  NAND2_X1 U709 ( .A1(n639), .A2(KEYINPUT2), .ZN(n641) );
  INV_X1 U710 ( .A(KEYINPUT70), .ZN(n640) );
  NAND2_X1 U711 ( .A1(n641), .A2(n640), .ZN(n642) );
  AND2_X1 U712 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U713 ( .A1(n645), .A2(n644), .ZN(n649) );
  INV_X1 U714 ( .A(n646), .ZN(n647) );
  INV_X1 U715 ( .A(KEYINPUT2), .ZN(n721) );
  NOR2_X1 U716 ( .A1(n647), .A2(n721), .ZN(n648) );
  NAND2_X1 U717 ( .A1(n679), .A2(n648), .ZN(n723) );
  BUF_X2 U718 ( .A(n667), .Z(n692) );
  XNOR2_X1 U719 ( .A(n651), .B(n650), .ZN(n653) );
  INV_X1 U720 ( .A(G952), .ZN(n652) );
  NAND2_X1 U721 ( .A1(n652), .A2(G953), .ZN(n672) );
  INV_X1 U722 ( .A(n672), .ZN(n697) );
  NOR2_X1 U723 ( .A1(n653), .A2(n697), .ZN(G66) );
  NAND2_X1 U724 ( .A1(n667), .A2(G475), .ZN(n657) );
  XOR2_X1 U725 ( .A(KEYINPUT69), .B(KEYINPUT59), .Z(n654) );
  XNOR2_X1 U726 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U727 ( .A(n657), .B(n656), .ZN(n658) );
  NAND2_X1 U728 ( .A1(n658), .A2(n672), .ZN(n660) );
  INV_X1 U729 ( .A(KEYINPUT60), .ZN(n659) );
  XNOR2_X1 U730 ( .A(n660), .B(n659), .ZN(G60) );
  NAND2_X1 U731 ( .A1(n667), .A2(G472), .ZN(n664) );
  XNOR2_X1 U732 ( .A(KEYINPUT120), .B(KEYINPUT62), .ZN(n661) );
  XNOR2_X1 U733 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U734 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U735 ( .A1(n665), .A2(n672), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n666), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U737 ( .A1(n667), .A2(G210), .ZN(n671) );
  XNOR2_X1 U738 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n668) );
  XNOR2_X1 U739 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U740 ( .A(n671), .B(n670), .ZN(n673) );
  NAND2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n675) );
  INV_X1 U742 ( .A(KEYINPUT56), .ZN(n674) );
  XNOR2_X1 U743 ( .A(n675), .B(n674), .ZN(G51) );
  INV_X1 U744 ( .A(n676), .ZN(n678) );
  NAND2_X1 U745 ( .A1(G953), .A2(n682), .ZN(n677) );
  NAND2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n687) );
  NAND2_X1 U747 ( .A1(n720), .A2(n766), .ZN(n685) );
  NAND2_X1 U748 ( .A1(G953), .A2(G224), .ZN(n680) );
  XOR2_X1 U749 ( .A(KEYINPUT61), .B(n680), .Z(n681) );
  NOR2_X1 U750 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U751 ( .A(KEYINPUT126), .B(n683), .Z(n684) );
  NAND2_X1 U752 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U753 ( .A(n687), .B(n686), .Z(G69) );
  NAND2_X1 U754 ( .A1(n692), .A2(G478), .ZN(n690) );
  XNOR2_X1 U755 ( .A(n688), .B(KEYINPUT125), .ZN(n689) );
  XNOR2_X1 U756 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U757 ( .A1(n691), .A2(n697), .ZN(G63) );
  NAND2_X1 U758 ( .A1(n692), .A2(G469), .ZN(n696) );
  XOR2_X1 U759 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n694) );
  XNOR2_X1 U760 ( .A(n693), .B(n694), .ZN(n695) );
  XNOR2_X1 U761 ( .A(n696), .B(n695), .ZN(n698) );
  NOR2_X1 U762 ( .A1(n698), .A2(n697), .ZN(G54) );
  XOR2_X1 U763 ( .A(G101), .B(n699), .Z(G3) );
  NAND2_X1 U764 ( .A1(n701), .A2(n489), .ZN(n700) );
  XNOR2_X1 U765 ( .A(n700), .B(G104), .ZN(G6) );
  XOR2_X1 U766 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n703) );
  NAND2_X1 U767 ( .A1(n701), .A2(n710), .ZN(n702) );
  XNOR2_X1 U768 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U769 ( .A(G107), .B(n704), .ZN(G9) );
  XOR2_X1 U770 ( .A(G128), .B(KEYINPUT29), .Z(n706) );
  NAND2_X1 U771 ( .A1(n707), .A2(n710), .ZN(n705) );
  XNOR2_X1 U772 ( .A(n706), .B(n705), .ZN(G30) );
  NAND2_X1 U773 ( .A1(n707), .A2(n489), .ZN(n708) );
  XNOR2_X1 U774 ( .A(n708), .B(G146), .ZN(G48) );
  NAND2_X1 U775 ( .A1(n489), .A2(n711), .ZN(n709) );
  XNOR2_X1 U776 ( .A(G113), .B(n709), .ZN(G15) );
  XOR2_X1 U777 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n713) );
  NAND2_X1 U778 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U779 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U780 ( .A(G116), .B(n714), .ZN(G18) );
  XNOR2_X1 U781 ( .A(G125), .B(n715), .ZN(n716) );
  XNOR2_X1 U782 ( .A(n716), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 U783 ( .A(n717), .ZN(n718) );
  XOR2_X1 U784 ( .A(G134), .B(n718), .Z(G36) );
  NAND2_X1 U785 ( .A1(n720), .A2(n765), .ZN(n722) );
  NAND2_X1 U786 ( .A1(n722), .A2(n721), .ZN(n724) );
  AND2_X1 U787 ( .A1(n724), .A2(n723), .ZN(n761) );
  NOR2_X1 U788 ( .A1(n727), .A2(n726), .ZN(n733) );
  NOR2_X1 U789 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U790 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U791 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U792 ( .A1(n413), .A2(n734), .ZN(n750) );
  NAND2_X1 U793 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U794 ( .A(KEYINPUT49), .B(n737), .Z(n739) );
  NAND2_X1 U795 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U796 ( .A(KEYINPUT123), .B(n740), .ZN(n743) );
  XNOR2_X1 U797 ( .A(KEYINPUT50), .B(n741), .ZN(n742) );
  NAND2_X1 U798 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U799 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U800 ( .A(KEYINPUT51), .B(n746), .ZN(n748) );
  INV_X1 U801 ( .A(n756), .ZN(n747) );
  NOR2_X1 U802 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U803 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U804 ( .A(n751), .B(KEYINPUT124), .ZN(n752) );
  XNOR2_X1 U805 ( .A(KEYINPUT52), .B(n752), .ZN(n753) );
  NOR2_X1 U806 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U807 ( .A1(G952), .A2(n755), .ZN(n759) );
  AND2_X1 U808 ( .A1(n725), .A2(n756), .ZN(n757) );
  NOR2_X1 U809 ( .A1(n757), .A2(G953), .ZN(n758) );
  NAND2_X1 U810 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U811 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U812 ( .A(n762), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U813 ( .A(n763), .B(n764), .ZN(n768) );
  XOR2_X1 U814 ( .A(n768), .B(n765), .Z(n767) );
  NAND2_X1 U815 ( .A1(n767), .A2(n766), .ZN(n773) );
  XNOR2_X1 U816 ( .A(G227), .B(n768), .ZN(n769) );
  NAND2_X1 U817 ( .A1(n769), .A2(G900), .ZN(n770) );
  XOR2_X1 U818 ( .A(KEYINPUT127), .B(n770), .Z(n771) );
  NAND2_X1 U819 ( .A1(G953), .A2(n771), .ZN(n772) );
  NAND2_X1 U820 ( .A1(n773), .A2(n772), .ZN(G72) );
  XOR2_X1 U821 ( .A(G131), .B(n774), .Z(G33) );
  XNOR2_X1 U822 ( .A(G143), .B(n775), .ZN(G45) );
endmodule

