

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591;

  XNOR2_X1 U323 ( .A(n416), .B(KEYINPUT107), .ZN(n417) );
  XNOR2_X1 U324 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U325 ( .A(KEYINPUT108), .B(n454), .ZN(n478) );
  XOR2_X1 U326 ( .A(n395), .B(n394), .Z(n291) );
  XNOR2_X1 U327 ( .A(KEYINPUT115), .B(KEYINPUT46), .ZN(n501) );
  XNOR2_X1 U328 ( .A(n502), .B(n501), .ZN(n505) );
  XNOR2_X1 U329 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n517) );
  XNOR2_X1 U330 ( .A(n518), .B(n517), .ZN(n550) );
  INV_X1 U331 ( .A(KEYINPUT37), .ZN(n416) );
  XNOR2_X1 U332 ( .A(n450), .B(n449), .ZN(n452) );
  XNOR2_X1 U333 ( .A(n396), .B(n291), .ZN(n397) );
  XNOR2_X1 U334 ( .A(n418), .B(n417), .ZN(n491) );
  XNOR2_X1 U335 ( .A(n398), .B(n397), .ZN(n399) );
  NOR2_X1 U336 ( .A1(n559), .A2(n558), .ZN(n570) );
  INV_X1 U337 ( .A(G29GAT), .ZN(n455) );
  XNOR2_X1 U338 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U339 ( .A(n458), .B(n457), .ZN(G1328GAT) );
  XOR2_X1 U340 ( .A(G85GAT), .B(G162GAT), .Z(n294) );
  XNOR2_X1 U341 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n292) );
  XNOR2_X1 U342 ( .A(n292), .B(KEYINPUT83), .ZN(n356) );
  XNOR2_X1 U343 ( .A(G134GAT), .B(n356), .ZN(n293) );
  XNOR2_X1 U344 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U345 ( .A(G29GAT), .B(n295), .ZN(n316) );
  XOR2_X1 U346 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n297) );
  XNOR2_X1 U347 ( .A(KEYINPUT95), .B(KEYINPUT94), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U349 ( .A(KEYINPUT4), .B(n298), .Z(n300) );
  NAND2_X1 U350 ( .A1(G225GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U352 ( .A(n301), .B(KEYINPUT1), .Z(n306) );
  XOR2_X1 U353 ( .A(KEYINPUT92), .B(KEYINPUT2), .Z(n303) );
  XNOR2_X1 U354 ( .A(KEYINPUT91), .B(G155GAT), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U356 ( .A(KEYINPUT3), .B(n304), .Z(n386) );
  XNOR2_X1 U357 ( .A(n386), .B(KEYINPUT98), .ZN(n305) );
  XNOR2_X1 U358 ( .A(n306), .B(n305), .ZN(n314) );
  XOR2_X1 U359 ( .A(KEYINPUT97), .B(G57GAT), .Z(n308) );
  XNOR2_X1 U360 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U362 ( .A(G148GAT), .B(G120GAT), .Z(n310) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(G141GAT), .ZN(n309) );
  XNOR2_X1 U364 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U365 ( .A(n312), .B(n311), .Z(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n316), .B(n315), .ZN(n552) );
  XOR2_X1 U368 ( .A(G29GAT), .B(G36GAT), .Z(n318) );
  XNOR2_X1 U369 ( .A(G50GAT), .B(G43GAT), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U371 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n320) );
  XNOR2_X1 U372 ( .A(KEYINPUT70), .B(KEYINPUT69), .ZN(n319) );
  XNOR2_X1 U373 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n451) );
  XOR2_X1 U375 ( .A(G218GAT), .B(G162GAT), .Z(n380) );
  XOR2_X1 U376 ( .A(KEYINPUT78), .B(n380), .Z(n324) );
  NAND2_X1 U377 ( .A1(G232GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U379 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n326) );
  XNOR2_X1 U380 ( .A(KEYINPUT66), .B(KEYINPUT9), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U382 ( .A(n328), .B(n327), .Z(n333) );
  XOR2_X1 U383 ( .A(G190GAT), .B(G134GAT), .Z(n355) );
  XOR2_X1 U384 ( .A(KEYINPUT75), .B(G92GAT), .Z(n330) );
  XNOR2_X1 U385 ( .A(G99GAT), .B(G85GAT), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U387 ( .A(G106GAT), .B(n331), .Z(n431) );
  XNOR2_X1 U388 ( .A(n355), .B(n431), .ZN(n332) );
  XNOR2_X1 U389 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n451), .B(n334), .ZN(n509) );
  INV_X1 U391 ( .A(n509), .ZN(n546) );
  XOR2_X1 U392 ( .A(KEYINPUT79), .B(n546), .Z(n571) );
  INV_X1 U393 ( .A(n571), .ZN(n459) );
  XNOR2_X1 U394 ( .A(KEYINPUT36), .B(n459), .ZN(n588) );
  XOR2_X1 U395 ( .A(G57GAT), .B(KEYINPUT13), .Z(n426) );
  XOR2_X1 U396 ( .A(G127GAT), .B(G71GAT), .Z(n336) );
  XNOR2_X1 U397 ( .A(G15GAT), .B(G183GAT), .ZN(n335) );
  XNOR2_X1 U398 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U399 ( .A(n426), .B(n337), .Z(n339) );
  NAND2_X1 U400 ( .A1(G231GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U401 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U402 ( .A(n340), .B(KEYINPUT80), .Z(n343) );
  XNOR2_X1 U403 ( .A(G1GAT), .B(KEYINPUT71), .ZN(n341) );
  XNOR2_X1 U404 ( .A(n341), .B(G8GAT), .ZN(n435) );
  XNOR2_X1 U405 ( .A(n435), .B(G64GAT), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n351) );
  XOR2_X1 U407 ( .A(G78GAT), .B(G211GAT), .Z(n345) );
  XNOR2_X1 U408 ( .A(G22GAT), .B(G155GAT), .ZN(n344) );
  XNOR2_X1 U409 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U410 ( .A(KEYINPUT12), .B(KEYINPUT81), .Z(n347) );
  XNOR2_X1 U411 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n346) );
  XNOR2_X1 U412 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U413 ( .A(n349), .B(n348), .Z(n350) );
  XNOR2_X1 U414 ( .A(n351), .B(n350), .ZN(n567) );
  INV_X1 U415 ( .A(n567), .ZN(n585) );
  XOR2_X1 U416 ( .A(KEYINPUT86), .B(KEYINPUT17), .Z(n353) );
  XNOR2_X1 U417 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U419 ( .A(KEYINPUT19), .B(n354), .Z(n400) );
  XOR2_X1 U420 ( .A(n356), .B(n355), .Z(n358) );
  XNOR2_X1 U421 ( .A(G43GAT), .B(G99GAT), .ZN(n357) );
  XNOR2_X1 U422 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n400), .B(n359), .ZN(n368) );
  XOR2_X1 U424 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n361) );
  NAND2_X1 U425 ( .A1(G227GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U427 ( .A(n362), .B(KEYINPUT84), .Z(n366) );
  XNOR2_X1 U428 ( .A(G169GAT), .B(G15GAT), .ZN(n363) );
  XNOR2_X1 U429 ( .A(n363), .B(G113GAT), .ZN(n444) );
  XNOR2_X1 U430 ( .A(G71GAT), .B(G176GAT), .ZN(n364) );
  XNOR2_X1 U431 ( .A(n364), .B(G120GAT), .ZN(n422) );
  XNOR2_X1 U432 ( .A(n444), .B(n422), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n559) );
  INV_X1 U435 ( .A(n559), .ZN(n521) );
  XOR2_X1 U436 ( .A(KEYINPUT24), .B(KEYINPUT88), .Z(n370) );
  NAND2_X1 U437 ( .A1(G228GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U438 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U439 ( .A(G204GAT), .B(n371), .ZN(n384) );
  XOR2_X1 U440 ( .A(KEYINPUT22), .B(KEYINPUT93), .Z(n373) );
  XNOR2_X1 U441 ( .A(KEYINPUT89), .B(KEYINPUT23), .ZN(n372) );
  XNOR2_X1 U442 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U443 ( .A(n374), .B(G106GAT), .Z(n376) );
  XOR2_X1 U444 ( .A(G148GAT), .B(G78GAT), .Z(n432) );
  XNOR2_X1 U445 ( .A(G50GAT), .B(n432), .ZN(n375) );
  XNOR2_X1 U446 ( .A(n376), .B(n375), .ZN(n379) );
  XOR2_X1 U447 ( .A(G211GAT), .B(KEYINPUT21), .Z(n378) );
  XNOR2_X1 U448 ( .A(G197GAT), .B(KEYINPUT90), .ZN(n377) );
  XNOR2_X1 U449 ( .A(n378), .B(n377), .ZN(n388) );
  XOR2_X1 U450 ( .A(n379), .B(n388), .Z(n382) );
  XOR2_X1 U451 ( .A(G141GAT), .B(G22GAT), .Z(n436) );
  XNOR2_X1 U452 ( .A(n436), .B(n380), .ZN(n381) );
  XNOR2_X1 U453 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U454 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U455 ( .A(n386), .B(n385), .ZN(n555) );
  NOR2_X1 U456 ( .A1(n521), .A2(n555), .ZN(n387) );
  XNOR2_X1 U457 ( .A(KEYINPUT26), .B(n387), .ZN(n576) );
  XOR2_X1 U458 ( .A(G204GAT), .B(G64GAT), .Z(n425) );
  XOR2_X1 U459 ( .A(n425), .B(G92GAT), .Z(n390) );
  XNOR2_X1 U460 ( .A(G218GAT), .B(n388), .ZN(n389) );
  XNOR2_X1 U461 ( .A(n390), .B(n389), .ZN(n398) );
  XOR2_X1 U462 ( .A(G190GAT), .B(G176GAT), .Z(n392) );
  XNOR2_X1 U463 ( .A(G169GAT), .B(G36GAT), .ZN(n391) );
  XNOR2_X1 U464 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U465 ( .A(G8GAT), .B(n393), .ZN(n396) );
  XOR2_X1 U466 ( .A(KEYINPUT99), .B(KEYINPUT80), .Z(n395) );
  NAND2_X1 U467 ( .A1(G226GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U468 ( .A(n400), .B(n399), .ZN(n549) );
  XOR2_X1 U469 ( .A(KEYINPUT27), .B(KEYINPUT100), .Z(n401) );
  XOR2_X1 U470 ( .A(n549), .B(n401), .Z(n409) );
  INV_X1 U471 ( .A(n409), .ZN(n402) );
  NAND2_X1 U472 ( .A1(n576), .A2(n402), .ZN(n407) );
  OR2_X1 U473 ( .A1(n559), .A2(n549), .ZN(n403) );
  NAND2_X1 U474 ( .A1(n403), .A2(n555), .ZN(n404) );
  XNOR2_X1 U475 ( .A(n404), .B(KEYINPUT102), .ZN(n405) );
  XOR2_X1 U476 ( .A(KEYINPUT25), .B(n405), .Z(n406) );
  NAND2_X1 U477 ( .A1(n407), .A2(n406), .ZN(n408) );
  NAND2_X1 U478 ( .A1(n408), .A2(n552), .ZN(n413) );
  NOR2_X1 U479 ( .A1(n552), .A2(n409), .ZN(n533) );
  XNOR2_X1 U480 ( .A(KEYINPUT28), .B(n555), .ZN(n497) );
  NAND2_X1 U481 ( .A1(n533), .A2(n497), .ZN(n519) );
  XNOR2_X1 U482 ( .A(n519), .B(KEYINPUT101), .ZN(n411) );
  XNOR2_X1 U483 ( .A(n521), .B(KEYINPUT87), .ZN(n410) );
  NAND2_X1 U484 ( .A1(n411), .A2(n410), .ZN(n412) );
  NAND2_X1 U485 ( .A1(n413), .A2(n412), .ZN(n462) );
  NAND2_X1 U486 ( .A1(n585), .A2(n462), .ZN(n414) );
  XNOR2_X1 U487 ( .A(KEYINPUT106), .B(n414), .ZN(n415) );
  NOR2_X1 U488 ( .A1(n588), .A2(n415), .ZN(n418) );
  XOR2_X1 U489 ( .A(KEYINPUT77), .B(KEYINPUT31), .Z(n424) );
  XOR2_X1 U490 ( .A(KEYINPUT32), .B(KEYINPUT74), .Z(n420) );
  XNOR2_X1 U491 ( .A(KEYINPUT33), .B(KEYINPUT76), .ZN(n419) );
  XNOR2_X1 U492 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U493 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U494 ( .A(n424), .B(n423), .ZN(n430) );
  XOR2_X1 U495 ( .A(n426), .B(n425), .Z(n428) );
  NAND2_X1 U496 ( .A1(G230GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U497 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U498 ( .A(n430), .B(n429), .Z(n434) );
  XNOR2_X1 U499 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U500 ( .A(n434), .B(n433), .ZN(n582) );
  NAND2_X1 U501 ( .A1(n436), .A2(n435), .ZN(n440) );
  INV_X1 U502 ( .A(n435), .ZN(n438) );
  INV_X1 U503 ( .A(n436), .ZN(n437) );
  NAND2_X1 U504 ( .A1(n438), .A2(n437), .ZN(n439) );
  NAND2_X1 U505 ( .A1(n440), .A2(n439), .ZN(n442) );
  AND2_X1 U506 ( .A1(G229GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U507 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U508 ( .A(KEYINPUT67), .B(n443), .Z(n450) );
  XNOR2_X1 U509 ( .A(n444), .B(KEYINPUT29), .ZN(n448) );
  XOR2_X1 U510 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n446) );
  XNOR2_X1 U511 ( .A(G197GAT), .B(KEYINPUT72), .ZN(n445) );
  XNOR2_X1 U512 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(n537) );
  INV_X1 U514 ( .A(n537), .ZN(n578) );
  XNOR2_X1 U515 ( .A(n578), .B(KEYINPUT73), .ZN(n560) );
  NAND2_X1 U516 ( .A1(n582), .A2(n560), .ZN(n464) );
  NOR2_X1 U517 ( .A1(n491), .A2(n464), .ZN(n453) );
  XOR2_X1 U518 ( .A(KEYINPUT38), .B(n453), .Z(n454) );
  NOR2_X1 U519 ( .A1(n552), .A2(n478), .ZN(n458) );
  XNOR2_X1 U520 ( .A(KEYINPUT105), .B(KEYINPUT39), .ZN(n456) );
  XOR2_X1 U521 ( .A(KEYINPUT16), .B(KEYINPUT82), .Z(n461) );
  NAND2_X1 U522 ( .A1(n459), .A2(n567), .ZN(n460) );
  XNOR2_X1 U523 ( .A(n461), .B(n460), .ZN(n463) );
  NAND2_X1 U524 ( .A1(n463), .A2(n462), .ZN(n481) );
  NOR2_X1 U525 ( .A1(n481), .A2(n464), .ZN(n465) );
  XNOR2_X1 U526 ( .A(n465), .B(KEYINPUT103), .ZN(n472) );
  NOR2_X1 U527 ( .A1(n552), .A2(n472), .ZN(n467) );
  XNOR2_X1 U528 ( .A(KEYINPUT34), .B(KEYINPUT104), .ZN(n466) );
  XNOR2_X1 U529 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U530 ( .A(G1GAT), .B(n468), .Z(G1324GAT) );
  NOR2_X1 U531 ( .A1(n549), .A2(n472), .ZN(n469) );
  XOR2_X1 U532 ( .A(G8GAT), .B(n469), .Z(G1325GAT) );
  NOR2_X1 U533 ( .A1(n559), .A2(n472), .ZN(n471) );
  XNOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n470) );
  XNOR2_X1 U535 ( .A(n471), .B(n470), .ZN(G1326GAT) );
  NOR2_X1 U536 ( .A1(n497), .A2(n472), .ZN(n473) );
  XOR2_X1 U537 ( .A(G22GAT), .B(n473), .Z(G1327GAT) );
  NOR2_X1 U538 ( .A1(n549), .A2(n478), .ZN(n474) );
  XOR2_X1 U539 ( .A(G36GAT), .B(n474), .Z(G1329GAT) );
  NOR2_X1 U540 ( .A1(n559), .A2(n478), .ZN(n476) );
  XNOR2_X1 U541 ( .A(KEYINPUT40), .B(KEYINPUT109), .ZN(n475) );
  XNOR2_X1 U542 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U543 ( .A(G43GAT), .B(n477), .ZN(G1330GAT) );
  NOR2_X1 U544 ( .A1(n497), .A2(n478), .ZN(n479) );
  XOR2_X1 U545 ( .A(G50GAT), .B(n479), .Z(G1331GAT) );
  XNOR2_X1 U546 ( .A(n582), .B(KEYINPUT41), .ZN(n541) );
  XNOR2_X1 U547 ( .A(KEYINPUT110), .B(n541), .ZN(n562) );
  NAND2_X1 U548 ( .A1(n562), .A2(n578), .ZN(n480) );
  XOR2_X1 U549 ( .A(KEYINPUT111), .B(n480), .Z(n490) );
  OR2_X1 U550 ( .A1(n490), .A2(n481), .ZN(n486) );
  NOR2_X1 U551 ( .A1(n552), .A2(n486), .ZN(n482) );
  XOR2_X1 U552 ( .A(n482), .B(KEYINPUT42), .Z(n483) );
  XNOR2_X1 U553 ( .A(G57GAT), .B(n483), .ZN(G1332GAT) );
  NOR2_X1 U554 ( .A1(n549), .A2(n486), .ZN(n484) );
  XOR2_X1 U555 ( .A(G64GAT), .B(n484), .Z(G1333GAT) );
  NOR2_X1 U556 ( .A1(n559), .A2(n486), .ZN(n485) );
  XOR2_X1 U557 ( .A(G71GAT), .B(n485), .Z(G1334GAT) );
  NOR2_X1 U558 ( .A1(n497), .A2(n486), .ZN(n488) );
  XNOR2_X1 U559 ( .A(KEYINPUT112), .B(KEYINPUT43), .ZN(n487) );
  XNOR2_X1 U560 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U561 ( .A(G78GAT), .B(n489), .ZN(G1335GAT) );
  OR2_X1 U562 ( .A1(n491), .A2(n490), .ZN(n496) );
  NOR2_X1 U563 ( .A1(n552), .A2(n496), .ZN(n493) );
  XNOR2_X1 U564 ( .A(G85GAT), .B(KEYINPUT113), .ZN(n492) );
  XNOR2_X1 U565 ( .A(n493), .B(n492), .ZN(G1336GAT) );
  NOR2_X1 U566 ( .A1(n549), .A2(n496), .ZN(n494) );
  XOR2_X1 U567 ( .A(G92GAT), .B(n494), .Z(G1337GAT) );
  NOR2_X1 U568 ( .A1(n559), .A2(n496), .ZN(n495) );
  XOR2_X1 U569 ( .A(G99GAT), .B(n495), .Z(G1338GAT) );
  NOR2_X1 U570 ( .A1(n497), .A2(n496), .ZN(n499) );
  XNOR2_X1 U571 ( .A(KEYINPUT44), .B(KEYINPUT114), .ZN(n498) );
  XNOR2_X1 U572 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U573 ( .A(G106GAT), .B(n500), .Z(G1339GAT) );
  NAND2_X1 U574 ( .A1(n541), .A2(n537), .ZN(n502) );
  OR2_X1 U575 ( .A1(n505), .A2(n567), .ZN(n504) );
  INV_X1 U576 ( .A(KEYINPUT116), .ZN(n503) );
  NAND2_X1 U577 ( .A1(n504), .A2(n503), .ZN(n508) );
  NOR2_X1 U578 ( .A1(n505), .A2(n567), .ZN(n506) );
  NAND2_X1 U579 ( .A1(KEYINPUT116), .A2(n506), .ZN(n507) );
  NAND2_X1 U580 ( .A1(n508), .A2(n507), .ZN(n510) );
  NAND2_X1 U581 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U582 ( .A(n511), .B(KEYINPUT47), .ZN(n516) );
  NOR2_X1 U583 ( .A1(n585), .A2(n588), .ZN(n512) );
  XNOR2_X1 U584 ( .A(KEYINPUT45), .B(n512), .ZN(n513) );
  NAND2_X1 U585 ( .A1(n513), .A2(n582), .ZN(n514) );
  NOR2_X1 U586 ( .A1(n560), .A2(n514), .ZN(n515) );
  NOR2_X1 U587 ( .A1(n516), .A2(n515), .ZN(n518) );
  BUF_X1 U588 ( .A(n550), .Z(n534) );
  NOR2_X1 U589 ( .A1(n534), .A2(n519), .ZN(n520) );
  NAND2_X1 U590 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n522), .B(KEYINPUT117), .ZN(n529) );
  NAND2_X1 U592 ( .A1(n560), .A2(n529), .ZN(n523) );
  XNOR2_X1 U593 ( .A(n523), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(G120GAT), .B(KEYINPUT49), .Z(n525) );
  NAND2_X1 U595 ( .A1(n529), .A2(n562), .ZN(n524) );
  XNOR2_X1 U596 ( .A(n525), .B(n524), .ZN(G1341GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n527) );
  NAND2_X1 U598 ( .A1(n529), .A2(n567), .ZN(n526) );
  XNOR2_X1 U599 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U600 ( .A(G127GAT), .B(n528), .Z(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n531) );
  NAND2_X1 U602 ( .A1(n529), .A2(n571), .ZN(n530) );
  XNOR2_X1 U603 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U604 ( .A(G134GAT), .B(n532), .Z(G1343GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n539) );
  NAND2_X1 U606 ( .A1(n533), .A2(n576), .ZN(n535) );
  NOR2_X1 U607 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U608 ( .A(n536), .B(KEYINPUT120), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n547), .A2(n537), .ZN(n538) );
  XNOR2_X1 U610 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(n540), .ZN(G1344GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n543) );
  NAND2_X1 U613 ( .A1(n547), .A2(n541), .ZN(n542) );
  XNOR2_X1 U614 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(n544), .ZN(G1345GAT) );
  NAND2_X1 U616 ( .A1(n547), .A2(n567), .ZN(n545) );
  XNOR2_X1 U617 ( .A(n545), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U618 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U619 ( .A(n548), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U620 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U621 ( .A(n551), .B(KEYINPUT54), .ZN(n553) );
  NAND2_X1 U622 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n554), .B(KEYINPUT65), .ZN(n577) );
  NAND2_X1 U624 ( .A1(n577), .A2(n555), .ZN(n557) );
  INV_X1 U625 ( .A(KEYINPUT55), .ZN(n556) );
  XNOR2_X1 U626 ( .A(n557), .B(n556), .ZN(n558) );
  NAND2_X1 U627 ( .A1(n560), .A2(n570), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U629 ( .A1(n562), .A2(n570), .ZN(n564) );
  XOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT123), .Z(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n566) );
  XOR2_X1 U632 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  NAND2_X1 U634 ( .A1(n567), .A2(n570), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(KEYINPUT124), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(G183GAT), .ZN(G1350GAT) );
  AND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n575) );
  XNOR2_X1 U638 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n572), .B(KEYINPUT125), .ZN(n573) );
  XNOR2_X1 U640 ( .A(KEYINPUT126), .B(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1351GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n587) );
  NOR2_X1 U643 ( .A1(n578), .A2(n587), .ZN(n580) );
  XNOR2_X1 U644 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(n581), .ZN(G1352GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n587), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n587), .ZN(n586) );
  XOR2_X1 U651 ( .A(G211GAT), .B(n586), .Z(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U653 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

