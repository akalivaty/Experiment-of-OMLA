//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  OAI21_X1  g004(.A(G128), .B1(new_n188), .B2(new_n190), .ZN(new_n191));
  OR3_X1    g005(.A1(new_n189), .A2(KEYINPUT65), .A3(G146), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT65), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n189), .A2(G146), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n198), .B(KEYINPUT68), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(new_n196), .A3(G128), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(new_n188), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT11), .B1(new_n204), .B2(G134), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G137), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n207), .A2(new_n208), .A3(new_n209), .A4(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT11), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(new_n210), .B2(G137), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n214), .A2(new_n215), .A3(new_n209), .A4(new_n211), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT66), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n210), .A2(G137), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n209), .B1(new_n220), .B2(new_n211), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n203), .A2(new_n218), .A3(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(G116), .B(G119), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT2), .B(G113), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n224), .B(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n214), .A2(new_n211), .A3(new_n215), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G131), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n216), .A2(KEYINPUT66), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n216), .A2(KEYINPUT66), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT69), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n235), .B(new_n230), .C1(new_n231), .C2(new_n232), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  XOR2_X1   g051(.A(KEYINPUT0), .B(G128), .Z(new_n238));
  AOI22_X1  g052(.A1(new_n197), .A2(new_n238), .B1(new_n201), .B2(KEYINPUT0), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n228), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n239), .ZN(new_n241));
  AOI211_X1 g055(.A(KEYINPUT70), .B(new_n241), .C1(new_n234), .C2(new_n236), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n227), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n243), .A2(new_n246), .A3(KEYINPUT30), .A4(new_n223), .ZN(new_n247));
  INV_X1    g061(.A(new_n236), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n235), .B1(new_n218), .B2(new_n230), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n239), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT70), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n237), .A2(new_n228), .A3(new_n239), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n251), .A2(KEYINPUT30), .A3(new_n223), .A4(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT71), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n247), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n233), .A2(new_n239), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n223), .A2(new_n256), .ZN(new_n257));
  XOR2_X1   g071(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n226), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n245), .B1(new_n255), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G210), .ZN(new_n264));
  NOR3_X1   g078(.A1(new_n264), .A2(G237), .A3(G953), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(G101), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n267));
  XOR2_X1   g081(.A(new_n266), .B(new_n267), .Z(new_n268));
  OAI21_X1  g082(.A(new_n187), .B1(new_n263), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n268), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n261), .B1(new_n254), .B2(new_n247), .ZN(new_n271));
  OAI211_X1 g085(.A(KEYINPUT72), .B(new_n270), .C1(new_n271), .C2(new_n245), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT28), .B1(new_n227), .B2(new_n250), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n257), .A2(new_n260), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n244), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n273), .B1(new_n275), .B2(KEYINPUT28), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT29), .B1(new_n276), .B2(new_n268), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n269), .A2(new_n272), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT73), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n244), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n243), .A2(new_n223), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n282), .A2(new_n260), .B1(new_n227), .B2(new_n243), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n281), .B1(new_n283), .B2(new_n280), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n273), .B1(new_n284), .B2(KEYINPUT28), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n268), .A2(KEYINPUT29), .ZN(new_n286));
  AOI21_X1  g100(.A(G902), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n269), .A2(new_n277), .A3(new_n288), .A4(new_n272), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n279), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G472), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n276), .A2(new_n268), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n255), .A2(new_n262), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n244), .A3(new_n268), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT31), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n263), .A2(KEYINPUT31), .A3(new_n268), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n292), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(G472), .A2(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT32), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT31), .B1(new_n263), .B2(new_n268), .ZN(new_n302));
  NOR4_X1   g116(.A1(new_n271), .A2(new_n295), .A3(new_n245), .A4(new_n270), .ZN(new_n303));
  OAI22_X1  g117(.A1(new_n302), .A2(new_n303), .B1(new_n276), .B2(new_n268), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT32), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(new_n299), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n291), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT75), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n291), .A2(new_n310), .A3(new_n307), .ZN(new_n311));
  XNOR2_X1  g125(.A(G125), .B(G140), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n312), .A2(new_n193), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G140), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT16), .B1(new_n315), .B2(G125), .ZN(new_n316));
  NAND2_X1  g130(.A1(KEYINPUT77), .A2(G125), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(G140), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n316), .B1(new_n318), .B2(KEYINPUT16), .ZN(new_n319));
  OR2_X1    g133(.A1(new_n319), .A2(new_n193), .ZN(new_n320));
  INV_X1    g134(.A(G128), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G119), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(KEYINPUT23), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n321), .A2(G119), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(G110), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n327), .B(KEYINPUT79), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n322), .ZN(new_n329));
  XOR2_X1   g143(.A(new_n329), .B(KEYINPUT76), .Z(new_n330));
  XOR2_X1   g144(.A(KEYINPUT24), .B(G110), .Z(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n314), .B(new_n320), .C1(new_n328), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n320), .A2(KEYINPUT78), .ZN(new_n334));
  OR3_X1    g148(.A1(new_n319), .A2(KEYINPUT78), .A3(new_n193), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n319), .A2(new_n193), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n330), .A2(new_n331), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n326), .A2(G110), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT22), .B(G137), .ZN(new_n342));
  INV_X1    g156(.A(G953), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n343), .A2(G221), .A3(G234), .ZN(new_n344));
  XOR2_X1   g158(.A(new_n342), .B(new_n344), .Z(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n345), .B1(new_n333), .B2(new_n340), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G902), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(KEYINPUT80), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n349), .B(new_n350), .C1(new_n354), .C2(KEYINPUT25), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G217), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(G234), .B2(new_n350), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n358), .A2(G902), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n349), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G221), .ZN(new_n365));
  XOR2_X1   g179(.A(KEYINPUT9), .B(G234), .Z(new_n366));
  AOI21_X1  g180(.A(new_n365), .B1(new_n366), .B2(new_n350), .ZN(new_n367));
  XNOR2_X1  g181(.A(G110), .B(G140), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n343), .A2(G227), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G104), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT3), .B1(new_n371), .B2(G107), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n373));
  INV_X1    g187(.A(G107), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(G104), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n372), .B(new_n375), .C1(G104), .C2(new_n374), .ZN(new_n376));
  OR2_X1    g190(.A1(new_n376), .A2(G101), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n374), .A2(G104), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n371), .A2(G107), .ZN(new_n379));
  OAI21_X1  g193(.A(G101), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n202), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n383));
  OR2_X1    g197(.A1(new_n383), .A2(KEYINPUT82), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n321), .B1(new_n383), .B2(KEYINPUT82), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n384), .A2(new_n385), .B1(new_n194), .B2(new_n196), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n381), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n387), .B1(new_n203), .B2(new_n381), .ZN(new_n388));
  XOR2_X1   g202(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n233), .A3(new_n389), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n388), .A2(new_n237), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n390), .B1(new_n391), .B2(KEYINPUT12), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n376), .A2(G101), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n377), .A2(KEYINPUT4), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n376), .A2(new_n395), .A3(G101), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n239), .A3(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(KEYINPUT81), .ZN(new_n398));
  INV_X1    g212(.A(new_n237), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT10), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n387), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n203), .A2(KEYINPUT10), .A3(new_n381), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n398), .A2(new_n399), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n370), .B1(new_n392), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n398), .A2(new_n401), .A3(new_n402), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n405), .A2(new_n237), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n370), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G469), .B1(new_n409), .B2(G902), .ZN(new_n410));
  INV_X1    g224(.A(new_n370), .ZN(new_n411));
  INV_X1    g225(.A(new_n403), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n411), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n390), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT12), .B1(new_n388), .B2(new_n237), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n413), .B1(new_n407), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G469), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n418), .A3(new_n350), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n367), .B1(new_n410), .B2(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n309), .A2(new_n311), .A3(new_n364), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n343), .A2(G952), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(G234), .B2(G237), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  XOR2_X1   g238(.A(KEYINPUT21), .B(G898), .Z(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT95), .ZN(new_n426));
  AOI211_X1 g240(.A(new_n350), .B(new_n343), .C1(G234), .C2(G237), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n424), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G214), .B1(G237), .B2(G902), .ZN(new_n430));
  XOR2_X1   g244(.A(KEYINPUT84), .B(KEYINPUT5), .Z(new_n431));
  INV_X1    g245(.A(G119), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(G116), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT85), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n431), .A2(KEYINPUT85), .A3(G116), .A4(new_n432), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n436), .A3(G113), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT88), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n224), .A2(KEYINPUT5), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n437), .A2(new_n438), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n224), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n443), .A2(new_n225), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT89), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n442), .A2(new_n447), .A3(new_n444), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n446), .A2(new_n381), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n443), .A2(new_n431), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n437), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n381), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n444), .ZN(new_n453));
  XOR2_X1   g267(.A(G110), .B(G122), .Z(new_n454));
  XOR2_X1   g268(.A(new_n454), .B(KEYINPUT8), .Z(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT90), .B1(new_n449), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G125), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n199), .A2(KEYINPUT87), .A3(new_n458), .A4(new_n202), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT87), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n203), .B2(G125), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n459), .B(new_n461), .C1(new_n458), .C2(new_n239), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT7), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n343), .A2(G224), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n462), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n451), .A2(new_n381), .A3(new_n444), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n394), .A2(new_n260), .A3(new_n396), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(new_n454), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n462), .A2(new_n465), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n470), .B1(new_n471), .B2(KEYINPUT7), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n446), .A2(new_n381), .A3(new_n448), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT90), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n473), .A2(new_n474), .A3(new_n455), .A4(new_n453), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n457), .A2(new_n466), .A3(new_n472), .A4(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G210), .B1(G237), .B2(G902), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n462), .B(new_n465), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n469), .A2(new_n454), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n479), .B1(KEYINPUT86), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n470), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n480), .A2(KEYINPUT86), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n469), .A2(new_n454), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(G902), .B1(new_n478), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n476), .A2(new_n477), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n477), .B1(new_n476), .B2(new_n486), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n429), .B(new_n430), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G237), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n343), .A3(G214), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(G143), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(new_n209), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT17), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n493), .B(new_n209), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n495), .B1(new_n496), .B2(KEYINPUT17), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n337), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n313), .B1(G146), .B2(new_n318), .ZN(new_n499));
  INV_X1    g313(.A(new_n493), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(KEYINPUT18), .B2(G131), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n494), .A2(KEYINPUT18), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT91), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n494), .A2(KEYINPUT91), .A3(KEYINPUT18), .ZN(new_n505));
  AOI211_X1 g319(.A(new_n499), .B(new_n501), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n498), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G113), .B(G122), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT93), .B(G104), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n496), .A2(new_n320), .ZN(new_n513));
  XOR2_X1   g327(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n514));
  AOI22_X1  g328(.A1(new_n318), .A2(KEYINPUT19), .B1(new_n514), .B2(new_n312), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n513), .B1(new_n193), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n510), .B1(new_n506), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G475), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n519), .A3(new_n350), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT20), .ZN(new_n521));
  OR2_X1    g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n507), .B(new_n510), .ZN(new_n523));
  OAI21_X1  g337(.A(G475), .B1(new_n523), .B2(G902), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n520), .A2(new_n521), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(G128), .B(G143), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n210), .B1(new_n528), .B2(KEYINPUT13), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n189), .A2(G128), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n529), .B1(KEYINPUT13), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(G116), .B(G122), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(new_n374), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n528), .A2(new_n210), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n528), .B(new_n210), .ZN(new_n536));
  INV_X1    g350(.A(G116), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT14), .A3(G122), .ZN(new_n538));
  INV_X1    g352(.A(new_n532), .ZN(new_n539));
  OAI211_X1 g353(.A(G107), .B(new_n538), .C1(new_n539), .C2(KEYINPUT14), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n532), .A2(new_n374), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT94), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n535), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n366), .A2(G217), .A3(new_n343), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n350), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT15), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G478), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n547), .B(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n527), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n490), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n421), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT96), .B(G101), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(G3));
  XOR2_X1   g370(.A(new_n546), .B(KEYINPUT33), .Z(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G478), .ZN(new_n558));
  NAND2_X1  g372(.A1(G478), .A2(G902), .ZN(new_n559));
  OR2_X1    g373(.A1(new_n547), .A2(G478), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n526), .A2(new_n562), .ZN(new_n563));
  OR3_X1    g377(.A1(new_n490), .A2(KEYINPUT97), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT97), .B1(new_n490), .B2(new_n563), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G472), .B1(new_n298), .B2(G902), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n304), .A2(new_n299), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n364), .A2(new_n567), .A3(new_n568), .A4(new_n420), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT34), .B(G104), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n570), .B(new_n571), .ZN(G6));
  INV_X1    g386(.A(new_n550), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n527), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n490), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT98), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(new_n569), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT35), .B(G107), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(G9));
  XOR2_X1   g393(.A(new_n341), .B(KEYINPUT99), .Z(new_n580));
  NOR2_X1   g394(.A1(new_n346), .A2(KEYINPUT36), .ZN(new_n581));
  OR2_X1    g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n581), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n361), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n359), .A2(new_n584), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n585), .A2(new_n420), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n552), .A2(new_n568), .A3(new_n567), .A4(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT37), .B(G110), .Z(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(G12));
  INV_X1    g403(.A(new_n430), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n476), .A2(new_n486), .ZN(new_n591));
  INV_X1    g405(.A(new_n477), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n590), .B1(new_n593), .B2(new_n487), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n594), .A2(new_n420), .ZN(new_n595));
  INV_X1    g409(.A(G900), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n427), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n424), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n574), .A2(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n309), .A2(new_n311), .A3(new_n585), .A4(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G128), .ZN(G30));
  OAI21_X1  g417(.A(new_n350), .B1(new_n284), .B2(new_n268), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n263), .A2(new_n270), .ZN(new_n605));
  OAI21_X1  g419(.A(G472), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n585), .B1(new_n307), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n593), .A2(new_n487), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(KEYINPUT38), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n526), .A2(new_n573), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n610), .A2(new_n590), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n607), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  XOR2_X1   g429(.A(new_n598), .B(KEYINPUT39), .Z(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n420), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n618), .B(KEYINPUT101), .Z(new_n619));
  OR2_X1    g433(.A1(new_n619), .A2(KEYINPUT40), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(KEYINPUT40), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n614), .A2(new_n615), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT102), .B(G143), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G45));
  INV_X1    g438(.A(new_n311), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n310), .B1(new_n291), .B2(new_n307), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n563), .A2(new_n599), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n627), .A2(new_n585), .A3(new_n595), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G146), .ZN(G48));
  NAND2_X1  g444(.A1(new_n417), .A2(new_n350), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(G469), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n419), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(new_n367), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n309), .A2(new_n311), .A3(new_n364), .A4(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n566), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT41), .B(G113), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G15));
  OR2_X1    g452(.A1(new_n635), .A2(new_n576), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G116), .ZN(G18));
  NAND4_X1  g454(.A1(new_n309), .A2(new_n552), .A3(new_n311), .A4(new_n585), .ZN(new_n641));
  INV_X1    g455(.A(new_n634), .ZN(new_n642));
  OR2_X1    g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G119), .ZN(G21));
  AND3_X1   g458(.A1(new_n359), .A2(KEYINPUT103), .A3(new_n362), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT103), .B1(new_n359), .B2(new_n362), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI22_X1  g461(.A1(new_n302), .A2(new_n303), .B1(new_n285), .B2(new_n268), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n299), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n647), .A2(new_n567), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n490), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n642), .A2(new_n610), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G122), .ZN(G24));
  NAND4_X1  g468(.A1(new_n567), .A2(new_n628), .A3(new_n649), .A4(new_n585), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n634), .A2(new_n594), .ZN(new_n656));
  OR3_X1    g470(.A1(new_n655), .A2(new_n656), .A3(KEYINPUT104), .ZN(new_n657));
  OAI21_X1  g471(.A(KEYINPUT104), .B1(new_n655), .B2(new_n656), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G125), .ZN(G27));
  NOR2_X1   g474(.A1(new_n608), .A2(new_n590), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n309), .A2(new_n311), .A3(new_n364), .A4(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n628), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n410), .A2(new_n419), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n664), .A2(KEYINPUT105), .ZN(new_n665));
  INV_X1    g479(.A(new_n367), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n664), .A2(KEYINPUT105), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n662), .A2(new_n663), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n661), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n663), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n671), .A2(new_n673), .A3(new_n308), .A4(new_n647), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  OAI22_X1  g491(.A1(new_n669), .A2(KEYINPUT42), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G131), .ZN(G33));
  NOR2_X1   g493(.A1(new_n662), .A2(new_n668), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n680), .A2(new_n600), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n210), .ZN(G36));
  NAND2_X1  g496(.A1(new_n567), .A2(new_n568), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n585), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n527), .A2(new_n562), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT43), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n684), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n672), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n687), .B1(new_n684), .B2(new_n686), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n411), .B1(new_n416), .B2(new_n412), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n691), .B(KEYINPUT45), .C1(new_n406), .C2(new_n407), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(new_n404), .B2(new_n408), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n692), .A2(new_n694), .A3(G469), .ZN(new_n695));
  NAND2_X1  g509(.A1(G469), .A2(G902), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT46), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n419), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n697), .A2(new_n698), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n666), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n616), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n689), .A2(new_n690), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G137), .ZN(G39));
  XNOR2_X1  g519(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n702), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n309), .A2(new_n311), .ZN(new_n708));
  INV_X1    g522(.A(new_n364), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n707), .A2(new_n708), .A3(new_n709), .A4(new_n673), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G140), .ZN(G42));
  OR2_X1    g525(.A1(G952), .A2(G953), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n713));
  AND4_X1   g527(.A1(new_n309), .A2(new_n311), .A3(new_n364), .A4(new_n634), .ZN(new_n714));
  INV_X1    g528(.A(new_n566), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(new_n639), .A3(new_n643), .A4(KEYINPUT111), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n574), .A2(new_n563), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n651), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n587), .B1(new_n569), .B2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n721), .B1(new_n421), .B2(new_n553), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n721), .B(KEYINPUT109), .C1(new_n421), .C2(new_n553), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n727));
  OAI22_X1  g541(.A1(new_n576), .A2(new_n635), .B1(new_n641), .B2(new_n642), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n653), .B1(new_n635), .B2(new_n566), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AND4_X1   g544(.A1(KEYINPUT53), .A2(new_n717), .A3(new_n726), .A4(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n309), .A2(new_n311), .A3(new_n585), .A4(new_n595), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n659), .B(new_n602), .C1(new_n732), .C2(new_n663), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n611), .A2(new_n608), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n668), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n607), .A3(new_n598), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT52), .B1(new_n733), .B2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n586), .A2(new_n550), .A3(new_n527), .A4(new_n598), .ZN(new_n739));
  OAI22_X1  g553(.A1(new_n708), .A2(new_n739), .B1(new_n655), .B2(new_n668), .ZN(new_n740));
  AOI22_X1  g554(.A1(new_n680), .A2(new_n600), .B1(new_n740), .B2(new_n661), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n659), .A2(new_n602), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n742), .A2(new_n629), .A3(new_n743), .A4(new_n736), .ZN(new_n744));
  AND4_X1   g558(.A1(new_n678), .A2(new_n738), .A3(new_n741), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n731), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n678), .A2(new_n738), .A3(new_n741), .A4(new_n744), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n728), .A2(new_n729), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n726), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n748), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n746), .A2(new_n747), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(KEYINPUT110), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n745), .A2(KEYINPUT53), .A3(new_n726), .A4(new_n750), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n756), .B(new_n748), .C1(new_n749), .C2(new_n751), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n753), .B1(new_n758), .B2(KEYINPUT54), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n686), .A2(new_n424), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n672), .A2(new_n642), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI211_X1 g576(.A(new_n646), .B(new_n645), .C1(new_n291), .C2(new_n307), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g578(.A(new_n764), .B(KEYINPUT48), .Z(new_n765));
  NAND2_X1  g579(.A1(new_n307), .A2(new_n606), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n767), .A2(new_n761), .A3(new_n423), .A4(new_n364), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n563), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n765), .A2(new_n422), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n633), .B(KEYINPUT108), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT112), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n666), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n773), .A2(new_n707), .ZN(new_n774));
  XOR2_X1   g588(.A(new_n774), .B(KEYINPUT114), .Z(new_n775));
  NAND2_X1  g589(.A1(new_n760), .A2(new_n650), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n672), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT51), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n776), .A2(new_n430), .A3(new_n609), .A4(new_n642), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT50), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n762), .A2(new_n567), .A3(new_n585), .A4(new_n649), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT113), .ZN(new_n783));
  INV_X1    g597(.A(new_n768), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n527), .A3(new_n561), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n781), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n770), .B1(new_n779), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n786), .B1(new_n777), .B2(new_n774), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(KEYINPUT51), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n759), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n776), .A2(new_n656), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n712), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n771), .B(KEYINPUT49), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n685), .A2(new_n590), .A3(new_n367), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n647), .A3(new_n795), .ZN(new_n796));
  OR3_X1    g610(.A1(new_n796), .A2(new_n766), .A3(new_n609), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n793), .A2(new_n797), .ZN(G75));
  INV_X1    g612(.A(new_n485), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(new_n478), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT55), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT56), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n801), .B1(KEYINPUT115), .B2(new_n802), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n264), .B(new_n350), .C1(new_n746), .C2(new_n752), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n803), .B1(new_n804), .B2(KEYINPUT56), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n343), .A2(G952), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n746), .A2(new_n752), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(G210), .A3(G902), .ZN(new_n809));
  INV_X1    g623(.A(new_n803), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n802), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n805), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n805), .A2(KEYINPUT116), .A3(new_n811), .A4(new_n807), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(G51));
  AOI21_X1  g630(.A(new_n747), .B1(new_n746), .B2(new_n752), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n753), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n696), .B(KEYINPUT57), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n417), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n808), .ZN(new_n821));
  OR3_X1    g635(.A1(new_n821), .A2(new_n350), .A3(new_n695), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n806), .B1(new_n820), .B2(new_n822), .ZN(G54));
  NOR2_X1   g637(.A1(new_n821), .A2(new_n350), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(KEYINPUT58), .A3(G475), .ZN(new_n825));
  INV_X1    g639(.A(new_n518), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n824), .A2(KEYINPUT58), .A3(G475), .A4(new_n518), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n827), .A2(new_n807), .A3(new_n828), .ZN(G60));
  XNOR2_X1  g643(.A(new_n559), .B(KEYINPUT59), .ZN(new_n830));
  XOR2_X1   g644(.A(KEYINPUT117), .B(KEYINPUT118), .Z(new_n831));
  XOR2_X1   g645(.A(new_n830), .B(new_n831), .Z(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n557), .B1(new_n759), .B2(new_n833), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n557), .A2(new_n833), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n808), .A2(KEYINPUT54), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n746), .A2(new_n747), .A3(new_n752), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT119), .B1(new_n838), .B2(new_n806), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n840), .B(new_n807), .C1(new_n818), .C2(new_n835), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n834), .A2(new_n839), .A3(new_n841), .ZN(G63));
  AND2_X1   g656(.A1(new_n582), .A2(new_n583), .ZN(new_n843));
  NAND2_X1  g657(.A1(G217), .A2(G902), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT60), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n808), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n807), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(KEYINPUT120), .A2(KEYINPUT61), .ZN(new_n850));
  OR2_X1    g664(.A1(KEYINPUT120), .A2(KEYINPUT61), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n349), .B1(new_n808), .B2(new_n846), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(KEYINPUT120), .B(KEYINPUT61), .C1(new_n848), .C2(new_n852), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(G66));
  AOI21_X1  g670(.A(new_n343), .B1(new_n426), .B2(G224), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n751), .B2(new_n343), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n799), .B1(G898), .B2(new_n343), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n858), .B(new_n859), .Z(G69));
  NAND2_X1  g674(.A1(new_n255), .A2(new_n259), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n861), .B(new_n515), .Z(new_n862));
  AOI21_X1  g676(.A(new_n343), .B1(G227), .B2(G900), .ZN(new_n863));
  XOR2_X1   g677(.A(KEYINPUT121), .B(KEYINPUT62), .Z(new_n864));
  OR3_X1    g678(.A1(new_n622), .A2(new_n733), .A3(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n704), .A2(new_n710), .ZN(new_n866));
  INV_X1    g680(.A(new_n662), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n619), .A3(new_n718), .ZN(new_n868));
  OAI22_X1  g682(.A1(new_n622), .A2(new_n733), .B1(KEYINPUT121), .B2(KEYINPUT62), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n865), .A2(new_n866), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  AOI211_X1 g684(.A(new_n862), .B(new_n863), .C1(new_n870), .C2(new_n343), .ZN(new_n871));
  INV_X1    g685(.A(new_n734), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n763), .A2(new_n703), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  AND4_X1   g690(.A1(new_n704), .A2(new_n875), .A3(new_n710), .A4(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n681), .A2(new_n733), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n878), .A3(new_n678), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n879), .A2(G953), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n880), .A2(new_n862), .ZN(new_n881));
  OAI21_X1  g695(.A(G953), .B1(new_n596), .B2(G227), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n871), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT123), .ZN(G72));
  INV_X1    g698(.A(KEYINPUT127), .ZN(new_n885));
  XOR2_X1   g699(.A(KEYINPUT124), .B(KEYINPUT63), .Z(new_n886));
  NAND2_X1  g700(.A1(G472), .A2(G902), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n886), .B(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(new_n879), .B2(new_n751), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n889), .A2(new_n270), .A3(new_n263), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n890), .A2(new_n891), .A3(new_n807), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n891), .B1(new_n890), .B2(new_n807), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n269), .A2(new_n294), .A3(new_n272), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n758), .A2(new_n888), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n888), .B1(new_n870), .B2(new_n751), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT125), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n899), .B(new_n888), .C1(new_n870), .C2(new_n751), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n898), .A2(new_n605), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n885), .B1(new_n894), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n890), .A2(new_n807), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT126), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n890), .A2(new_n891), .A3(new_n807), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n907), .A2(KEYINPUT127), .A3(new_n896), .A4(new_n901), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n903), .A2(new_n908), .ZN(G57));
endmodule


