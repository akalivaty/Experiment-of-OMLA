//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT9), .ZN(new_n203));
  INV_X1    g002(.A(G71gat), .ZN(new_n204));
  INV_X1    g003(.A(G78gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G71gat), .B(G78gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n202), .A2(new_n208), .A3(new_n206), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n210), .A2(KEYINPUT95), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT95), .B1(new_n210), .B2(new_n211), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT21), .ZN(new_n216));
  INV_X1    g015(.A(G127gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(G127gat), .B1(new_n214), .B2(KEYINPUT21), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G15gat), .B(G22gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT16), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(G1gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(G1gat), .B2(new_n221), .ZN(new_n224));
  XOR2_X1   g023(.A(new_n224), .B(G8gat), .Z(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(new_n215), .B2(new_n216), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n220), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n219), .A3(new_n218), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n231));
  XNOR2_X1  g030(.A(G155gat), .B(G183gat), .ZN(new_n232));
  XOR2_X1   g031(.A(new_n231), .B(new_n232), .Z(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G231gat), .A2(G233gat), .ZN(new_n236));
  INV_X1    g035(.A(G211gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n230), .A2(new_n233), .ZN(new_n240));
  OR3_X1    g039(.A1(new_n235), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n239), .B1(new_n235), .B2(new_n240), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G85gat), .A2(G92gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT7), .ZN(new_n245));
  NAND2_X1  g044(.A1(G99gat), .A2(G106gat), .ZN(new_n246));
  INV_X1    g045(.A(G85gat), .ZN(new_n247));
  INV_X1    g046(.A(G92gat), .ZN(new_n248));
  AOI22_X1  g047(.A1(KEYINPUT8), .A2(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n245), .A2(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(G99gat), .B(G106gat), .Z(new_n251));
  AND3_X1   g050(.A1(new_n250), .A2(KEYINPUT96), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT96), .B1(new_n250), .B2(new_n251), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n250), .A2(new_n251), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G43gat), .B(G50gat), .ZN(new_n256));
  INV_X1    g055(.A(G29gat), .ZN(new_n257));
  INV_X1    g056(.A(G36gat), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT14), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n258), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT14), .B1(new_n257), .B2(new_n258), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n262), .A2(KEYINPUT15), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(KEYINPUT15), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n256), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(KEYINPUT15), .ZN(new_n266));
  INV_X1    g065(.A(new_n256), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n255), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n265), .A2(new_n268), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT93), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT17), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(KEYINPUT93), .A2(KEYINPUT17), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n273), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n265), .A2(new_n268), .A3(new_n275), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n269), .B(new_n270), .C1(new_n279), .C2(new_n255), .ZN(new_n280));
  XNOR2_X1  g079(.A(G190gat), .B(G218gat), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n280), .A2(new_n281), .ZN(new_n283));
  XNOR2_X1  g082(.A(G134gat), .B(G162gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT97), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  OR3_X1    g087(.A1(new_n282), .A2(new_n283), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n288), .B1(new_n282), .B2(new_n283), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT98), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n243), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n241), .A2(new_n242), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT98), .B1(new_n295), .B2(new_n291), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G197gat), .B(G204gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT22), .ZN(new_n299));
  NAND2_X1  g098(.A1(G211gat), .A2(G218gat), .ZN(new_n300));
  INV_X1    g099(.A(G218gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n237), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT79), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT22), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n300), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(new_n298), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT79), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n299), .A2(new_n308), .A3(new_n300), .A4(new_n302), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n304), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT80), .ZN(new_n312));
  NAND2_X1  g111(.A1(G226gat), .A2(G233gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT69), .ZN(new_n314));
  OR2_X1    g113(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n315), .A2(KEYINPUT27), .A3(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(G190gat), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n321));
  OAI21_X1  g120(.A(new_n314), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n321), .ZN(new_n323));
  AND2_X1   g122(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n318), .B1(new_n326), .B2(KEYINPUT27), .ZN(new_n327));
  OAI211_X1 g126(.A(KEYINPUT69), .B(new_n323), .C1(new_n327), .C2(G190gat), .ZN(new_n328));
  INV_X1    g127(.A(G190gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n319), .A2(KEYINPUT70), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT70), .B1(new_n319), .B2(new_n330), .ZN(new_n332));
  OAI211_X1 g131(.A(KEYINPUT28), .B(new_n329), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n322), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n335), .A2(KEYINPUT71), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT26), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G169gat), .ZN(new_n339));
  INV_X1    g138(.A(G176gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n341), .B1(new_n336), .B2(new_n337), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n338), .A2(new_n342), .B1(G183gat), .B2(G190gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT24), .ZN(new_n344));
  INV_X1    g143(.A(G183gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n344), .B1(new_n345), .B2(new_n329), .ZN(new_n346));
  NAND3_X1  g145(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT67), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n315), .A2(new_n316), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(new_n329), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n349), .B(new_n329), .C1(new_n324), .C2(new_n325), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n348), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n335), .A2(KEYINPUT23), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n355), .A2(new_n341), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n335), .A2(KEYINPUT23), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n354), .A2(KEYINPUT25), .A3(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(KEYINPUT65), .B(G176gat), .Z(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(KEYINPUT23), .A3(new_n339), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n346), .B(new_n347), .C1(G183gat), .C2(G190gat), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n356), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT25), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n334), .A2(new_n343), .B1(new_n359), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n313), .B1(new_n366), .B2(KEYINPUT29), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n334), .A2(new_n343), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n359), .A2(new_n365), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n313), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n312), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT80), .B1(new_n375), .B2(new_n313), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n311), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT88), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n313), .B1(new_n368), .B2(new_n369), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n380), .B1(new_n375), .B2(new_n313), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n310), .ZN(new_n382));
  OAI211_X1 g181(.A(KEYINPUT88), .B(new_n311), .C1(new_n373), .C2(new_n376), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n379), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT37), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT89), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  XOR2_X1   g186(.A(G8gat), .B(G36gat), .Z(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(G64gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(new_n248), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n310), .B1(new_n373), .B2(new_n376), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n367), .A2(new_n311), .A3(new_n372), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT37), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n391), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT38), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT89), .A3(KEYINPUT37), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n387), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT90), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT5), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT73), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT1), .ZN(new_n405));
  INV_X1    g204(.A(G113gat), .ZN(new_n406));
  INV_X1    g205(.A(G120gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT72), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT72), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(G120gat), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n406), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n407), .A2(G113gat), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n404), .B(new_n405), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G127gat), .B(G134gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(G113gat), .B(G120gat), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n414), .A2(new_n415), .A3(KEYINPUT1), .ZN(new_n416));
  OAI211_X1 g215(.A(KEYINPUT73), .B(new_n405), .C1(new_n411), .C2(new_n412), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n413), .A2(new_n416), .B1(new_n417), .B2(new_n414), .ZN(new_n418));
  INV_X1    g217(.A(G155gat), .ZN(new_n419));
  INV_X1    g218(.A(G162gat), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT83), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G141gat), .ZN(new_n422));
  INV_X1    g221(.A(G148gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G141gat), .A2(G148gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT2), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n427), .B1(G155gat), .B2(G162gat), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n421), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G155gat), .B(G162gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT2), .B1(new_n419), .B2(new_n420), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(new_n424), .A3(new_n425), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n430), .B1(new_n434), .B2(new_n421), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT3), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT84), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n429), .A2(new_n431), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n434), .A2(new_n430), .A3(new_n421), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT3), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n438), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI211_X1 g242(.A(KEYINPUT84), .B(KEYINPUT3), .C1(new_n439), .C2(new_n440), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n418), .B(new_n437), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT4), .B1(new_n418), .B2(new_n436), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n413), .A2(new_n416), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n417), .A2(new_n414), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT4), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n450), .A3(new_n441), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(G225gat), .A2(G233gat), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n445), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n453), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n449), .A2(new_n441), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n418), .A2(new_n436), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n403), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n461));
  XNOR2_X1  g260(.A(G1gat), .B(G29gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G57gat), .B(G85gat), .ZN(new_n464));
  XOR2_X1   g263(.A(new_n463), .B(new_n464), .Z(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n454), .A2(new_n403), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n460), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n467), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n465), .B1(new_n469), .B2(new_n459), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n460), .A2(KEYINPUT6), .A3(new_n466), .A4(new_n467), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n367), .A2(new_n312), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(new_n381), .B2(new_n312), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n393), .B1(new_n476), .B2(new_n310), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT37), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n398), .B1(new_n397), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT91), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n474), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n390), .B1(new_n392), .B2(new_n394), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(new_n479), .B2(KEYINPUT91), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT90), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n387), .A2(new_n399), .A3(new_n485), .A4(new_n400), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n402), .A2(new_n482), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  XOR2_X1   g286(.A(G78gat), .B(G106gat), .Z(new_n488));
  OAI21_X1  g287(.A(new_n442), .B1(new_n432), .B2(new_n435), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT84), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n441), .A2(new_n438), .A3(new_n442), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT29), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT86), .B1(new_n492), .B2(new_n310), .ZN(new_n493));
  NAND2_X1  g292(.A1(G228gat), .A2(G233gat), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n374), .B1(new_n443), .B2(new_n444), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT86), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(new_n496), .A3(new_n311), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT29), .B1(new_n303), .B2(new_n307), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n436), .B1(new_n498), .B2(KEYINPUT3), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n493), .A2(new_n494), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT31), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n490), .A2(new_n491), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n310), .B1(new_n502), .B2(new_n374), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n310), .A2(new_n374), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n441), .B1(new_n504), .B2(new_n442), .ZN(new_n505));
  OAI211_X1 g304(.A(G228gat), .B(G233gat), .C1(new_n503), .C2(new_n505), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n500), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n501), .B1(new_n500), .B2(new_n506), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n488), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n500), .A2(new_n506), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT31), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n500), .A2(new_n501), .A3(new_n506), .ZN(new_n512));
  INV_X1    g311(.A(new_n488), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G22gat), .B(G50gat), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n509), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n515), .B1(new_n509), .B2(new_n514), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n445), .A2(new_n452), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n455), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n520), .B(KEYINPUT87), .Z(new_n521));
  INV_X1    g320(.A(KEYINPUT39), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n520), .B(KEYINPUT87), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n456), .A2(new_n457), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n522), .B1(new_n525), .B2(new_n453), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n523), .A2(new_n527), .A3(new_n465), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT40), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n523), .A2(new_n527), .A3(KEYINPUT40), .A4(new_n465), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n530), .A2(new_n468), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n392), .A2(new_n394), .A3(new_n390), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT81), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n392), .A2(new_n394), .A3(KEYINPUT81), .A4(new_n390), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT82), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n538), .B(new_n539), .C1(new_n477), .C2(new_n390), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT30), .B1(new_n483), .B2(KEYINPUT82), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n537), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n518), .B1(new_n532), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n487), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n537), .A2(new_n474), .A3(new_n540), .A4(new_n541), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n518), .A2(new_n545), .ZN(new_n546));
  AND4_X1   g345(.A1(KEYINPUT74), .A2(new_n368), .A3(new_n449), .A4(new_n369), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT74), .B1(new_n366), .B2(new_n449), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT34), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n370), .A2(new_n418), .ZN(new_n551));
  NAND2_X1  g350(.A1(G227gat), .A2(G233gat), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n552), .B(KEYINPUT64), .Z(new_n553));
  NAND4_X1  g352(.A1(new_n549), .A2(new_n550), .A3(new_n551), .A4(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n368), .A2(new_n449), .A3(new_n369), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT74), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n366), .A2(KEYINPUT74), .A3(new_n449), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n557), .A2(new_n551), .A3(new_n558), .A4(new_n552), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT34), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n554), .A2(KEYINPUT76), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT76), .B1(new_n554), .B2(new_n560), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n557), .A2(new_n551), .A3(new_n558), .ZN(new_n564));
  INV_X1    g363(.A(new_n553), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT32), .ZN(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT75), .B(KEYINPUT33), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G15gat), .B(G43gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(G71gat), .B(G99gat), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n571), .B(new_n572), .Z(new_n573));
  NAND3_X1  g372(.A1(new_n567), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT32), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n575), .B1(new_n564), .B2(new_n565), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n568), .B1(new_n564), .B2(new_n565), .ZN(new_n577));
  INV_X1    g376(.A(new_n573), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT78), .B1(new_n563), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n563), .A2(new_n580), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT76), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n559), .A2(KEYINPUT34), .ZN(new_n584));
  NOR3_X1   g383(.A1(new_n564), .A2(KEYINPUT34), .A3(new_n565), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n554), .A2(KEYINPUT76), .A3(new_n560), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT78), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n588), .A2(new_n589), .A3(new_n579), .A4(new_n574), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n581), .A2(new_n582), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT36), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR3_X1   g392(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n594));
  AOI221_X4 g393(.A(new_n575), .B1(new_n568), .B2(new_n573), .C1(new_n564), .C2(new_n565), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT77), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n563), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n588), .A2(new_n580), .A3(KEYINPUT77), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT36), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n593), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n544), .A2(new_n546), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n591), .ZN(new_n603));
  NOR3_X1   g402(.A1(new_n518), .A2(new_n545), .A3(KEYINPUT35), .ZN(new_n604));
  AND4_X1   g403(.A1(new_n474), .A2(new_n537), .A3(new_n540), .A4(new_n541), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n509), .A2(new_n514), .ZN(new_n606));
  INV_X1    g405(.A(new_n515), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n509), .A2(new_n514), .A3(new_n515), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n605), .A2(new_n599), .A3(new_n610), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n603), .A2(new_n604), .B1(new_n611), .B2(KEYINPUT35), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n297), .B1(new_n602), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n251), .A2(KEYINPUT99), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n250), .B(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(new_n210), .A3(new_n211), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT10), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n617), .B(new_n618), .C1(new_n214), .C2(new_n255), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n214), .A2(new_n255), .A3(KEYINPUT10), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n617), .B1(new_n214), .B2(new_n255), .ZN(new_n624));
  INV_X1    g423(.A(new_n622), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G120gat), .B(G148gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT100), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G176gat), .ZN(new_n629));
  INV_X1    g428(.A(G204gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n623), .A2(new_n626), .A3(new_n632), .ZN(new_n633));
  AOI211_X1 g432(.A(KEYINPUT101), .B(new_n625), .C1(new_n619), .C2(new_n620), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n635), .B1(new_n621), .B2(new_n622), .ZN(new_n636));
  AOI211_X1 g435(.A(new_n634), .B(new_n636), .C1(new_n625), .C2(new_n624), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n633), .B1(new_n637), .B2(new_n632), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n278), .A2(new_n225), .ZN(new_n640));
  NAND2_X1  g439(.A1(G229gat), .A2(G233gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n225), .A2(new_n271), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT18), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT94), .B1(new_n225), .B2(new_n271), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(new_n642), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n641), .B(KEYINPUT13), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n642), .B1(new_n278), .B2(new_n225), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(KEYINPUT18), .A3(new_n641), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n646), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G169gat), .B(G197gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G113gat), .B(G141gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT92), .B(KEYINPUT11), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT12), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n646), .A2(new_n651), .A3(new_n660), .A4(new_n653), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n639), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n614), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n474), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n542), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT16), .B(G8gat), .Z(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT102), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n675), .A2(KEYINPUT42), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n672), .A2(G8gat), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(KEYINPUT42), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(G1325gat));
  INV_X1    g478(.A(new_n601), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n668), .A2(G15gat), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(G15gat), .B1(new_n668), .B2(new_n603), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(KEYINPUT103), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(KEYINPUT103), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(G1326gat));
  NOR2_X1   g484(.A1(new_n667), .A2(new_n610), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT43), .B(G22gat), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  AOI21_X1  g487(.A(new_n292), .B1(new_n602), .B2(new_n613), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n666), .A2(new_n295), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(G29gat), .A3(new_n474), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT45), .Z(new_n694));
  NAND2_X1  g493(.A1(new_n601), .A2(new_n546), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n695), .B1(new_n543), .B2(new_n487), .ZN(new_n696));
  OAI211_X1 g495(.A(KEYINPUT44), .B(new_n291), .C1(new_n696), .C2(new_n612), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT104), .B1(new_n605), .B2(new_n610), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n518), .A2(new_n700), .A3(new_n545), .ZN(new_n701));
  AOI22_X1  g500(.A1(new_n699), .A2(new_n701), .B1(new_n593), .B2(new_n600), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n612), .B1(new_n544), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n698), .B1(new_n703), .B2(new_n292), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n697), .A2(new_n704), .A3(new_n691), .ZN(new_n705));
  OAI21_X1  g504(.A(G29gat), .B1(new_n705), .B2(new_n474), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n694), .A2(new_n706), .ZN(G1328gat));
  INV_X1    g506(.A(new_n542), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n692), .A2(G36gat), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT46), .ZN(new_n710));
  OAI21_X1  g509(.A(G36gat), .B1(new_n705), .B2(new_n708), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1329gat));
  NOR2_X1   g511(.A1(new_n692), .A2(new_n591), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n680), .A2(G43gat), .ZN(new_n714));
  OAI22_X1  g513(.A1(new_n713), .A2(G43gat), .B1(new_n705), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g515(.A(G50gat), .B1(new_n705), .B2(new_n610), .ZN(new_n717));
  OR3_X1    g516(.A1(new_n692), .A2(G50gat), .A3(new_n610), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT48), .Z(G1331gat));
  INV_X1    g519(.A(new_n664), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n294), .A2(new_n721), .A3(new_n296), .A4(new_n638), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT105), .Z(new_n723));
  OR3_X1    g522(.A1(new_n723), .A2(KEYINPUT106), .A3(new_n703), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT106), .B1(new_n723), .B2(new_n703), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n474), .B(KEYINPUT107), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g529(.A(KEYINPUT49), .B(G64gat), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n727), .A2(new_n542), .A3(new_n731), .ZN(new_n732));
  OAI22_X1  g531(.A1(new_n726), .A2(new_n708), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(G1333gat));
  OAI21_X1  g533(.A(G71gat), .B1(new_n726), .B2(new_n601), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n591), .B(KEYINPUT108), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n204), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n726), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n735), .B(new_n739), .C1(new_n726), .C2(new_n737), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1334gat));
  NOR2_X1   g542(.A1(new_n726), .A2(new_n610), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT110), .B(G78gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1335gat));
  NOR2_X1   g545(.A1(new_n243), .A2(new_n664), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n639), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n697), .A2(new_n704), .A3(new_n749), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n750), .A2(new_n247), .A3(new_n474), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n544), .A2(new_n702), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n292), .B1(new_n753), .B2(new_n613), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n752), .B1(new_n754), .B2(new_n747), .ZN(new_n755));
  NOR4_X1   g554(.A1(new_n703), .A2(KEYINPUT51), .A3(new_n292), .A4(new_n748), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n755), .A2(new_n756), .A3(new_n639), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n669), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n751), .B1(new_n758), .B2(new_n247), .ZN(G1336gat));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n755), .A2(new_n756), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n761), .A2(new_n248), .A3(new_n638), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n762), .B2(new_n708), .ZN(new_n763));
  OAI21_X1  g562(.A(G92gat), .B1(new_n750), .B2(new_n708), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n762), .B2(new_n708), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n763), .A2(new_n765), .A3(KEYINPUT52), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  OAI221_X1 g566(.A(new_n764), .B1(new_n760), .B2(new_n767), .C1(new_n762), .C2(new_n708), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(G1337gat));
  INV_X1    g568(.A(G99gat), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n757), .A2(new_n770), .A3(new_n603), .ZN(new_n771));
  OAI21_X1  g570(.A(G99gat), .B1(new_n750), .B2(new_n601), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(G1338gat));
  NAND2_X1  g572(.A1(new_n753), .A2(new_n613), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(new_n291), .A3(new_n747), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT51), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n754), .A2(new_n752), .A3(new_n747), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n610), .A2(G106gat), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n776), .A2(new_n638), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n761), .A2(KEYINPUT113), .A3(new_n638), .A4(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n697), .A2(new_n704), .A3(new_n518), .A4(new_n749), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G106gat), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n784), .A2(KEYINPUT112), .A3(G106gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT53), .B1(new_n783), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n779), .A2(new_n785), .A3(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n779), .A2(new_n785), .A3(KEYINPUT114), .A4(new_n791), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n790), .A2(new_n796), .ZN(G1339gat));
  OR3_X1    g596(.A1(new_n652), .A2(KEYINPUT116), .A3(new_n641), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT116), .B1(new_n652), .B2(new_n641), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n798), .B(new_n799), .C1(new_n650), .C2(new_n648), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n659), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n638), .A2(new_n801), .A3(new_n663), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n621), .A2(new_n622), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT115), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n623), .A2(KEYINPUT115), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n804), .B(KEYINPUT54), .C1(new_n805), .C2(new_n803), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n636), .B2(new_n634), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n806), .A2(KEYINPUT55), .A3(new_n631), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n664), .A2(new_n633), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n806), .A2(new_n631), .A3(new_n808), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n802), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n292), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n291), .A2(new_n663), .A3(new_n801), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n811), .A2(new_n812), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n817), .A2(new_n633), .A3(new_n809), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n243), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n294), .A2(new_n721), .A3(new_n296), .A4(new_n639), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(new_n610), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n542), .A2(new_n474), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n603), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(G113gat), .B1(new_n826), .B2(new_n721), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n823), .A2(new_n708), .A3(new_n728), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n599), .A2(new_n610), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n664), .A2(new_n406), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n827), .B1(new_n831), .B2(new_n832), .ZN(G1340gat));
  OAI21_X1  g632(.A(G120gat), .B1(new_n826), .B2(new_n639), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n408), .A2(new_n410), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n638), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n834), .B1(new_n831), .B2(new_n836), .ZN(G1341gat));
  NOR3_X1   g636(.A1(new_n826), .A2(new_n217), .A3(new_n295), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n838), .A2(KEYINPUT117), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n217), .B1(new_n831), .B2(new_n295), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(KEYINPUT117), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(G1342gat));
  NOR3_X1   g641(.A1(new_n831), .A2(G134gat), .A3(new_n292), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT56), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  OAI21_X1  g645(.A(G134gat), .B1(new_n826), .B2(new_n292), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(G1343gat));
  NAND2_X1  g647(.A1(new_n601), .A2(new_n825), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n823), .A2(new_n518), .ZN(new_n850));
  XNOR2_X1  g649(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n817), .A2(KEYINPUT119), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n809), .A2(new_n633), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n811), .A2(new_n856), .A3(new_n812), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n854), .A2(new_n855), .A3(new_n664), .A4(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n291), .B1(new_n858), .B2(new_n802), .ZN(new_n859));
  INV_X1    g658(.A(new_n819), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n295), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n610), .B1(new_n861), .B2(new_n821), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(KEYINPUT57), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n849), .B1(new_n853), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n422), .B1(new_n864), .B2(new_n664), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n680), .A2(new_n610), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n828), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n721), .A2(G141gat), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(KEYINPUT120), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n868), .A2(KEYINPUT120), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT58), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n853), .A2(new_n863), .ZN(new_n873));
  INV_X1    g672(.A(new_n849), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n664), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(KEYINPUT121), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n877), .B1(new_n864), .B2(new_n664), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n876), .A2(new_n422), .A3(new_n878), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n871), .A2(KEYINPUT58), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n872), .B1(new_n879), .B2(new_n880), .ZN(G1344gat));
  INV_X1    g680(.A(new_n867), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n423), .A3(new_n638), .ZN(new_n883));
  AOI211_X1 g682(.A(new_n639), .B(new_n849), .C1(new_n853), .C2(new_n863), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n423), .A2(KEYINPUT59), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT122), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n864), .A2(new_n638), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n889), .A3(new_n885), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n518), .B(new_n851), .C1(new_n820), .C2(new_n822), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n893), .B1(new_n862), .B2(KEYINPUT57), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n638), .A3(new_n874), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n892), .B1(new_n895), .B2(G148gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n883), .B1(new_n891), .B2(new_n896), .ZN(G1345gat));
  AOI21_X1  g696(.A(G155gat), .B1(new_n882), .B2(new_n243), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n295), .A2(new_n419), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n864), .B2(new_n899), .ZN(G1346gat));
  AOI21_X1  g699(.A(G162gat), .B1(new_n882), .B2(new_n291), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n292), .A2(new_n420), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n864), .B2(new_n902), .ZN(G1347gat));
  NOR2_X1   g702(.A1(new_n728), .A2(new_n708), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n824), .A2(new_n736), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(G169gat), .B1(new_n905), .B2(new_n721), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n823), .A2(new_n474), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n542), .A3(new_n830), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n664), .A2(new_n339), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(G1348gat));
  NOR3_X1   g709(.A1(new_n905), .A2(new_n639), .A3(new_n360), .ZN(new_n911));
  INV_X1    g710(.A(new_n908), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n638), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n911), .B1(new_n340), .B2(new_n913), .ZN(G1349gat));
  OAI211_X1 g713(.A(new_n912), .B(new_n243), .C1(new_n332), .C2(new_n331), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n326), .B1(new_n905), .B2(new_n295), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT60), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n915), .A2(new_n919), .A3(new_n916), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1350gat));
  NAND3_X1  g720(.A1(new_n912), .A2(new_n329), .A3(new_n291), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n905), .A2(new_n292), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n923), .A2(new_n924), .A3(G190gat), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n923), .B2(G190gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n922), .B1(new_n925), .B2(new_n926), .ZN(G1351gat));
  NAND2_X1  g726(.A1(new_n601), .A2(new_n904), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n601), .A2(KEYINPUT123), .A3(new_n904), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n931), .B1(new_n930), .B2(new_n932), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n894), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(G197gat), .B1(new_n935), .B2(new_n721), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n907), .A2(new_n542), .A3(new_n866), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n721), .A2(G197gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(G1352gat));
  NOR3_X1   g738(.A1(new_n937), .A2(G204gat), .A3(new_n639), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT62), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n935), .A2(new_n639), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n941), .B1(new_n630), .B2(new_n943), .ZN(G1353gat));
  OR3_X1    g743(.A1(new_n937), .A2(G211gat), .A3(new_n295), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n295), .B1(new_n930), .B2(new_n932), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n894), .A2(new_n946), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n947), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n948));
  AOI21_X1  g747(.A(KEYINPUT63), .B1(new_n947), .B2(G211gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G1354gat));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT125), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n291), .A2(KEYINPUT126), .A3(G218gat), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n894), .B(new_n953), .C1(new_n933), .C2(new_n934), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n955), .B1(new_n292), .B2(new_n301), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n951), .A2(new_n952), .A3(new_n954), .A4(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n301), .B1(new_n937), .B2(new_n292), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n957), .A2(KEYINPUT127), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1355gat));
endmodule


