

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U554 ( .A(KEYINPUT31), .ZN(n726) );
  NOR2_X1 U555 ( .A1(G164), .A2(G1384), .ZN(n775) );
  NOR2_X1 U556 ( .A1(G651), .A2(n619), .ZN(n644) );
  AND2_X1 U557 ( .A1(G2105), .A2(G2104), .ZN(n869) );
  NAND2_X1 U558 ( .A1(G114), .A2(n869), .ZN(n520) );
  INV_X1 U559 ( .A(G2105), .ZN(n522) );
  NOR2_X1 U560 ( .A1(G2104), .A2(n522), .ZN(n870) );
  NAND2_X1 U561 ( .A1(G126), .A2(n870), .ZN(n519) );
  NAND2_X1 U562 ( .A1(n520), .A2(n519), .ZN(n528) );
  NOR2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n521), .Z(n867) );
  NAND2_X1 U565 ( .A1(G138), .A2(n867), .ZN(n524) );
  AND2_X1 U566 ( .A1(n522), .A2(G2104), .ZN(n875) );
  NAND2_X1 U567 ( .A1(G102), .A2(n875), .ZN(n523) );
  NAND2_X1 U568 ( .A1(n524), .A2(n523), .ZN(n526) );
  INV_X1 U569 ( .A(KEYINPUT91), .ZN(n525) );
  XNOR2_X1 U570 ( .A(n526), .B(n525), .ZN(n527) );
  NOR2_X1 U571 ( .A1(n528), .A2(n527), .ZN(G164) );
  INV_X1 U572 ( .A(G651), .ZN(n534) );
  NOR2_X1 U573 ( .A1(G543), .A2(n534), .ZN(n529) );
  XOR2_X1 U574 ( .A(KEYINPUT1), .B(n529), .Z(n643) );
  NAND2_X1 U575 ( .A1(G64), .A2(n643), .ZN(n531) );
  XOR2_X1 U576 ( .A(G543), .B(KEYINPUT0), .Z(n619) );
  NAND2_X1 U577 ( .A1(G52), .A2(n644), .ZN(n530) );
  NAND2_X1 U578 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U579 ( .A(KEYINPUT66), .B(n532), .ZN(n539) );
  NOR2_X1 U580 ( .A1(G651), .A2(G543), .ZN(n639) );
  NAND2_X1 U581 ( .A1(n639), .A2(G90), .ZN(n533) );
  XOR2_X1 U582 ( .A(KEYINPUT67), .B(n533), .Z(n536) );
  NOR2_X1 U583 ( .A1(n619), .A2(n534), .ZN(n638) );
  NAND2_X1 U584 ( .A1(n638), .A2(G77), .ZN(n535) );
  NAND2_X1 U585 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U586 ( .A(KEYINPUT9), .B(n537), .Z(n538) );
  NOR2_X1 U587 ( .A1(n539), .A2(n538), .ZN(G171) );
  AND2_X1 U588 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U589 ( .A(G57), .ZN(G237) );
  INV_X1 U590 ( .A(G132), .ZN(G219) );
  INV_X1 U591 ( .A(G82), .ZN(G220) );
  NAND2_X1 U592 ( .A1(n639), .A2(G89), .ZN(n540) );
  XNOR2_X1 U593 ( .A(n540), .B(KEYINPUT4), .ZN(n542) );
  NAND2_X1 U594 ( .A1(G76), .A2(n638), .ZN(n541) );
  NAND2_X1 U595 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U596 ( .A(n543), .B(KEYINPUT5), .ZN(n549) );
  XNOR2_X1 U597 ( .A(KEYINPUT77), .B(KEYINPUT6), .ZN(n547) );
  NAND2_X1 U598 ( .A1(G63), .A2(n643), .ZN(n545) );
  NAND2_X1 U599 ( .A1(G51), .A2(n644), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U601 ( .A(n547), .B(n546), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U603 ( .A(KEYINPUT7), .B(n550), .ZN(G168) );
  XOR2_X1 U604 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U605 ( .A(KEYINPUT70), .B(KEYINPUT10), .Z(n552) );
  NAND2_X1 U606 ( .A1(G7), .A2(G661), .ZN(n551) );
  XNOR2_X1 U607 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U608 ( .A(KEYINPUT69), .B(n553), .ZN(G223) );
  INV_X1 U609 ( .A(G223), .ZN(n825) );
  NAND2_X1 U610 ( .A1(n825), .A2(G567), .ZN(n554) );
  XOR2_X1 U611 ( .A(KEYINPUT11), .B(n554), .Z(G234) );
  NAND2_X1 U612 ( .A1(n643), .A2(G56), .ZN(n555) );
  XNOR2_X1 U613 ( .A(n555), .B(KEYINPUT14), .ZN(n563) );
  NAND2_X1 U614 ( .A1(n638), .A2(G68), .ZN(n556) );
  XNOR2_X1 U615 ( .A(KEYINPUT71), .B(n556), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n639), .A2(G81), .ZN(n557) );
  XOR2_X1 U617 ( .A(n557), .B(KEYINPUT12), .Z(n558) );
  NOR2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U619 ( .A(KEYINPUT72), .B(n560), .Z(n561) );
  XNOR2_X1 U620 ( .A(KEYINPUT13), .B(n561), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U622 ( .A(n564), .B(KEYINPUT73), .ZN(n566) );
  NAND2_X1 U623 ( .A1(G43), .A2(n644), .ZN(n565) );
  NAND2_X1 U624 ( .A1(n566), .A2(n565), .ZN(n955) );
  INV_X1 U625 ( .A(G860), .ZN(n590) );
  OR2_X1 U626 ( .A1(n955), .A2(n590), .ZN(G153) );
  INV_X1 U627 ( .A(G171), .ZN(G301) );
  INV_X1 U628 ( .A(G868), .ZN(n661) );
  NOR2_X1 U629 ( .A1(G301), .A2(n661), .ZN(n577) );
  NAND2_X1 U630 ( .A1(G92), .A2(n639), .ZN(n568) );
  NAND2_X1 U631 ( .A1(G66), .A2(n643), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT74), .B(n569), .ZN(n573) );
  NAND2_X1 U634 ( .A1(G79), .A2(n638), .ZN(n571) );
  NAND2_X1 U635 ( .A1(G54), .A2(n644), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT15), .B(n574), .Z(n575) );
  XNOR2_X1 U639 ( .A(KEYINPUT75), .B(n575), .ZN(n940) );
  NOR2_X1 U640 ( .A1(G868), .A2(n940), .ZN(n576) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT76), .B(n578), .ZN(G284) );
  NAND2_X1 U643 ( .A1(G78), .A2(n638), .ZN(n580) );
  NAND2_X1 U644 ( .A1(G91), .A2(n639), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U646 ( .A1(n643), .A2(G65), .ZN(n581) );
  XOR2_X1 U647 ( .A(KEYINPUT68), .B(n581), .Z(n582) );
  NOR2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U649 ( .A1(n644), .A2(G53), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(G299) );
  NOR2_X1 U651 ( .A1(G868), .A2(G299), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n586), .B(KEYINPUT78), .ZN(n588) );
  NOR2_X1 U653 ( .A1(n661), .A2(G286), .ZN(n587) );
  NOR2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U655 ( .A(KEYINPUT79), .B(n589), .Z(G297) );
  NAND2_X1 U656 ( .A1(n590), .A2(G559), .ZN(n591) );
  INV_X1 U657 ( .A(n940), .ZN(n897) );
  NAND2_X1 U658 ( .A1(n591), .A2(n897), .ZN(n592) );
  XNOR2_X1 U659 ( .A(n592), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U660 ( .A1(G868), .A2(n955), .ZN(n595) );
  NAND2_X1 U661 ( .A1(G868), .A2(n897), .ZN(n593) );
  NOR2_X1 U662 ( .A1(G559), .A2(n593), .ZN(n594) );
  NOR2_X1 U663 ( .A1(n595), .A2(n594), .ZN(G282) );
  NAND2_X1 U664 ( .A1(G99), .A2(n875), .ZN(n597) );
  NAND2_X1 U665 ( .A1(G111), .A2(n869), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U667 ( .A(KEYINPUT80), .B(n598), .ZN(n603) );
  NAND2_X1 U668 ( .A1(G123), .A2(n870), .ZN(n599) );
  XNOR2_X1 U669 ( .A(n599), .B(KEYINPUT18), .ZN(n601) );
  NAND2_X1 U670 ( .A1(n867), .A2(G135), .ZN(n600) );
  NAND2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U672 ( .A1(n603), .A2(n602), .ZN(n1010) );
  XNOR2_X1 U673 ( .A(n1010), .B(G2096), .ZN(n605) );
  INV_X1 U674 ( .A(G2100), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n605), .A2(n604), .ZN(G156) );
  NAND2_X1 U676 ( .A1(G80), .A2(n638), .ZN(n607) );
  NAND2_X1 U677 ( .A1(G93), .A2(n639), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U679 ( .A1(G67), .A2(n643), .ZN(n608) );
  XNOR2_X1 U680 ( .A(KEYINPUT81), .B(n608), .ZN(n609) );
  NOR2_X1 U681 ( .A1(n610), .A2(n609), .ZN(n612) );
  NAND2_X1 U682 ( .A1(n644), .A2(G55), .ZN(n611) );
  NAND2_X1 U683 ( .A1(n612), .A2(n611), .ZN(n660) );
  NAND2_X1 U684 ( .A1(n897), .A2(G559), .ZN(n658) );
  XNOR2_X1 U685 ( .A(n955), .B(n658), .ZN(n613) );
  NOR2_X1 U686 ( .A1(G860), .A2(n613), .ZN(n614) );
  XOR2_X1 U687 ( .A(n660), .B(n614), .Z(G145) );
  NAND2_X1 U688 ( .A1(G49), .A2(n644), .ZN(n616) );
  NAND2_X1 U689 ( .A1(G74), .A2(G651), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U691 ( .A(KEYINPUT82), .B(n617), .ZN(n618) );
  NOR2_X1 U692 ( .A1(n643), .A2(n618), .ZN(n621) );
  NAND2_X1 U693 ( .A1(n619), .A2(G87), .ZN(n620) );
  NAND2_X1 U694 ( .A1(n621), .A2(n620), .ZN(G288) );
  NAND2_X1 U695 ( .A1(G86), .A2(n639), .ZN(n623) );
  NAND2_X1 U696 ( .A1(G61), .A2(n643), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U698 ( .A1(n638), .A2(G73), .ZN(n624) );
  XOR2_X1 U699 ( .A(KEYINPUT2), .B(n624), .Z(n625) );
  NOR2_X1 U700 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U701 ( .A(KEYINPUT83), .B(n627), .Z(n629) );
  NAND2_X1 U702 ( .A1(n644), .A2(G48), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(G305) );
  NAND2_X1 U704 ( .A1(G62), .A2(n643), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G50), .A2(n644), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U707 ( .A(KEYINPUT84), .B(n632), .Z(n634) );
  NAND2_X1 U708 ( .A1(n639), .A2(G88), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U710 ( .A1(G75), .A2(n638), .ZN(n635) );
  XNOR2_X1 U711 ( .A(KEYINPUT85), .B(n635), .ZN(n636) );
  NOR2_X1 U712 ( .A1(n637), .A2(n636), .ZN(G166) );
  NAND2_X1 U713 ( .A1(G72), .A2(n638), .ZN(n641) );
  NAND2_X1 U714 ( .A1(G85), .A2(n639), .ZN(n640) );
  NAND2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U716 ( .A(KEYINPUT65), .B(n642), .ZN(n648) );
  NAND2_X1 U717 ( .A1(G60), .A2(n643), .ZN(n646) );
  NAND2_X1 U718 ( .A1(G47), .A2(n644), .ZN(n645) );
  AND2_X1 U719 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U720 ( .A1(n648), .A2(n647), .ZN(G290) );
  INV_X1 U721 ( .A(G299), .ZN(n696) );
  XOR2_X1 U722 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n650) );
  XNOR2_X1 U723 ( .A(KEYINPUT88), .B(KEYINPUT19), .ZN(n649) );
  XNOR2_X1 U724 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U725 ( .A(n651), .B(G288), .ZN(n652) );
  XNOR2_X1 U726 ( .A(n652), .B(n660), .ZN(n653) );
  XNOR2_X1 U727 ( .A(n696), .B(n653), .ZN(n656) );
  XOR2_X1 U728 ( .A(G166), .B(G290), .Z(n654) );
  XNOR2_X1 U729 ( .A(G305), .B(n654), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n955), .B(n657), .ZN(n895) );
  XNOR2_X1 U732 ( .A(n658), .B(n895), .ZN(n659) );
  NAND2_X1 U733 ( .A1(n659), .A2(G868), .ZN(n663) );
  NAND2_X1 U734 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U735 ( .A1(n663), .A2(n662), .ZN(G295) );
  NAND2_X1 U736 ( .A1(G2078), .A2(G2084), .ZN(n664) );
  XOR2_X1 U737 ( .A(KEYINPUT20), .B(n664), .Z(n665) );
  NAND2_X1 U738 ( .A1(G2090), .A2(n665), .ZN(n666) );
  XNOR2_X1 U739 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U740 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U741 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U742 ( .A1(G661), .A2(G483), .ZN(n676) );
  NOR2_X1 U743 ( .A1(G220), .A2(G219), .ZN(n668) );
  XOR2_X1 U744 ( .A(KEYINPUT22), .B(n668), .Z(n669) );
  NOR2_X1 U745 ( .A1(G218), .A2(n669), .ZN(n670) );
  XOR2_X1 U746 ( .A(KEYINPUT89), .B(n670), .Z(n671) );
  NAND2_X1 U747 ( .A1(G96), .A2(n671), .ZN(n829) );
  NAND2_X1 U748 ( .A1(n829), .A2(G2106), .ZN(n675) );
  NAND2_X1 U749 ( .A1(G69), .A2(G120), .ZN(n672) );
  NOR2_X1 U750 ( .A1(G237), .A2(n672), .ZN(n673) );
  NAND2_X1 U751 ( .A1(G108), .A2(n673), .ZN(n830) );
  NAND2_X1 U752 ( .A1(n830), .A2(G567), .ZN(n674) );
  NAND2_X1 U753 ( .A1(n675), .A2(n674), .ZN(n850) );
  NOR2_X1 U754 ( .A1(n676), .A2(n850), .ZN(n677) );
  XNOR2_X1 U755 ( .A(n677), .B(KEYINPUT90), .ZN(n828) );
  NAND2_X1 U756 ( .A1(G36), .A2(n828), .ZN(G176) );
  NAND2_X1 U757 ( .A1(n869), .A2(G113), .ZN(n680) );
  NAND2_X1 U758 ( .A1(G101), .A2(n875), .ZN(n678) );
  XOR2_X1 U759 ( .A(KEYINPUT23), .B(n678), .Z(n679) );
  NAND2_X1 U760 ( .A1(n680), .A2(n679), .ZN(n684) );
  NAND2_X1 U761 ( .A1(G137), .A2(n867), .ZN(n682) );
  NAND2_X1 U762 ( .A1(G125), .A2(n870), .ZN(n681) );
  NAND2_X1 U763 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U764 ( .A1(n684), .A2(n683), .ZN(G160) );
  XOR2_X1 U765 ( .A(KEYINPUT92), .B(G166), .Z(G303) );
  NOR2_X1 U766 ( .A1(G1981), .A2(G305), .ZN(n685) );
  XNOR2_X1 U767 ( .A(KEYINPUT24), .B(n685), .ZN(n688) );
  NAND2_X1 U768 ( .A1(G160), .A2(G40), .ZN(n774) );
  INV_X1 U769 ( .A(n774), .ZN(n686) );
  NAND2_X1 U770 ( .A1(n686), .A2(n775), .ZN(n687) );
  XNOR2_X2 U771 ( .A(n687), .B(KEYINPUT64), .ZN(n732) );
  NAND2_X1 U772 ( .A1(n732), .A2(G8), .ZN(n757) );
  INV_X1 U773 ( .A(n757), .ZN(n758) );
  NAND2_X1 U774 ( .A1(n688), .A2(n758), .ZN(n752) );
  NOR2_X1 U775 ( .A1(n732), .A2(G2084), .ZN(n718) );
  NAND2_X1 U776 ( .A1(G8), .A2(n718), .ZN(n731) );
  NOR2_X1 U777 ( .A1(G1966), .A2(n757), .ZN(n729) );
  INV_X1 U778 ( .A(n732), .ZN(n702) );
  XNOR2_X1 U779 ( .A(G2078), .B(KEYINPUT25), .ZN(n924) );
  NAND2_X1 U780 ( .A1(n702), .A2(n924), .ZN(n690) );
  XNOR2_X1 U781 ( .A(KEYINPUT97), .B(G1961), .ZN(n966) );
  NAND2_X1 U782 ( .A1(n732), .A2(n966), .ZN(n689) );
  NAND2_X1 U783 ( .A1(n690), .A2(n689), .ZN(n723) );
  NAND2_X1 U784 ( .A1(n723), .A2(G171), .ZN(n717) );
  XNOR2_X1 U785 ( .A(KEYINPUT29), .B(KEYINPUT99), .ZN(n715) );
  NAND2_X1 U786 ( .A1(G2072), .A2(n702), .ZN(n691) );
  XNOR2_X1 U787 ( .A(n691), .B(KEYINPUT27), .ZN(n693) );
  INV_X1 U788 ( .A(G1956), .ZN(n969) );
  NOR2_X1 U789 ( .A1(n702), .A2(n969), .ZN(n692) );
  NOR2_X1 U790 ( .A1(n693), .A2(n692), .ZN(n697) );
  NOR2_X1 U791 ( .A1(n697), .A2(n696), .ZN(n695) );
  XOR2_X1 U792 ( .A(KEYINPUT98), .B(KEYINPUT28), .Z(n694) );
  XNOR2_X1 U793 ( .A(n695), .B(n694), .ZN(n713) );
  NAND2_X1 U794 ( .A1(n697), .A2(n696), .ZN(n711) );
  NAND2_X1 U795 ( .A1(n702), .A2(G1996), .ZN(n698) );
  XNOR2_X1 U796 ( .A(n698), .B(KEYINPUT26), .ZN(n700) );
  NAND2_X1 U797 ( .A1(n732), .A2(G1341), .ZN(n699) );
  NAND2_X1 U798 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U799 ( .A1(n955), .A2(n701), .ZN(n706) );
  NAND2_X1 U800 ( .A1(G2067), .A2(n702), .ZN(n704) );
  NAND2_X1 U801 ( .A1(n732), .A2(G1348), .ZN(n703) );
  NAND2_X1 U802 ( .A1(n704), .A2(n703), .ZN(n707) );
  NOR2_X1 U803 ( .A1(n940), .A2(n707), .ZN(n705) );
  OR2_X1 U804 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U805 ( .A1(n940), .A2(n707), .ZN(n708) );
  NAND2_X1 U806 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U807 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U809 ( .A(n715), .B(n714), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n717), .A2(n716), .ZN(n738) );
  NOR2_X1 U811 ( .A1(n729), .A2(n718), .ZN(n719) );
  XNOR2_X1 U812 ( .A(KEYINPUT100), .B(n719), .ZN(n720) );
  NAND2_X1 U813 ( .A1(n720), .A2(G8), .ZN(n721) );
  XNOR2_X1 U814 ( .A(n721), .B(KEYINPUT30), .ZN(n722) );
  NOR2_X1 U815 ( .A1(G168), .A2(n722), .ZN(n725) );
  NOR2_X1 U816 ( .A1(G171), .A2(n723), .ZN(n724) );
  NOR2_X1 U817 ( .A1(n725), .A2(n724), .ZN(n727) );
  XNOR2_X1 U818 ( .A(n727), .B(n726), .ZN(n740) );
  AND2_X1 U819 ( .A1(n738), .A2(n740), .ZN(n728) );
  NOR2_X1 U820 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U821 ( .A1(n731), .A2(n730), .ZN(n747) );
  INV_X1 U822 ( .A(G8), .ZN(n737) );
  NOR2_X1 U823 ( .A1(n732), .A2(G2090), .ZN(n734) );
  NOR2_X1 U824 ( .A1(G1971), .A2(n757), .ZN(n733) );
  NOR2_X1 U825 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U826 ( .A1(n735), .A2(G303), .ZN(n736) );
  OR2_X1 U827 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U828 ( .A1(n738), .A2(n741), .ZN(n739) );
  NAND2_X1 U829 ( .A1(n740), .A2(n739), .ZN(n744) );
  INV_X1 U830 ( .A(n741), .ZN(n742) );
  OR2_X1 U831 ( .A1(n742), .A2(G286), .ZN(n743) );
  NAND2_X1 U832 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U833 ( .A(n745), .B(KEYINPUT32), .ZN(n746) );
  NAND2_X1 U834 ( .A1(n747), .A2(n746), .ZN(n755) );
  NOR2_X1 U835 ( .A1(G2090), .A2(G303), .ZN(n748) );
  NAND2_X1 U836 ( .A1(G8), .A2(n748), .ZN(n749) );
  NAND2_X1 U837 ( .A1(n755), .A2(n749), .ZN(n750) );
  NAND2_X1 U838 ( .A1(n757), .A2(n750), .ZN(n751) );
  NAND2_X1 U839 ( .A1(n752), .A2(n751), .ZN(n772) );
  NOR2_X1 U840 ( .A1(G303), .A2(G1971), .ZN(n753) );
  NOR2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n943) );
  NOR2_X1 U842 ( .A1(n753), .A2(n943), .ZN(n754) );
  AND2_X1 U843 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U844 ( .A1(n757), .A2(n756), .ZN(n764) );
  NAND2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n949) );
  INV_X1 U846 ( .A(KEYINPUT33), .ZN(n766) );
  NAND2_X1 U847 ( .A1(n758), .A2(n943), .ZN(n759) );
  NOR2_X1 U848 ( .A1(n766), .A2(n759), .ZN(n760) );
  XNOR2_X1 U849 ( .A(n760), .B(KEYINPUT101), .ZN(n765) );
  AND2_X1 U850 ( .A1(n949), .A2(n765), .ZN(n762) );
  XNOR2_X1 U851 ( .A(G1981), .B(G305), .ZN(n961) );
  INV_X1 U852 ( .A(n961), .ZN(n761) );
  AND2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n770) );
  INV_X1 U855 ( .A(n765), .ZN(n767) );
  OR2_X1 U856 ( .A1(n767), .A2(n766), .ZN(n768) );
  OR2_X1 U857 ( .A1(n961), .A2(n768), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U859 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U860 ( .A(n773), .B(KEYINPUT102), .ZN(n809) );
  NOR2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n820) );
  XNOR2_X1 U862 ( .A(G2067), .B(KEYINPUT37), .ZN(n810) );
  XNOR2_X1 U863 ( .A(KEYINPUT94), .B(KEYINPUT34), .ZN(n779) );
  NAND2_X1 U864 ( .A1(G104), .A2(n875), .ZN(n777) );
  NAND2_X1 U865 ( .A1(G140), .A2(n867), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U867 ( .A(n779), .B(n778), .ZN(n785) );
  NAND2_X1 U868 ( .A1(n869), .A2(G116), .ZN(n780) );
  XOR2_X1 U869 ( .A(KEYINPUT95), .B(n780), .Z(n782) );
  NAND2_X1 U870 ( .A1(n870), .A2(G128), .ZN(n781) );
  NAND2_X1 U871 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U872 ( .A(KEYINPUT35), .B(n783), .Z(n784) );
  NOR2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U874 ( .A(KEYINPUT36), .B(n786), .ZN(n892) );
  NOR2_X1 U875 ( .A1(n810), .A2(n892), .ZN(n1017) );
  NAND2_X1 U876 ( .A1(n820), .A2(n1017), .ZN(n816) );
  NAND2_X1 U877 ( .A1(G95), .A2(n875), .ZN(n788) );
  NAND2_X1 U878 ( .A1(G131), .A2(n867), .ZN(n787) );
  NAND2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n792) );
  NAND2_X1 U880 ( .A1(G107), .A2(n869), .ZN(n790) );
  NAND2_X1 U881 ( .A1(G119), .A2(n870), .ZN(n789) );
  NAND2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n791) );
  OR2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n880) );
  AND2_X1 U884 ( .A1(n880), .A2(G1991), .ZN(n802) );
  XOR2_X1 U885 ( .A(KEYINPUT96), .B(KEYINPUT38), .Z(n794) );
  NAND2_X1 U886 ( .A1(G105), .A2(n875), .ZN(n793) );
  XNOR2_X1 U887 ( .A(n794), .B(n793), .ZN(n798) );
  NAND2_X1 U888 ( .A1(G117), .A2(n869), .ZN(n796) );
  NAND2_X1 U889 ( .A1(G129), .A2(n870), .ZN(n795) );
  NAND2_X1 U890 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n800) );
  NAND2_X1 U892 ( .A1(n867), .A2(G141), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n885) );
  AND2_X1 U894 ( .A1(n885), .A2(G1996), .ZN(n801) );
  NOR2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n1007) );
  INV_X1 U896 ( .A(n820), .ZN(n803) );
  NOR2_X1 U897 ( .A1(n1007), .A2(n803), .ZN(n813) );
  INV_X1 U898 ( .A(n813), .ZN(n804) );
  AND2_X1 U899 ( .A1(n816), .A2(n804), .ZN(n807) );
  XOR2_X1 U900 ( .A(G1986), .B(KEYINPUT93), .Z(n805) );
  XNOR2_X1 U901 ( .A(G290), .B(n805), .ZN(n942) );
  NAND2_X1 U902 ( .A1(n942), .A2(n820), .ZN(n806) );
  NAND2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n808) );
  OR2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n823) );
  NAND2_X1 U905 ( .A1(n810), .A2(n892), .ZN(n1026) );
  NOR2_X1 U906 ( .A1(G1996), .A2(n885), .ZN(n1005) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n811) );
  NOR2_X1 U908 ( .A1(G1991), .A2(n880), .ZN(n1009) );
  NOR2_X1 U909 ( .A1(n811), .A2(n1009), .ZN(n812) );
  NOR2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U911 ( .A1(n1005), .A2(n814), .ZN(n815) );
  XNOR2_X1 U912 ( .A(n815), .B(KEYINPUT39), .ZN(n817) );
  NAND2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n1026), .A2(n818), .ZN(n819) );
  XOR2_X1 U915 ( .A(KEYINPUT103), .B(n819), .Z(n821) );
  NAND2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U918 ( .A(n824), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n825), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n826) );
  NAND2_X1 U921 ( .A1(G661), .A2(n826), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U923 ( .A1(n828), .A2(n827), .ZN(G188) );
  XOR2_X1 U924 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  INV_X1 U926 ( .A(G120), .ZN(G236) );
  INV_X1 U927 ( .A(G69), .ZN(G235) );
  NOR2_X1 U928 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U929 ( .A(G325), .ZN(G261) );
  XOR2_X1 U930 ( .A(G2100), .B(G2096), .Z(n832) );
  XNOR2_X1 U931 ( .A(KEYINPUT42), .B(G2678), .ZN(n831) );
  XNOR2_X1 U932 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U933 ( .A(KEYINPUT43), .B(G2090), .Z(n834) );
  XNOR2_X1 U934 ( .A(G2067), .B(G2072), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U936 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U937 ( .A(G2078), .B(G2084), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(G227) );
  XOR2_X1 U939 ( .A(KEYINPUT108), .B(G1956), .Z(n840) );
  XNOR2_X1 U940 ( .A(G1996), .B(G1991), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U942 ( .A(n841), .B(KEYINPUT41), .Z(n843) );
  XNOR2_X1 U943 ( .A(G1966), .B(G1961), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U945 ( .A(G1976), .B(G1981), .Z(n845) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1971), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U948 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U949 ( .A(KEYINPUT107), .B(G2474), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(G229) );
  INV_X1 U951 ( .A(n850), .ZN(G319) );
  NAND2_X1 U952 ( .A1(G124), .A2(n870), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n851), .B(KEYINPUT44), .ZN(n854) );
  NAND2_X1 U954 ( .A1(G136), .A2(n867), .ZN(n852) );
  XOR2_X1 U955 ( .A(KEYINPUT109), .B(n852), .Z(n853) );
  NAND2_X1 U956 ( .A1(n854), .A2(n853), .ZN(n858) );
  NAND2_X1 U957 ( .A1(G100), .A2(n875), .ZN(n856) );
  NAND2_X1 U958 ( .A1(G112), .A2(n869), .ZN(n855) );
  NAND2_X1 U959 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U960 ( .A1(n858), .A2(n857), .ZN(G162) );
  NAND2_X1 U961 ( .A1(G118), .A2(n869), .ZN(n860) );
  NAND2_X1 U962 ( .A1(G130), .A2(n870), .ZN(n859) );
  NAND2_X1 U963 ( .A1(n860), .A2(n859), .ZN(n866) );
  NAND2_X1 U964 ( .A1(G106), .A2(n875), .ZN(n862) );
  NAND2_X1 U965 ( .A1(G142), .A2(n867), .ZN(n861) );
  NAND2_X1 U966 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U967 ( .A(KEYINPUT110), .B(n863), .Z(n864) );
  XNOR2_X1 U968 ( .A(KEYINPUT45), .B(n864), .ZN(n865) );
  NOR2_X1 U969 ( .A1(n866), .A2(n865), .ZN(n884) );
  XOR2_X1 U970 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n882) );
  NAND2_X1 U971 ( .A1(n867), .A2(G139), .ZN(n868) );
  XNOR2_X1 U972 ( .A(KEYINPUT111), .B(n868), .ZN(n879) );
  NAND2_X1 U973 ( .A1(G115), .A2(n869), .ZN(n872) );
  NAND2_X1 U974 ( .A1(G127), .A2(n870), .ZN(n871) );
  NAND2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n873), .B(KEYINPUT47), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n874), .B(KEYINPUT112), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n875), .A2(G103), .ZN(n876) );
  NAND2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n1019) );
  XOR2_X1 U981 ( .A(n880), .B(n1019), .Z(n881) );
  XNOR2_X1 U982 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U983 ( .A(n884), .B(n883), .Z(n887) );
  XOR2_X1 U984 ( .A(G160), .B(n885), .Z(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U986 ( .A(n888), .B(G162), .Z(n890) );
  XNOR2_X1 U987 ( .A(G164), .B(n1010), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U989 ( .A(n892), .B(n891), .Z(n893) );
  NOR2_X1 U990 ( .A1(G37), .A2(n893), .ZN(n894) );
  XOR2_X1 U991 ( .A(KEYINPUT113), .B(n894), .Z(G395) );
  XNOR2_X1 U992 ( .A(G286), .B(G301), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U995 ( .A1(G37), .A2(n899), .ZN(G397) );
  XNOR2_X1 U996 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n901) );
  NOR2_X1 U997 ( .A1(G227), .A2(G229), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n914) );
  XNOR2_X1 U999 ( .A(G2446), .B(KEYINPUT104), .ZN(n911) );
  XOR2_X1 U1000 ( .A(G2430), .B(G2427), .Z(n903) );
  XNOR2_X1 U1001 ( .A(KEYINPUT105), .B(G2438), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n907) );
  XOR2_X1 U1003 ( .A(G2435), .B(G2454), .Z(n905) );
  XNOR2_X1 U1004 ( .A(G1341), .B(G1348), .ZN(n904) );
  XNOR2_X1 U1005 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1006 ( .A(n907), .B(n906), .Z(n909) );
  XNOR2_X1 U1007 ( .A(G2443), .B(G2451), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  NAND2_X1 U1010 ( .A1(n912), .A2(G14), .ZN(n917) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n917), .ZN(n913) );
  NOR2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  INV_X1 U1017 ( .A(n917), .ZN(G401) );
  XOR2_X1 U1018 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n1029) );
  XNOR2_X1 U1019 ( .A(KEYINPUT119), .B(G2090), .ZN(n918) );
  XNOR2_X1 U1020 ( .A(n918), .B(G35), .ZN(n935) );
  XNOR2_X1 U1021 ( .A(G2084), .B(G34), .ZN(n919) );
  XNOR2_X1 U1022 ( .A(n919), .B(KEYINPUT54), .ZN(n933) );
  XOR2_X1 U1023 ( .A(G25), .B(G1991), .Z(n920) );
  NAND2_X1 U1024 ( .A1(n920), .A2(G28), .ZN(n930) );
  XNOR2_X1 U1025 ( .A(G2067), .B(G26), .ZN(n922) );
  XNOR2_X1 U1026 ( .A(G2072), .B(G33), .ZN(n921) );
  NOR2_X1 U1027 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1028 ( .A(KEYINPUT120), .B(n923), .ZN(n928) );
  XOR2_X1 U1029 ( .A(n924), .B(G27), .Z(n926) );
  XNOR2_X1 U1030 ( .A(G1996), .B(G32), .ZN(n925) );
  NOR2_X1 U1031 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1032 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1033 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1034 ( .A(n931), .B(KEYINPUT53), .ZN(n932) );
  NOR2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(n1029), .B(n936), .ZN(n938) );
  INV_X1 U1038 ( .A(G29), .ZN(n937) );
  NAND2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1040 ( .A1(G11), .A2(n939), .ZN(n994) );
  XNOR2_X1 U1041 ( .A(G1348), .B(n940), .ZN(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n954) );
  XNOR2_X1 U1043 ( .A(G171), .B(G1961), .ZN(n946) );
  INV_X1 U1044 ( .A(n943), .ZN(n944) );
  XNOR2_X1 U1045 ( .A(n944), .B(KEYINPUT122), .ZN(n945) );
  NAND2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(n948) );
  XNOR2_X1 U1047 ( .A(G1956), .B(G299), .ZN(n947) );
  NOR2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n950) );
  NAND2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n952) );
  XNOR2_X1 U1050 ( .A(G1971), .B(G303), .ZN(n951) );
  NOR2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n958) );
  XOR2_X1 U1053 ( .A(G1341), .B(n955), .Z(n956) );
  XNOR2_X1 U1054 ( .A(KEYINPUT123), .B(n956), .ZN(n957) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1056 ( .A(KEYINPUT124), .B(n959), .Z(n965) );
  XOR2_X1 U1057 ( .A(G168), .B(G1966), .Z(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1059 ( .A(KEYINPUT57), .B(n962), .Z(n963) );
  XNOR2_X1 U1060 ( .A(KEYINPUT121), .B(n963), .ZN(n964) );
  NOR2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n997) );
  NOR2_X1 U1062 ( .A1(KEYINPUT56), .A2(n997), .ZN(n991) );
  XNOR2_X1 U1063 ( .A(n966), .B(G5), .ZN(n988) );
  XOR2_X1 U1064 ( .A(G1966), .B(G21), .Z(n979) );
  XOR2_X1 U1065 ( .A(G4), .B(KEYINPUT126), .Z(n968) );
  XNOR2_X1 U1066 ( .A(G1348), .B(KEYINPUT59), .ZN(n967) );
  XNOR2_X1 U1067 ( .A(n968), .B(n967), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(G20), .B(n969), .ZN(n973) );
  XNOR2_X1 U1069 ( .A(G1341), .B(G19), .ZN(n971) );
  XNOR2_X1 U1070 ( .A(G6), .B(G1981), .ZN(n970) );
  NOR2_X1 U1071 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1072 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1073 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1074 ( .A(KEYINPUT60), .B(n976), .Z(n977) );
  XNOR2_X1 U1075 ( .A(KEYINPUT127), .B(n977), .ZN(n978) );
  NAND2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(G1971), .B(G22), .ZN(n981) );
  XNOR2_X1 U1078 ( .A(G23), .B(G1976), .ZN(n980) );
  NOR2_X1 U1079 ( .A1(n981), .A2(n980), .ZN(n983) );
  XOR2_X1 U1080 ( .A(G1986), .B(G24), .Z(n982) );
  NAND2_X1 U1081 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1082 ( .A(KEYINPUT58), .B(n984), .ZN(n985) );
  NOR2_X1 U1083 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1084 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1085 ( .A(n989), .B(KEYINPUT61), .ZN(n995) );
  NOR2_X1 U1086 ( .A1(KEYINPUT125), .A2(n995), .ZN(n990) );
  NOR2_X1 U1087 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1088 ( .A1(G16), .A2(n992), .ZN(n993) );
  NOR2_X1 U1089 ( .A1(n994), .A2(n993), .ZN(n1003) );
  INV_X1 U1090 ( .A(n995), .ZN(n996) );
  NAND2_X1 U1091 ( .A1(KEYINPUT125), .A2(n996), .ZN(n1000) );
  INV_X1 U1092 ( .A(n997), .ZN(n998) );
  NAND2_X1 U1093 ( .A1(KEYINPUT56), .A2(n998), .ZN(n999) );
  NAND2_X1 U1094 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1095 ( .A1(n1001), .A2(G16), .ZN(n1002) );
  AND2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1033) );
  XOR2_X1 U1097 ( .A(G2090), .B(G162), .Z(n1004) );
  NOR2_X1 U1098 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1099 ( .A(KEYINPUT51), .B(n1006), .Z(n1015) );
  XNOR2_X1 U1100 ( .A(G160), .B(G2084), .ZN(n1008) );
  NAND2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1103 ( .A(KEYINPUT115), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1107 ( .A(KEYINPUT116), .B(n1018), .Z(n1024) );
  XOR2_X1 U1108 ( .A(G2072), .B(n1019), .Z(n1021) );
  XOR2_X1 U1109 ( .A(G164), .B(G2078), .Z(n1020) );
  NOR2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1111 ( .A(KEYINPUT50), .B(n1022), .Z(n1023) );
  NOR2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1114 ( .A(n1027), .B(KEYINPUT117), .ZN(n1028) );
  XNOR2_X1 U1115 ( .A(KEYINPUT52), .B(n1028), .ZN(n1030) );
  NAND2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1117 ( .A1(n1031), .A2(G29), .ZN(n1032) );
  NAND2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1034), .Z(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

