//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n434, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n549, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1226, new_n1227,
    new_n1228, new_n1229;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(new_n434));
  INV_X1    g009(.A(new_n434), .ZN(G218));
  INV_X1    g010(.A(G132), .ZN(G219));
  XNOR2_X1  g011(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G221), .A3(G219), .A4(G220), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n463), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n468), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n471), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n467), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n478), .A2(new_n479), .A3(G124), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  OAI21_X1  g058(.A(KEYINPUT69), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n468), .A2(G136), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n477), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n480), .A2(new_n484), .A3(new_n485), .A4(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND4_X1  g064(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n477), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n481), .A2(G138), .A3(new_n477), .A4(new_n492), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G114), .C2(new_n477), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n464), .A2(new_n466), .A3(G126), .A4(G2105), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n508), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n514), .A2(new_n507), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n510), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n514), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G62), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n503), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n518), .A2(new_n522), .ZN(G166));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n514), .B(new_n524), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n515), .A2(G89), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n509), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n526), .A2(new_n531), .ZN(G168));
  AOI22_X1  g107(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n503), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n509), .A2(G52), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n516), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G171));
  AOI22_X1  g113(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n503), .ZN(new_n540));
  XOR2_X1   g115(.A(KEYINPUT73), .B(G81), .Z(new_n541));
  AOI22_X1  g116(.A1(new_n515), .A2(new_n541), .B1(new_n509), .B2(G43), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT74), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  XOR2_X1   g126(.A(new_n551), .B(KEYINPUT75), .Z(G188));
  INV_X1    g127(.A(new_n507), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n553), .A2(G53), .A3(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT77), .ZN(new_n557));
  XOR2_X1   g132(.A(KEYINPUT76), .B(KEYINPUT9), .Z(new_n558));
  NAND3_X1  g133(.A1(new_n509), .A2(G53), .A3(new_n558), .ZN(new_n559));
  AND3_X1   g134(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n557), .B1(new_n556), .B2(new_n559), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n514), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT78), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n565), .A2(new_n568), .A3(G651), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n567), .A2(new_n569), .B1(G91), .B2(new_n515), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n562), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  INV_X1    g148(.A(G166), .ZN(G303));
  NAND2_X1  g149(.A1(new_n509), .A2(G49), .ZN(new_n575));
  INV_X1    g150(.A(G87), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n516), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n525), .A2(G74), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n577), .B1(new_n579), .B2(G651), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(new_n515), .A2(G86), .ZN(new_n582));
  INV_X1    g157(.A(G48), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n553), .A2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n519), .A2(G61), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n503), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n585), .A2(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n503), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n509), .A2(G47), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n516), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G290));
  XOR2_X1   g171(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n516), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n514), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(new_n509), .B2(G54), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n515), .A2(G92), .A3(new_n597), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n600), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G171), .B2(new_n608), .ZN(G284));
  OAI21_X1  g185(.A(new_n609), .B1(G171), .B2(new_n608), .ZN(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  INV_X1    g187(.A(G299), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT80), .Z(G297));
  XNOR2_X1  g190(.A(new_n614), .B(KEYINPUT81), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n606), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n543), .A2(new_n608), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n607), .A2(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n608), .B2(new_n620), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n481), .A2(new_n469), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT82), .B(G2100), .Z(new_n626));
  INV_X1    g201(.A(KEYINPUT83), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n625), .B(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(G123), .ZN(new_n630));
  OR3_X1    g205(.A1(new_n482), .A2(KEYINPUT84), .A3(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(KEYINPUT84), .B1(new_n482), .B2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n468), .A2(G135), .ZN(new_n633));
  OR2_X1    g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G111), .C2(new_n477), .ZN(new_n635));
  NAND4_X1  g210(.A1(new_n631), .A2(new_n632), .A3(new_n633), .A4(new_n635), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n636), .A2(G2096), .B1(new_n627), .B2(new_n626), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n629), .B(new_n637), .C1(G2096), .C2(new_n636), .ZN(G156));
  XNOR2_X1  g213(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n639));
  INV_X1    g214(.A(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  INV_X1    g220(.A(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2427), .B(G2430), .Z(new_n648));
  OAI21_X1  g223(.A(KEYINPUT14), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT86), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI211_X1 g226(.A(KEYINPUT86), .B(KEYINPUT14), .C1(new_n647), .C2(new_n648), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(G1341), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n647), .A2(new_n648), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n654), .B1(new_n653), .B2(new_n655), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n644), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n660), .A2(new_n656), .A3(new_n643), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n659), .A2(new_n661), .A3(new_n663), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(G14), .A3(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(G2067), .B(G2678), .Z(new_n669));
  XNOR2_X1  g244(.A(G2084), .B(G2090), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2072), .B(G2078), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT18), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n669), .A2(new_n670), .ZN(new_n675));
  AND3_X1   g250(.A1(new_n675), .A2(KEYINPUT17), .A3(new_n672), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n672), .B1(new_n675), .B2(KEYINPUT17), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n676), .A2(new_n677), .A3(new_n671), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2096), .B(G2100), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1961), .B(G1966), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  INV_X1    g266(.A(new_n686), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(new_n688), .ZN(new_n693));
  INV_X1    g268(.A(new_n689), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n692), .A2(new_n693), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT88), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G1991), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n696), .A2(new_n698), .ZN(new_n701));
  INV_X1    g276(.A(G1991), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AND3_X1   g278(.A1(new_n700), .A2(G1996), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(G1996), .B1(new_n700), .B2(new_n703), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1981), .B(G1986), .ZN(new_n706));
  NOR3_X1   g281(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n706), .ZN(new_n708));
  INV_X1    g283(.A(G1996), .ZN(new_n709));
  INV_X1    g284(.A(new_n703), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n701), .A2(new_n702), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n700), .A2(G1996), .A3(new_n703), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n708), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n683), .B1(new_n707), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n706), .B1(new_n704), .B2(new_n705), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n712), .A2(new_n708), .A3(new_n713), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n716), .A2(new_n682), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n715), .A2(new_n718), .ZN(G229));
  AND2_X1   g294(.A1(KEYINPUT90), .A2(G16), .ZN(new_n720));
  NOR2_X1   g295(.A1(KEYINPUT90), .A2(G16), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(G24), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n595), .B2(new_n722), .ZN(new_n724));
  INV_X1    g299(.A(G1986), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G25), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n478), .A2(G119), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n468), .A2(G131), .ZN(new_n730));
  OR2_X1    g305(.A1(G95), .A2(G2105), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n731), .B(G2104), .C1(G107), .C2(new_n477), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n728), .B1(new_n734), .B2(new_n727), .ZN(new_n735));
  MUX2_X1   g310(.A(new_n728), .B(new_n735), .S(KEYINPUT89), .Z(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT35), .B(G1991), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n736), .B(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G16), .A2(G23), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n580), .B2(G16), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT33), .B(G1976), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n722), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G22), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G166), .B2(new_n744), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1971), .ZN(new_n747));
  INV_X1    g322(.A(G16), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G6), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n585), .A2(new_n588), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(new_n748), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT32), .B(G1981), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT91), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n751), .B(new_n753), .Z(new_n754));
  NOR3_X1   g329(.A1(new_n743), .A2(new_n747), .A3(new_n754), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n755), .A2(KEYINPUT34), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n755), .A2(KEYINPUT34), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n726), .B(new_n739), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT36), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G28), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(KEYINPUT30), .ZN(new_n762));
  AOI21_X1  g337(.A(G29), .B1(new_n761), .B2(KEYINPUT30), .ZN(new_n763));
  OR2_X1    g338(.A1(KEYINPUT31), .A2(G11), .ZN(new_n764));
  NAND2_X1  g339(.A1(KEYINPUT31), .A2(G11), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n762), .A2(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n636), .B2(new_n727), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT24), .ZN(new_n768));
  INV_X1    g343(.A(G34), .ZN(new_n769));
  AOI21_X1  g344(.A(G29), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n768), .B2(new_n769), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G160), .B2(new_n727), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n772), .A2(G2084), .ZN(new_n773));
  NAND2_X1  g348(.A1(G168), .A2(G16), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G16), .B2(G21), .ZN(new_n775));
  INV_X1    g350(.A(G1966), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n767), .B(new_n773), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  OAI22_X1  g352(.A1(KEYINPUT96), .A2(G2072), .B1(G29), .B2(G33), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n481), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(new_n477), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n468), .A2(G139), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n469), .A2(G103), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(KEYINPUT25), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(KEYINPUT25), .ZN(new_n784));
  AND4_X1   g359(.A1(new_n780), .A2(new_n781), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n778), .B1(new_n785), .B2(G29), .ZN(new_n786));
  NAND2_X1  g361(.A1(KEYINPUT96), .A2(G2072), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n777), .B(new_n788), .C1(G2084), .C2(new_n772), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n775), .A2(new_n776), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n727), .A2(G27), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G164), .B2(new_n727), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2078), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n789), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT92), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n744), .A2(G19), .ZN(new_n796));
  AOI211_X1 g371(.A(new_n795), .B(new_n796), .C1(new_n543), .C2(new_n722), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n795), .B2(new_n796), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(new_n654), .ZN(new_n799));
  OAI21_X1  g374(.A(KEYINPUT93), .B1(G104), .B2(G2105), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NOR3_X1   g376(.A1(KEYINPUT93), .A2(G104), .A3(G2105), .ZN(new_n802));
  OAI221_X1 g377(.A(G2104), .B1(G116), .B2(new_n477), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(KEYINPUT94), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(KEYINPUT94), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n468), .ZN(new_n807));
  INV_X1    g382(.A(G140), .ZN(new_n808));
  INV_X1    g383(.A(G128), .ZN(new_n809));
  OAI22_X1  g384(.A1(new_n807), .A2(new_n808), .B1(new_n809), .B2(new_n482), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(new_n727), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT95), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n727), .A2(G26), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT28), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G2067), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n794), .A2(new_n799), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n727), .A2(G35), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G162), .B2(new_n727), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT29), .Z(new_n822));
  INV_X1    g397(.A(G2090), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n824), .A2(KEYINPUT99), .B1(KEYINPUT98), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n744), .A2(G20), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT23), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n613), .B2(new_n748), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT100), .B(G1956), .Z(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n748), .A2(G4), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n606), .B2(new_n748), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(G1348), .ZN(new_n834));
  NOR2_X1   g409(.A1(G29), .A2(G32), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n478), .A2(G129), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n468), .A2(G141), .ZN(new_n837));
  NAND3_X1  g412(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT26), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n840), .A2(new_n841), .B1(G105), .B2(new_n469), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n836), .A2(new_n837), .A3(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n843), .A2(KEYINPUT97), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(KEYINPUT97), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n835), .B1(new_n847), .B2(G29), .ZN(new_n848));
  XOR2_X1   g423(.A(KEYINPUT27), .B(G1996), .Z(new_n849));
  AOI21_X1  g424(.A(new_n834), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(G1348), .B2(new_n833), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n826), .A2(new_n831), .A3(new_n850), .A4(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(G5), .A2(G16), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(G171), .B2(G16), .ZN(new_n855));
  INV_X1    g430(.A(G1961), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n824), .B2(KEYINPUT99), .ZN(new_n858));
  OAI22_X1  g433(.A1(new_n825), .A2(KEYINPUT98), .B1(new_n829), .B2(new_n830), .ZN(new_n859));
  NOR4_X1   g434(.A1(new_n819), .A2(new_n853), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n760), .A2(new_n861), .ZN(G311));
  OAI21_X1  g437(.A(KEYINPUT101), .B1(new_n760), .B2(new_n861), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n759), .A2(new_n864), .A3(new_n860), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(G150));
  NAND2_X1  g441(.A1(new_n525), .A2(G67), .ZN(new_n867));
  NAND2_X1  g442(.A1(G80), .A2(G543), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n503), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n509), .A2(G55), .ZN(new_n870));
  INV_X1    g445(.A(G93), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n870), .B1(new_n516), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(G860), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT37), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n606), .A2(G559), .ZN(new_n877));
  XOR2_X1   g452(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n878));
  XOR2_X1   g453(.A(new_n877), .B(new_n878), .Z(new_n879));
  NAND2_X1  g454(.A1(new_n543), .A2(new_n873), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n540), .B(new_n542), .C1(new_n869), .C2(new_n872), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n874), .B1(new_n879), .B2(new_n882), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n876), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT102), .ZN(G145));
  XNOR2_X1  g461(.A(new_n488), .B(new_n475), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n636), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n844), .A2(new_n785), .A3(new_n845), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n785), .B1(new_n844), .B2(new_n845), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n811), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n494), .A2(new_n495), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n893), .B1(new_n494), .B2(new_n495), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n500), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n785), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n846), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n811), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n899), .A2(new_n900), .A3(new_n889), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n892), .A2(new_n897), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n897), .B1(new_n892), .B2(new_n901), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n468), .A2(G142), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n477), .A2(G118), .ZN(new_n906));
  OAI21_X1  g481(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n908), .B1(G130), .B2(new_n478), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(new_n624), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(new_n733), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n903), .A2(new_n904), .A3(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n910), .B(new_n734), .ZN(new_n913));
  INV_X1    g488(.A(new_n901), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n900), .B1(new_n899), .B2(new_n889), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n896), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n913), .B1(new_n916), .B2(new_n902), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n888), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(G37), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n911), .B1(new_n903), .B2(new_n904), .ZN(new_n921));
  XOR2_X1   g496(.A(new_n888), .B(KEYINPUT106), .Z(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT104), .B1(new_n903), .B2(new_n904), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n916), .A2(new_n925), .A3(new_n902), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n911), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n923), .B1(new_n927), .B2(KEYINPUT105), .ZN(new_n928));
  INV_X1    g503(.A(new_n926), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n925), .B1(new_n916), .B2(new_n902), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n913), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n920), .B1(new_n928), .B2(new_n933), .ZN(new_n934));
  XOR2_X1   g509(.A(new_n934), .B(KEYINPUT40), .Z(G395));
  INV_X1    g510(.A(KEYINPUT42), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n882), .B(KEYINPUT107), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(G559), .B2(new_n607), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n882), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n620), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n613), .A2(new_n607), .ZN(new_n942));
  NAND2_X1  g517(.A1(G299), .A2(new_n606), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT41), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n942), .A2(new_n943), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n938), .A2(new_n941), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n944), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n952), .B1(new_n938), .B2(new_n941), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n936), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n938), .A2(new_n941), .ZN(new_n955));
  OAI211_X1 g530(.A(KEYINPUT42), .B(new_n950), .C1(new_n955), .C2(new_n952), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n750), .B(G166), .ZN(new_n957));
  NAND2_X1  g532(.A1(G290), .A2(new_n580), .ZN(new_n958));
  NAND2_X1  g533(.A1(G288), .A2(new_n595), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n957), .A3(new_n959), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(KEYINPUT109), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n954), .A2(new_n956), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n964), .B1(new_n954), .B2(new_n956), .ZN(new_n966));
  OAI21_X1  g541(.A(G868), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(G868), .B2(new_n873), .ZN(G295));
  OAI21_X1  g543(.A(new_n967), .B1(G868), .B2(new_n873), .ZN(G331));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n970));
  INV_X1    g545(.A(new_n962), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n970), .B1(new_n971), .B2(new_n960), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n961), .A2(KEYINPUT110), .A3(new_n962), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(G301), .A2(G168), .ZN(new_n975));
  NAND2_X1  g550(.A1(G171), .A2(G286), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n882), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n975), .A2(new_n880), .A3(new_n881), .A4(new_n976), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n947), .B1(new_n942), .B2(new_n943), .ZN(new_n981));
  OAI22_X1  g556(.A1(new_n981), .A2(KEYINPUT111), .B1(new_n944), .B2(new_n945), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n981), .A2(KEYINPUT111), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n978), .A2(new_n944), .A3(new_n979), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n974), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n949), .A2(new_n980), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n988), .A2(new_n963), .A3(new_n985), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n989), .A2(new_n919), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n987), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n974), .B1(new_n988), .B2(new_n985), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n989), .A2(new_n919), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT43), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n993), .A2(new_n994), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n987), .A2(new_n990), .A3(KEYINPUT112), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(new_n986), .B2(new_n994), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1000), .B1(new_n1004), .B2(KEYINPUT43), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n998), .B1(new_n1005), .B2(new_n997), .ZN(G397));
  INV_X1    g581(.A(G1384), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT45), .B1(new_n896), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n470), .A2(G40), .A3(new_n474), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n811), .B(G2067), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n847), .A2(new_n709), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n846), .A2(G1996), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n733), .B(new_n737), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1011), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1011), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n595), .B(G1986), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n1020), .B(KEYINPUT113), .Z(new_n1021));
  INV_X1    g596(.A(G40), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n1007), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(G160), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1008), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT119), .B1(new_n1025), .B2(G1966), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1023), .A2(G160), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n496), .A2(KEYINPUT103), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n494), .A2(new_n495), .A3(new_n893), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1384), .B1(new_n1030), .B2(new_n500), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1027), .B(G40), .C1(new_n1031), .C2(KEYINPUT45), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(new_n1033), .A3(new_n776), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT50), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n896), .A2(new_n1035), .A3(new_n1007), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n501), .A2(new_n1007), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1010), .B1(new_n1037), .B2(KEYINPUT50), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  OR2_X1    g614(.A1(new_n1039), .A2(G2084), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1026), .A2(new_n1034), .A3(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1041), .A2(G8), .A3(G168), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n896), .A2(KEYINPUT45), .A3(new_n1007), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT45), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1010), .B1(new_n1037), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1971), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(KEYINPUT114), .A3(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1036), .A2(new_n1038), .A3(new_n823), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT114), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1043), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1054), .B1(new_n1055), .B2(G1971), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1056), .A2(KEYINPUT115), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1057));
  NAND2_X1  g632(.A1(G303), .A2(G8), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT117), .ZN(new_n1061));
  NAND4_X1  g636(.A1(G303), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1058), .A2(new_n1065), .A3(new_n1059), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .A4(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1053), .A2(new_n1057), .A3(G8), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1067), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1010), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1037), .B2(KEYINPUT50), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1070), .A2(G2090), .A3(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1055), .A2(G1971), .ZN(new_n1074));
  OAI21_X1  g649(.A(G8), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1069), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n580), .A2(G1976), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1031), .A2(new_n1071), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(G8), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n580), .B2(G1976), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1079), .A2(KEYINPUT52), .ZN(new_n1083));
  NAND2_X1  g658(.A1(G305), .A2(G1981), .ZN(new_n1084));
  INV_X1    g659(.A(G1981), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n750), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT49), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1084), .A2(KEYINPUT49), .A3(new_n1086), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1089), .A2(G8), .A3(new_n1078), .A4(new_n1090), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1082), .A2(new_n1083), .A3(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1042), .A2(new_n1068), .A3(new_n1076), .A4(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT63), .B1(new_n1093), .B2(KEYINPUT120), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1068), .A2(new_n1092), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(new_n1076), .A4(new_n1042), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1053), .A2(G8), .A3(new_n1057), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n1069), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1095), .A2(KEYINPUT63), .A3(new_n1042), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1103), .B(G8), .C1(new_n1041), .C2(G286), .ZN(new_n1104));
  INV_X1    g679(.A(G8), .ZN(new_n1105));
  NOR2_X1   g680(.A1(G168), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1041), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  AOI211_X1 g683(.A(new_n1103), .B(new_n1106), .C1(new_n1041), .C2(G8), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1036), .A2(new_n1038), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1111), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n856), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1047), .B2(G2078), .ZN(new_n1116));
  NAND2_X1  g691(.A1(G301), .A2(KEYINPUT54), .ZN(new_n1117));
  OR3_X1    g692(.A1(new_n534), .A2(KEYINPUT54), .A3(new_n537), .ZN(new_n1118));
  AND4_X1   g693(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n474), .B1(new_n470), .B2(KEYINPUT123), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1120), .B1(KEYINPUT123), .B2(new_n470), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1009), .A2(G40), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT124), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1115), .A2(G2078), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1009), .A2(new_n1125), .A3(G40), .A4(new_n1121), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1123), .A2(new_n1044), .A3(new_n1124), .A4(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(G2078), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1025), .A2(KEYINPUT53), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1114), .A2(new_n1129), .A3(new_n1116), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1119), .A2(new_n1127), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1132), .A2(new_n1076), .A3(new_n1068), .A4(new_n1092), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1110), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(G1956), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT56), .B(G2072), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1055), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT57), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n556), .A2(new_n1140), .A3(new_n559), .ZN(new_n1141));
  AOI22_X1  g716(.A1(G299), .A2(KEYINPUT57), .B1(new_n570), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1136), .A2(new_n1138), .A3(new_n1142), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1145), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT58), .B(G1341), .Z(new_n1149));
  NAND2_X1  g724(.A1(new_n1078), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(G1996), .B2(new_n1047), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n544), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n1147), .A2(new_n1148), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n640), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1078), .A2(G2067), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT60), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1162), .B1(new_n1163), .B2(new_n606), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT60), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1165), .A2(KEYINPUT122), .A3(new_n607), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1161), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1163), .A2(new_n1162), .A3(new_n606), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1161), .ZN(new_n1169));
  OAI21_X1  g744(.A(KEYINPUT122), .B1(new_n1165), .B2(new_n607), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1155), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1146), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1159), .A2(new_n606), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1173), .B1(new_n1174), .B2(new_n1144), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1134), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(G288), .A2(G1976), .ZN(new_n1177));
  AOI22_X1  g752(.A1(new_n1091), .A2(new_n1177), .B1(new_n1085), .B2(new_n750), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT118), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n1180), .A2(G8), .A3(new_n1078), .ZN(new_n1181));
  OR2_X1    g756(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1068), .ZN(new_n1183));
  AOI22_X1  g758(.A1(new_n1181), .A2(new_n1182), .B1(new_n1183), .B2(new_n1092), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1102), .A2(new_n1176), .A3(new_n1184), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1130), .A2(G171), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1068), .A2(new_n1186), .A3(new_n1092), .A4(new_n1076), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1041), .A2(G8), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1106), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1188), .A2(KEYINPUT51), .A3(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1190), .A2(new_n1107), .A3(new_n1104), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1187), .B1(new_n1191), .B2(KEYINPUT62), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT62), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1190), .A2(new_n1193), .A3(new_n1107), .A4(new_n1104), .ZN(new_n1194));
  AOI21_X1  g769(.A(KEYINPUT125), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(KEYINPUT62), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1187), .ZN(new_n1197));
  AND4_X1   g772(.A1(KEYINPUT125), .A2(new_n1196), .A3(new_n1194), .A4(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1195), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1021), .B1(new_n1185), .B2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1011), .A2(KEYINPUT48), .A3(new_n725), .A4(new_n595), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT48), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n595), .A2(new_n725), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1202), .B1(new_n1018), .B2(new_n1203), .ZN(new_n1204));
  AND3_X1   g779(.A1(new_n1017), .A2(new_n1201), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1018), .B1(new_n847), .B2(new_n1012), .ZN(new_n1206));
  AND3_X1   g781(.A1(new_n1011), .A2(KEYINPUT46), .A3(new_n709), .ZN(new_n1207));
  AOI21_X1  g782(.A(KEYINPUT46), .B1(new_n1011), .B2(new_n709), .ZN(new_n1208));
  NOR3_X1   g783(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT47), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n734), .A2(new_n738), .ZN(new_n1211));
  OAI22_X1  g786(.A1(new_n1015), .A2(new_n1211), .B1(G2067), .B2(new_n900), .ZN(new_n1212));
  AOI211_X1 g787(.A(new_n1205), .B(new_n1210), .C1(new_n1011), .C2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1200), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g789(.A(KEYINPUT126), .ZN(new_n1216));
  NOR2_X1   g790(.A1(new_n461), .A2(G227), .ZN(new_n1217));
  NAND3_X1  g791(.A1(new_n667), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g792(.A(new_n1218), .ZN(new_n1219));
  AOI21_X1  g793(.A(new_n1216), .B1(new_n667), .B2(new_n1217), .ZN(new_n1220));
  OAI211_X1 g794(.A(new_n715), .B(new_n718), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1221));
  NOR2_X1   g795(.A1(new_n934), .A2(new_n1221), .ZN(new_n1222));
  AND3_X1   g796(.A1(new_n1222), .A2(KEYINPUT127), .A3(new_n996), .ZN(new_n1223));
  AOI21_X1  g797(.A(KEYINPUT127), .B1(new_n1222), .B2(new_n996), .ZN(new_n1224));
  NOR2_X1   g798(.A1(new_n1223), .A2(new_n1224), .ZN(G308));
  NAND2_X1  g799(.A1(new_n1222), .A2(new_n996), .ZN(new_n1226));
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n1227));
  NAND2_X1  g801(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g802(.A1(new_n1222), .A2(new_n996), .A3(KEYINPUT127), .ZN(new_n1229));
  NAND2_X1  g803(.A1(new_n1228), .A2(new_n1229), .ZN(G225));
endmodule


