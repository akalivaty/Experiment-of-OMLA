//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957;
  AND2_X1   g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203));
  XOR2_X1   g002(.A(G113gat), .B(G120gat), .Z(new_n204));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT68), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(KEYINPUT69), .B(KEYINPUT1), .Z(new_n209));
  NAND3_X1  g008(.A1(new_n204), .A2(new_n209), .A3(new_n203), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT70), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n216), .B2(KEYINPUT26), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT26), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n217), .A2(KEYINPUT67), .B1(new_n218), .B2(new_n213), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n214), .B(new_n220), .C1(new_n216), .C2(KEYINPUT26), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(KEYINPUT27), .B(G183gat), .Z(new_n225));
  INV_X1    g024(.A(KEYINPUT28), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n225), .A2(new_n226), .A3(G190gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT27), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G183gat), .ZN(new_n229));
  AOI21_X1  g028(.A(G190gat), .B1(new_n229), .B2(KEYINPUT66), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT65), .B(G183gat), .ZN(new_n231));
  OAI221_X1 g030(.A(new_n230), .B1(KEYINPUT66), .B2(new_n229), .C1(new_n228), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n227), .B1(new_n232), .B2(new_n226), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n224), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT25), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n223), .A2(KEYINPUT24), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT24), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(G183gat), .A3(G190gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(G183gat), .B2(G190gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n213), .B1(KEYINPUT23), .B2(new_n215), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT64), .B(G176gat), .ZN(new_n243));
  INV_X1    g042(.A(G169gat), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n244), .A2(KEYINPUT23), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n240), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G176gat), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n249), .A2(new_n235), .A3(new_n241), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n239), .B1(new_n231), .B2(G190gat), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n235), .A2(new_n247), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n212), .B1(new_n234), .B2(new_n252), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n219), .A2(new_n221), .B1(G183gat), .B2(G190gat), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n232), .A2(new_n226), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n255), .B2(new_n227), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n206), .B(KEYINPUT68), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n210), .B(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n252), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n256), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n202), .B1(new_n253), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(KEYINPUT73), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n253), .A2(new_n202), .A3(new_n262), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT32), .ZN(new_n267));
  XNOR2_X1  g066(.A(G15gat), .B(G43gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT72), .ZN(new_n269));
  XNOR2_X1  g068(.A(G71gat), .B(G99gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT33), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n273), .B1(new_n266), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n266), .A2(new_n273), .A3(new_n274), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n272), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n271), .A2(KEYINPUT33), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n266), .A2(KEYINPUT32), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n278), .A2(KEYINPUT34), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT34), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n266), .A2(new_n273), .A3(new_n274), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n267), .B(new_n271), .C1(new_n284), .C2(new_n275), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n283), .B1(new_n285), .B2(new_n280), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n265), .B1(new_n282), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT34), .B1(new_n278), .B2(new_n281), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(new_n283), .A3(new_n280), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n264), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G1gat), .B(G29gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(KEYINPUT0), .ZN(new_n293));
  XNOR2_X1  g092(.A(G57gat), .B(G85gat), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n293), .B(new_n294), .Z(new_n295));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n257), .A2(new_n259), .A3(KEYINPUT78), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT78), .B1(new_n257), .B2(new_n259), .ZN(new_n299));
  XNOR2_X1  g098(.A(G141gat), .B(G148gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n300), .B1(KEYINPUT2), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT76), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n303), .B1(new_n304), .B2(new_n301), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n305), .B1(new_n304), .B2(new_n301), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G155gat), .B(G162gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n302), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NOR3_X1   g112(.A1(new_n298), .A2(new_n299), .A3(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n260), .A2(new_n312), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n297), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n298), .A2(new_n299), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n312), .B(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT4), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n212), .A2(new_n320), .A3(new_n313), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT4), .B1(new_n260), .B2(new_n312), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n317), .A2(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n316), .A2(KEYINPUT5), .B1(new_n323), .B2(new_n296), .ZN(new_n324));
  INV_X1    g123(.A(new_n299), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n212), .A2(KEYINPUT78), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n319), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n321), .A2(new_n322), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT5), .ZN(new_n330));
  NOR3_X1   g129(.A1(new_n329), .A2(new_n330), .A3(new_n297), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n295), .B1(new_n324), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n295), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n323), .A2(KEYINPUT5), .A3(new_n296), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n326), .A2(new_n325), .A3(new_n312), .ZN(new_n335));
  INV_X1    g134(.A(new_n315), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n330), .B1(new_n337), .B2(new_n297), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n329), .A2(new_n297), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n333), .B(new_n334), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT6), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n332), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n324), .A2(new_n331), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n343), .A2(KEYINPUT6), .A3(new_n333), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G8gat), .B(G36gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(G64gat), .B(G92gat), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n346), .B(new_n347), .Z(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  AND2_X1   g148(.A1(G226gat), .A2(G233gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n350), .A2(KEYINPUT29), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n351), .B1(new_n234), .B2(new_n252), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT75), .B1(new_n234), .B2(new_n252), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n256), .A2(new_n261), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n353), .B1(new_n357), .B2(new_n350), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT74), .B(G197gat), .ZN(new_n359));
  INV_X1    g158(.A(G204gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT22), .ZN(new_n362));
  INV_X1    g161(.A(G211gat), .ZN(new_n363));
  INV_X1    g162(.A(G218gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(G211gat), .B(G218gat), .Z(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n367), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n361), .A2(new_n369), .A3(new_n365), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n358), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n354), .A2(new_n356), .A3(new_n351), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n256), .A2(new_n261), .A3(new_n350), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n349), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n376), .B(new_n348), .C1(new_n358), .C2(new_n372), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(KEYINPUT30), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n373), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT30), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n381), .A2(new_n382), .A3(new_n376), .A4(new_n348), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(G22gat), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT29), .B1(new_n368), .B2(new_n370), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n312), .B1(new_n387), .B2(KEYINPUT3), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT79), .ZN(new_n389));
  INV_X1    g188(.A(G228gat), .ZN(new_n390));
  INV_X1    g189(.A(G233gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n386), .B1(new_n389), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  AOI211_X1 g194(.A(G22gat), .B(new_n392), .C1(new_n388), .C2(KEYINPUT79), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT31), .B(G50gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n398), .B1(new_n394), .B2(new_n396), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT29), .B1(new_n313), .B2(new_n318), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n388), .B1(new_n371), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G78gat), .B(G106gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n402), .B(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n291), .A2(new_n345), .A3(new_n385), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT35), .ZN(new_n410));
  INV_X1    g209(.A(new_n345), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(new_n384), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n282), .A2(new_n286), .A3(new_n265), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n264), .B1(new_n288), .B2(new_n289), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n287), .A2(KEYINPUT82), .A3(new_n290), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n402), .B(new_n406), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n418), .A2(KEYINPUT35), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n412), .A2(new_n416), .A3(new_n417), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n410), .A2(new_n420), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n323), .A2(KEYINPUT39), .A3(new_n296), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(new_n333), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n329), .A2(new_n297), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n424), .B(KEYINPUT39), .C1(new_n297), .C2(new_n337), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n423), .A2(new_n425), .A3(KEYINPUT40), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT40), .B1(new_n423), .B2(new_n425), .ZN(new_n427));
  INV_X1    g226(.A(new_n340), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n418), .B1(new_n429), .B2(new_n384), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n342), .A2(new_n344), .A3(new_n379), .ZN(new_n431));
  XOR2_X1   g230(.A(KEYINPUT80), .B(KEYINPUT37), .Z(new_n432));
  OAI211_X1 g231(.A(new_n376), .B(new_n432), .C1(new_n358), .C2(new_n372), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT81), .ZN(new_n434));
  OR2_X1    g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n434), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n348), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT37), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n374), .A2(new_n375), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n438), .B1(new_n439), .B2(new_n371), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n358), .A2(new_n371), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT38), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n431), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT38), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT37), .B1(new_n373), .B2(new_n377), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n445), .B1(new_n437), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n430), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n385), .A2(new_n345), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n418), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n291), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT36), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT36), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n291), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n421), .B1(new_n451), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G190gat), .B(G218gat), .ZN(new_n458));
  AND2_X1   g257(.A1(G43gat), .A2(G50gat), .ZN(new_n459));
  NOR2_X1   g258(.A1(G43gat), .A2(G50gat), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT15), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT83), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT83), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n465), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT84), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT14), .ZN(new_n469));
  INV_X1    g268(.A(G29gat), .ZN(new_n470));
  INV_X1    g269(.A(G36gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n467), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(G29gat), .A2(G36gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n468), .B1(new_n467), .B2(new_n472), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n462), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OR4_X1    g276(.A1(KEYINPUT86), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n472), .A2(KEYINPUT86), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n467), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n461), .A2(new_n474), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT15), .ZN(new_n483));
  NAND2_X1  g282(.A1(G43gat), .A2(G50gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT85), .B(G50gat), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n483), .B(new_n484), .C1(new_n485), .C2(G43gat), .ZN(new_n486));
  AND4_X1   g285(.A1(KEYINPUT87), .A2(new_n480), .A3(new_n482), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n483), .ZN(new_n488));
  AND2_X1   g287(.A1(KEYINPUT85), .A2(G50gat), .ZN(new_n489));
  NOR2_X1   g288(.A1(KEYINPUT85), .A2(G50gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(G43gat), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n488), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n493), .A2(new_n481), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT87), .B1(new_n494), .B2(new_n480), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n477), .B(KEYINPUT17), .C1(new_n487), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(G99gat), .A2(G106gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT8), .ZN(new_n498));
  NAND2_X1  g297(.A1(G85gat), .A2(G92gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT7), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(G85gat), .ZN(new_n502));
  INV_X1    g301(.A(G92gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n498), .A2(new_n501), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  OR2_X1    g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n497), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g309(.A1(KEYINPUT8), .A2(new_n497), .B1(new_n502), .B2(new_n503), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n511), .A2(new_n508), .A3(new_n501), .A4(new_n505), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT93), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n510), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n506), .A2(new_n509), .A3(KEYINPUT93), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n482), .A2(new_n486), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n467), .A2(new_n479), .A3(new_n478), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n494), .A2(KEYINPUT87), .A3(new_n480), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n467), .A2(new_n472), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT84), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(new_n474), .A3(new_n473), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n520), .A2(new_n521), .B1(new_n524), .B2(new_n462), .ZN(new_n525));
  XOR2_X1   g324(.A(KEYINPUT88), .B(KEYINPUT17), .Z(new_n526));
  OAI211_X1 g325(.A(new_n496), .B(new_n516), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT94), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n477), .B1(new_n487), .B2(new_n495), .ZN(new_n530));
  INV_X1    g329(.A(new_n526), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n532), .A2(KEYINPUT94), .A3(new_n496), .A4(new_n516), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT41), .ZN(new_n535));
  NAND2_X1  g334(.A1(G232gat), .A2(G233gat), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n536), .B(KEYINPUT91), .Z(new_n537));
  OAI22_X1  g336(.A1(new_n525), .A2(new_n516), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n458), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n538), .B1(new_n529), .B2(new_n533), .ZN(new_n540));
  INV_X1    g339(.A(new_n458), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT95), .B1(new_n540), .B2(new_n541), .ZN(new_n543));
  XOR2_X1   g342(.A(G134gat), .B(G162gat), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT92), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n537), .A2(new_n535), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n539), .A2(new_n542), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n540), .A2(new_n541), .ZN(new_n549));
  AOI211_X1 g348(.A(new_n458), .B(new_n538), .C1(new_n529), .C2(new_n533), .ZN(new_n550));
  INV_X1    g349(.A(new_n547), .ZN(new_n551));
  NOR4_X1   g350(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT95), .A4(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(G71gat), .A2(G78gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(G71gat), .A2(G78gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G57gat), .B(G64gat), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G57gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(G64gat), .ZN(new_n561));
  INV_X1    g360(.A(G64gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(G57gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G71gat), .B(G78gat), .ZN(new_n565));
  INV_X1    g364(.A(new_n558), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n559), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT21), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(G127gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(G15gat), .B(G22gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT16), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n574), .B1(new_n575), .B2(G1gat), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n576), .B1(G1gat), .B2(new_n574), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(G8gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n579), .B1(new_n569), .B2(new_n568), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n573), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n582));
  INV_X1    g381(.A(G155gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G183gat), .B(G211gat), .Z(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n581), .B(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n553), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n496), .B(new_n579), .C1(new_n525), .C2(new_n526), .ZN(new_n590));
  NAND2_X1  g389(.A1(G229gat), .A2(G233gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n530), .A2(new_n578), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT18), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n591), .B(KEYINPUT13), .Z(new_n596));
  INV_X1    g395(.A(new_n592), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n530), .A2(new_n578), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n590), .A2(KEYINPUT18), .A3(new_n591), .A4(new_n592), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT89), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n601), .A2(KEYINPUT89), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G113gat), .B(G141gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(G197gat), .ZN(new_n606));
  XOR2_X1   g405(.A(KEYINPUT11), .B(G169gat), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n608), .B(KEYINPUT12), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n599), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n601), .A2(KEYINPUT89), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n601), .A2(KEYINPUT89), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n593), .A2(KEYINPUT90), .A3(new_n594), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT90), .B1(new_n593), .B2(new_n594), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI22_X1  g416(.A1(new_n604), .A2(new_n610), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n514), .A2(new_n515), .A3(new_n568), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n512), .A2(new_n559), .A3(new_n567), .ZN(new_n622));
  INV_X1    g421(.A(new_n497), .ZN(new_n623));
  NOR2_X1   g422(.A1(G99gat), .A2(G106gat), .ZN(new_n624));
  OAI21_X1  g423(.A(KEYINPUT96), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT96), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n507), .A2(new_n627), .A3(new_n497), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n506), .A2(new_n625), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n506), .A2(new_n625), .A3(new_n628), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT97), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n622), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT98), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n622), .A2(new_n631), .A3(KEYINPUT98), .A4(new_n629), .ZN(new_n635));
  AOI211_X1 g434(.A(KEYINPUT10), .B(new_n621), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT10), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n516), .A2(new_n637), .A3(new_n568), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n620), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n621), .B1(new_n634), .B2(new_n635), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n639), .B1(new_n620), .B2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G120gat), .B(G148gat), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT99), .ZN(new_n643));
  XNOR2_X1  g442(.A(G176gat), .B(G204gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n643), .B(new_n644), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n641), .A2(new_n646), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n589), .A2(new_n619), .A3(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n457), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n411), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G1gat), .ZN(G1324gat));
  INV_X1    g453(.A(KEYINPUT42), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n384), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT16), .B(G8gat), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT101), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n655), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(G8gat), .ZN(new_n662));
  OR3_X1    g461(.A1(new_n656), .A2(new_n655), .A3(new_n660), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(G1325gat));
  INV_X1    g463(.A(new_n652), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n453), .A2(new_n455), .ZN(new_n666));
  OAI21_X1  g465(.A(G15gat), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(G15gat), .ZN(new_n668));
  INV_X1    g467(.A(new_n416), .ZN(new_n669));
  INV_X1    g468(.A(new_n417), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n652), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n667), .A2(new_n672), .ZN(G1326gat));
  NAND2_X1  g472(.A1(new_n652), .A2(new_n418), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT43), .B(G22gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  INV_X1    g475(.A(new_n587), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n619), .A2(new_n677), .A3(new_n650), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n457), .A2(new_n553), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n470), .A3(new_n411), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT45), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n437), .A2(new_n446), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n443), .B(new_n431), .C1(new_n683), .C2(new_n445), .ZN(new_n684));
  AOI22_X1  g483(.A1(new_n684), .A2(new_n430), .B1(new_n449), .B2(new_n418), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n666), .A2(new_n685), .B1(new_n410), .B2(new_n420), .ZN(new_n686));
  INV_X1    g485(.A(new_n553), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n682), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n457), .A2(KEYINPUT44), .A3(new_n553), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n678), .B(KEYINPUT102), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(G29gat), .B1(new_n691), .B2(new_n345), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n681), .A2(new_n692), .ZN(G1328gat));
  NAND3_X1  g492(.A1(new_n679), .A2(new_n471), .A3(new_n384), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT46), .Z(new_n695));
  OAI21_X1  g494(.A(G36gat), .B1(new_n691), .B2(new_n385), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(G1329gat));
  NOR2_X1   g496(.A1(KEYINPUT104), .A2(KEYINPUT47), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n688), .A2(new_n456), .A3(new_n689), .A4(new_n690), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(G43gat), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n669), .A2(new_n670), .A3(G43gat), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n457), .A2(new_n553), .A3(new_n678), .A4(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(new_n707));
  AOI211_X1 g506(.A(new_n698), .B(new_n701), .C1(new_n703), .C2(new_n707), .ZN(new_n708));
  AND4_X1   g507(.A1(new_n699), .A2(new_n703), .A3(new_n707), .A4(new_n700), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(G1330gat));
  OAI21_X1  g509(.A(new_n485), .B1(new_n691), .B2(new_n408), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n408), .A2(new_n485), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT48), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n679), .A2(new_n712), .B1(KEYINPUT105), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n713), .A2(KEYINPUT105), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1331gat));
  INV_X1    g516(.A(new_n650), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n589), .A2(new_n618), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n457), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n345), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(new_n560), .ZN(G1332gat));
  NOR2_X1   g521(.A1(new_n720), .A2(new_n385), .ZN(new_n723));
  NOR2_X1   g522(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n724));
  AND2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(new_n723), .B2(new_n724), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n720), .B2(new_n666), .ZN(new_n728));
  INV_X1    g527(.A(G71gat), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n671), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n720), .B2(new_n730), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g531(.A1(new_n720), .A2(new_n408), .ZN(new_n733));
  XNOR2_X1  g532(.A(KEYINPUT106), .B(G78gat), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1335gat));
  NOR2_X1   g534(.A1(new_n618), .A2(new_n677), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n688), .A2(new_n650), .A3(new_n689), .A4(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G85gat), .B1(new_n737), .B2(new_n345), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n457), .A2(new_n553), .A3(new_n736), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT51), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n457), .A2(new_n741), .A3(new_n553), .A4(new_n736), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n740), .A2(new_n650), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n411), .A2(new_n502), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n738), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n738), .B(KEYINPUT107), .C1(new_n743), .C2(new_n744), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(G1336gat));
  OAI21_X1  g548(.A(G92gat), .B1(new_n737), .B2(new_n385), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n384), .A2(new_n503), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n743), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT52), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n750), .B(new_n754), .C1(new_n743), .C2(new_n751), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(G1337gat));
  OAI21_X1  g555(.A(G99gat), .B1(new_n737), .B2(new_n666), .ZN(new_n757));
  INV_X1    g556(.A(G99gat), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n671), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n759), .B2(new_n743), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT108), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n757), .B(new_n762), .C1(new_n743), .C2(new_n759), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(G1338gat));
  OAI21_X1  g563(.A(G106gat), .B1(new_n737), .B2(new_n408), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n408), .A2(G106gat), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n740), .A2(new_n650), .A3(new_n742), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n765), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n765), .A2(KEYINPUT109), .A3(new_n767), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT53), .B1(new_n765), .B2(KEYINPUT109), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(G1339gat));
  INV_X1    g571(.A(new_n620), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n634), .A2(new_n635), .ZN(new_n774));
  INV_X1    g573(.A(new_n621), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(new_n637), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n638), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n773), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n645), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n776), .A2(new_n773), .A3(new_n777), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n639), .A2(KEYINPUT54), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n780), .A2(new_n782), .A3(KEYINPUT55), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n780), .A2(new_n782), .A3(KEYINPUT111), .A4(KEYINPUT55), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT55), .B1(new_n780), .B2(new_n782), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n647), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n618), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n591), .B1(new_n590), .B2(new_n592), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n597), .A2(new_n598), .A3(new_n596), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n608), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  XOR2_X1   g592(.A(new_n793), .B(KEYINPUT112), .Z(new_n794));
  OR2_X1    g593(.A1(new_n614), .A2(new_n617), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n795), .A3(new_n650), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n553), .B1(new_n790), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n539), .A2(new_n542), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n543), .A2(new_n547), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n539), .A2(new_n543), .A3(new_n542), .A4(new_n547), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n787), .A2(new_n800), .A3(new_n801), .A4(new_n789), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n794), .A2(new_n795), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n587), .B1(new_n797), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n588), .A2(new_n619), .A3(new_n718), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n345), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n452), .A2(new_n384), .A3(new_n418), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(G113gat), .B1(new_n810), .B2(new_n618), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n418), .B1(new_n805), .B2(new_n806), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n345), .A2(new_n384), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n671), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n618), .A2(G113gat), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n811), .B1(new_n816), .B2(new_n817), .ZN(G1340gat));
  AOI21_X1  g617(.A(G120gat), .B1(new_n810), .B2(new_n650), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n650), .A2(G120gat), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n816), .B2(new_n820), .ZN(G1341gat));
  INV_X1    g620(.A(new_n816), .ZN(new_n822));
  OAI21_X1  g621(.A(G127gat), .B1(new_n822), .B2(new_n587), .ZN(new_n823));
  INV_X1    g622(.A(G127gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n810), .A2(new_n824), .A3(new_n677), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(G1342gat));
  OR3_X1    g625(.A1(new_n809), .A2(G134gat), .A3(new_n687), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n827), .A2(KEYINPUT56), .ZN(new_n828));
  OAI21_X1  g627(.A(G134gat), .B1(new_n822), .B2(new_n687), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(KEYINPUT56), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(G1343gat));
  NAND2_X1  g630(.A1(new_n666), .A2(new_n814), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n408), .B1(new_n805), .B2(new_n806), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n805), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n806), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n838), .B1(new_n805), .B2(new_n836), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n408), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n835), .B1(new_n840), .B2(new_n834), .ZN(new_n841));
  INV_X1    g640(.A(G141gat), .ZN(new_n842));
  OR3_X1    g641(.A1(new_n841), .A2(new_n842), .A3(new_n619), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n844), .A2(KEYINPUT115), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT114), .B1(new_n666), .B2(new_n418), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n453), .A2(KEYINPUT114), .A3(new_n455), .A4(new_n418), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n846), .A2(new_n384), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n618), .A3(new_n807), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n850), .A2(new_n842), .B1(KEYINPUT115), .B2(new_n844), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n843), .A2(new_n845), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n845), .B1(new_n843), .B2(new_n851), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(G1344gat));
  NAND2_X1  g653(.A1(new_n849), .A2(new_n807), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(G148gat), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n856), .A2(new_n857), .A3(new_n650), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n418), .A2(new_n834), .ZN(new_n860));
  OR3_X1    g659(.A1(new_n797), .A2(new_n804), .A3(KEYINPUT117), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT117), .B1(new_n797), .B2(new_n804), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n587), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n860), .B1(new_n863), .B2(new_n806), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n833), .A2(new_n834), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n666), .A2(new_n650), .A3(new_n814), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n867), .A2(KEYINPUT118), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n857), .B1(new_n867), .B2(KEYINPUT118), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n859), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n835), .B(new_n650), .C1(new_n840), .C2(new_n834), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n857), .A2(KEYINPUT59), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n871), .A2(KEYINPUT116), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT116), .B1(new_n871), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n858), .B1(new_n870), .B2(new_n875), .ZN(G1345gat));
  OAI21_X1  g675(.A(G155gat), .B1(new_n841), .B2(new_n587), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n677), .A2(new_n583), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n855), .B2(new_n878), .ZN(G1346gat));
  INV_X1    g678(.A(G162gat), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n841), .A2(new_n880), .A3(new_n687), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n856), .A2(new_n553), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n880), .B2(new_n882), .ZN(G1347gat));
  NAND2_X1  g682(.A1(new_n345), .A2(new_n384), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n345), .A2(new_n384), .A3(KEYINPUT120), .ZN(new_n887));
  AND4_X1   g686(.A1(new_n417), .A2(new_n886), .A3(new_n416), .A4(new_n887), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n812), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n619), .A2(new_n244), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n418), .B1(new_n287), .B2(new_n290), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n891), .A2(new_n892), .A3(new_n384), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n891), .B2(new_n384), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n411), .B1(new_n805), .B2(new_n806), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n895), .A2(new_n896), .A3(new_n618), .ZN(new_n897));
  AOI22_X1  g696(.A1(new_n889), .A2(new_n890), .B1(new_n897), .B2(new_n244), .ZN(G1348gat));
  NOR2_X1   g697(.A1(new_n718), .A2(new_n243), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n895), .A2(new_n896), .A3(new_n650), .ZN(new_n900));
  AOI22_X1  g699(.A1(new_n889), .A2(new_n899), .B1(new_n900), .B2(new_n248), .ZN(G1349gat));
  NOR2_X1   g700(.A1(new_n587), .A2(new_n225), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n895), .A2(new_n896), .A3(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n231), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n805), .A2(new_n806), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n905), .A2(new_n408), .A3(new_n677), .A4(new_n888), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n812), .A2(KEYINPUT121), .A3(new_n677), .A4(new_n888), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n903), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g709(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n906), .A2(new_n907), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n231), .A3(new_n909), .ZN(new_n916));
  INV_X1    g715(.A(new_n903), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n914), .B1(new_n918), .B2(KEYINPUT122), .ZN(new_n919));
  AOI211_X1 g718(.A(KEYINPUT122), .B(new_n903), .C1(new_n908), .C2(new_n909), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n913), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT60), .B1(new_n910), .B2(new_n923), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n924), .A2(KEYINPUT123), .A3(new_n920), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n912), .B1(new_n922), .B2(new_n925), .ZN(G1350gat));
  NOR2_X1   g725(.A1(new_n687), .A2(G190gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n895), .A2(new_n896), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n889), .A2(new_n553), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n929), .A2(new_n930), .A3(G190gat), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n929), .B2(G190gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(G1351gat));
  NAND4_X1  g732(.A1(new_n896), .A2(new_n666), .A3(new_n384), .A4(new_n418), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n934), .A2(G197gat), .A3(new_n619), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT125), .Z(new_n936));
  NAND3_X1  g735(.A1(new_n666), .A2(new_n886), .A3(new_n887), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT126), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n864), .A2(new_n865), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n939), .A3(new_n618), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT127), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G197gat), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n940), .A2(KEYINPUT127), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n936), .B1(new_n942), .B2(new_n943), .ZN(G1352gat));
  NOR3_X1   g743(.A1(new_n934), .A2(G204gat), .A3(new_n718), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT62), .ZN(new_n946));
  INV_X1    g745(.A(new_n938), .ZN(new_n947));
  INV_X1    g746(.A(new_n939), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n947), .A2(new_n948), .A3(new_n718), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n946), .B1(new_n949), .B2(new_n360), .ZN(G1353gat));
  NAND3_X1  g749(.A1(new_n938), .A2(new_n939), .A3(new_n677), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n951), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT63), .B1(new_n951), .B2(G211gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n677), .A2(new_n363), .ZN(new_n954));
  OAI22_X1  g753(.A1(new_n952), .A2(new_n953), .B1(new_n934), .B2(new_n954), .ZN(G1354gat));
  NOR3_X1   g754(.A1(new_n947), .A2(new_n948), .A3(new_n687), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n553), .A2(new_n364), .ZN(new_n957));
  OAI22_X1  g756(.A1(new_n956), .A2(new_n364), .B1(new_n934), .B2(new_n957), .ZN(G1355gat));
endmodule


