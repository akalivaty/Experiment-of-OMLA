//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n575, new_n576, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n634, new_n635, new_n638, new_n639,
    new_n641, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1215, new_n1216, new_n1217;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT66), .B(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G137), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND3_X1   g038(.A1(KEYINPUT68), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT3), .B1(KEYINPUT68), .B2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n463), .A2(new_n467), .B1(G101), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  XOR2_X1   g046(.A(KEYINPUT66), .B(G2105), .Z(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OR2_X1    g051(.A1(new_n476), .A2(KEYINPUT67), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(KEYINPUT67), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n471), .B1(new_n477), .B2(new_n478), .ZN(G160));
  NOR2_X1   g054(.A1(new_n472), .A2(new_n466), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OAI221_X1 g056(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n472), .C2(G112), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n466), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(G126), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT4), .A2(G138), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n461), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n489), .B1(new_n492), .B2(new_n467), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n472), .A2(G138), .A3(new_n473), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT69), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n493), .A2(new_n499), .A3(new_n496), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n503), .B1(KEYINPUT6), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n509), .A2(KEYINPUT70), .ZN(new_n510));
  OAI21_X1  g085(.A(G651), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT71), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(KEYINPUT70), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(G651), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n506), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G62), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n518), .A2(G50), .B1(G651), .B2(new_n524), .ZN(new_n525));
  OR2_X1    g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n528), .B1(new_n509), .B2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n529), .B1(new_n512), .B2(new_n517), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G88), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n525), .A2(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  AOI21_X1  g108(.A(new_n522), .B1(KEYINPUT6), .B2(new_n504), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n516), .B1(new_n515), .B2(G651), .ZN(new_n535));
  AOI211_X1 g110(.A(KEYINPUT71), .B(new_n504), .C1(new_n513), .C2(new_n514), .ZN(new_n536));
  OAI211_X1 g111(.A(G89), .B(new_n534), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  OAI211_X1 g112(.A(G51), .B(new_n505), .C1(new_n535), .C2(new_n536), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n528), .A2(KEYINPUT72), .A3(G63), .A4(G651), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT72), .ZN(new_n540));
  NAND2_X1  g115(.A1(G63), .A2(G651), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n522), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT7), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n543), .A2(KEYINPUT7), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n539), .A2(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n537), .A2(new_n538), .A3(new_n546), .ZN(G286));
  INV_X1    g122(.A(G286), .ZN(G168));
  OAI211_X1 g123(.A(G52), .B(new_n505), .C1(new_n535), .C2(new_n536), .ZN(new_n549));
  OAI211_X1 g124(.A(G90), .B(new_n534), .C1(new_n535), .C2(new_n536), .ZN(new_n550));
  NAND2_X1  g125(.A1(G77), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G64), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n522), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n549), .A2(new_n550), .A3(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  OAI211_X1 g131(.A(G81), .B(new_n534), .C1(new_n535), .C2(new_n536), .ZN(new_n557));
  OAI211_X1 g132(.A(G43), .B(new_n505), .C1(new_n535), .C2(new_n536), .ZN(new_n558));
  INV_X1    g133(.A(G56), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n559), .B1(new_n526), .B2(new_n527), .ZN(new_n560));
  NAND2_X1  g135(.A1(G68), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT73), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n564), .B(new_n561), .C1(new_n522), .C2(new_n559), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(G651), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n557), .A2(new_n558), .A3(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n557), .A2(new_n558), .A3(new_n566), .A4(KEYINPUT74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G860), .ZN(G153));
  NAND4_X1  g148(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g149(.A1(G1), .A2(G3), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT8), .ZN(new_n576));
  NAND4_X1  g151(.A1(G319), .A2(G483), .A3(G661), .A4(new_n576), .ZN(G188));
  NAND3_X1  g152(.A1(new_n530), .A2(KEYINPUT75), .A3(G91), .ZN(new_n578));
  OAI211_X1 g153(.A(G91), .B(new_n534), .C1(new_n535), .C2(new_n536), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(G78), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G65), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n522), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n578), .A2(new_n581), .B1(G651), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g160(.A(G53), .B(new_n505), .C1(new_n535), .C2(new_n536), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT9), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(G299));
  NAND2_X1  g163(.A1(new_n530), .A2(G87), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n518), .A2(G49), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G288));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  OAI21_X1  g168(.A(KEYINPUT76), .B1(new_n522), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G73), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(new_n503), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT76), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n528), .A2(new_n597), .A3(G61), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n518), .A2(G48), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n530), .A2(G86), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G305));
  INV_X1    g179(.A(G60), .ZN(new_n605));
  INV_X1    g180(.A(G72), .ZN(new_n606));
  OAI22_X1  g181(.A1(new_n522), .A2(new_n605), .B1(new_n606), .B2(new_n503), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI221_X1 g184(.A(KEYINPUT77), .B1(new_n606), .B2(new_n503), .C1(new_n522), .C2(new_n605), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n609), .A2(G651), .A3(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  AOI22_X1  g189(.A1(G47), .A2(new_n518), .B1(new_n530), .B2(G85), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(G290));
  NAND2_X1  g191(.A1(G301), .A2(G868), .ZN(new_n617));
  OAI211_X1 g192(.A(G92), .B(new_n534), .C1(new_n535), .C2(new_n536), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT10), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(G54), .ZN(new_n621));
  AOI211_X1 g196(.A(new_n621), .B(new_n506), .C1(new_n512), .C2(new_n517), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n528), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n623), .A2(new_n504), .ZN(new_n624));
  NOR3_X1   g199(.A1(new_n622), .A2(KEYINPUT79), .A3(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT79), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n518), .A2(G54), .ZN(new_n627));
  INV_X1    g202(.A(new_n624), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n620), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n617), .B1(new_n631), .B2(G868), .ZN(G284));
  OAI21_X1  g207(.A(new_n617), .B1(new_n631), .B2(G868), .ZN(G321));
  INV_X1    g208(.A(G868), .ZN(new_n634));
  NAND2_X1  g209(.A1(G299), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(new_n634), .B2(G168), .ZN(G297));
  OAI21_X1  g211(.A(new_n635), .B1(new_n634), .B2(G168), .ZN(G280));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n631), .B1(new_n638), .B2(G860), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT80), .ZN(G148));
  NAND2_X1  g215(.A1(new_n631), .A2(new_n638), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(G868), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n572), .B2(G868), .ZN(G323));
  XNOR2_X1  g218(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g219(.A1(new_n473), .A2(new_n469), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT12), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT13), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2100), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n480), .A2(G123), .ZN(new_n649));
  OAI221_X1 g224(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n472), .C2(G111), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n483), .A2(G135), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2096), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n648), .A2(new_n653), .ZN(G156));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT81), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2427), .B(G2430), .Z(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(KEYINPUT14), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2451), .B(G2454), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n661), .B(new_n665), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2443), .B(G2446), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(G14), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n669), .B2(new_n667), .ZN(G401));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT17), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT82), .ZN(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n675), .B2(new_n672), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n676), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n677), .B2(new_n679), .ZN(new_n681));
  INV_X1    g256(.A(new_n672), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n682), .A2(new_n678), .A3(new_n674), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT18), .Z(new_n684));
  NAND3_X1  g259(.A1(new_n673), .A2(new_n678), .A3(new_n675), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G2096), .B(G2100), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G227));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT83), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1956), .B(G2474), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT19), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT20), .Z(new_n697));
  NOR2_X1   g272(.A1(new_n690), .A2(new_n692), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n699), .A2(new_n695), .A3(new_n693), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n697), .B(new_n700), .C1(new_n695), .C2(new_n699), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1991), .B(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT84), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1981), .B(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(G229));
  NAND2_X1  g284(.A1(new_n480), .A2(G119), .ZN(new_n710));
  OAI221_X1 g285(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n472), .C2(G107), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n483), .A2(G131), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  MUX2_X1   g288(.A(G25), .B(new_n713), .S(G29), .Z(new_n714));
  XOR2_X1   g289(.A(KEYINPUT35), .B(G1991), .Z(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(G290), .A2(G16), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G24), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT85), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G1986), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n719), .A2(G23), .ZN(new_n724));
  INV_X1    g299(.A(G288), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(new_n719), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT33), .B(G1976), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n726), .A2(new_n728), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT86), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n719), .A2(G6), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n602), .A2(new_n603), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n719), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT32), .B(G1981), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n729), .A2(KEYINPUT86), .A3(new_n730), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n719), .A2(G22), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G166), .B2(new_n719), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(G1971), .Z(new_n742));
  NAND4_X1  g317(.A1(new_n733), .A2(new_n738), .A3(new_n739), .A4(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT34), .ZN(new_n745));
  AOI211_X1 g320(.A(new_n717), .B(new_n723), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT88), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n743), .A2(KEYINPUT34), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT87), .B(KEYINPUT36), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n746), .A2(new_n747), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n744), .A2(new_n745), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n723), .A2(new_n717), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n751), .A2(new_n748), .A3(new_n752), .A4(new_n749), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(KEYINPUT88), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n751), .A2(new_n748), .A3(new_n752), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(KEYINPUT36), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n750), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT25), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n483), .A2(G139), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(new_n472), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G29), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n765), .B2(G33), .ZN(new_n767));
  INV_X1    g342(.A(G2072), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n480), .A2(G129), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n483), .A2(G141), .ZN(new_n770));
  NAND3_X1  g345(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT26), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n773), .A2(new_n774), .B1(G105), .B2(new_n469), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n769), .A2(new_n770), .A3(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(new_n765), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n765), .B2(G32), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT27), .B(G1996), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n767), .A2(new_n768), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT91), .B(KEYINPUT24), .Z(new_n782));
  AOI21_X1  g357(.A(G29), .B1(new_n782), .B2(G34), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G34), .B2(new_n782), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT92), .Z(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G160), .B2(G29), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G2084), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n781), .B(new_n787), .C1(new_n768), .C2(new_n767), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT93), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n719), .A2(G19), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n572), .B2(new_n719), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT89), .B(G1341), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT30), .B(G28), .ZN(new_n794));
  OR2_X1    g369(.A1(KEYINPUT31), .A2(G11), .ZN(new_n795));
  NAND2_X1  g370(.A1(KEYINPUT31), .A2(G11), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n794), .A2(new_n765), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n652), .B2(new_n765), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n765), .A2(G26), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT28), .ZN(new_n800));
  OAI221_X1 g375(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n472), .C2(G116), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT90), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  AOI22_X1  g378(.A1(G128), .A2(new_n480), .B1(new_n483), .B2(G140), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n800), .B1(new_n806), .B2(new_n765), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n798), .B1(new_n807), .B2(G2067), .ZN(new_n808));
  INV_X1    g383(.A(G2078), .ZN(new_n809));
  NAND2_X1  g384(.A1(G164), .A2(G29), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G27), .B2(G29), .ZN(new_n811));
  OAI221_X1 g386(.A(new_n808), .B1(G2067), .B2(new_n807), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n719), .A2(G21), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G168), .B2(new_n719), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT94), .B(G1966), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G1961), .ZN(new_n817));
  NOR2_X1   g392(.A1(G5), .A2(G16), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT95), .Z(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G301), .B2(new_n719), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n765), .A2(G35), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G162), .B2(new_n765), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT29), .ZN(new_n823));
  OAI221_X1 g398(.A(new_n816), .B1(new_n817), .B2(new_n820), .C1(new_n823), .C2(G2090), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n811), .A2(new_n809), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(G2090), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OR4_X1    g402(.A1(new_n793), .A2(new_n812), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n786), .A2(G2084), .B1(new_n779), .B2(new_n780), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n817), .B2(new_n820), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT96), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n719), .A2(G20), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT23), .Z(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(G299), .B2(G16), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(G1956), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n719), .A2(G4), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n631), .B2(new_n719), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G1348), .ZN(new_n839));
  NOR4_X1   g414(.A1(new_n789), .A2(new_n828), .A3(new_n836), .A4(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n757), .A2(new_n840), .ZN(G311));
  AND3_X1   g416(.A1(new_n757), .A2(KEYINPUT97), .A3(new_n840), .ZN(new_n842));
  AOI21_X1  g417(.A(KEYINPUT97), .B1(new_n757), .B2(new_n840), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(G150));
  XNOR2_X1  g419(.A(KEYINPUT98), .B(G93), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n534), .B(new_n845), .C1(new_n535), .C2(new_n536), .ZN(new_n846));
  OAI211_X1 g421(.A(G55), .B(new_n505), .C1(new_n535), .C2(new_n536), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n848), .A2(new_n504), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G860), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT37), .Z(new_n852));
  NOR2_X1   g427(.A1(new_n850), .A2(new_n567), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n571), .B2(new_n850), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT38), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n638), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT99), .Z(new_n860));
  INV_X1    g435(.A(G860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n857), .B2(new_n858), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n852), .B1(new_n860), .B2(new_n862), .ZN(G145));
  OR2_X1    g438(.A1(new_n805), .A2(new_n497), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n805), .A2(new_n497), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n776), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n776), .B1(new_n864), .B2(new_n865), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n763), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n870), .A2(new_n764), .A3(new_n866), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n713), .B(new_n646), .ZN(new_n872));
  OR3_X1    g447(.A1(new_n472), .A2(KEYINPUT100), .A3(G118), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT100), .B1(new_n472), .B2(G118), .ZN(new_n874));
  OR2_X1    g449(.A1(G106), .A2(G2105), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n873), .A2(G2104), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  AOI22_X1  g451(.A1(G130), .A2(new_n480), .B1(new_n483), .B2(G142), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n872), .B(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n869), .A2(new_n871), .A3(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n485), .B(new_n652), .Z(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G160), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n879), .ZN(new_n885));
  INV_X1    g460(.A(new_n871), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n764), .B1(new_n870), .B2(new_n866), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(G37), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n880), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n888), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n891), .B(new_n885), .C1(new_n886), .C2(new_n887), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n890), .B1(new_n895), .B2(new_n882), .ZN(new_n896));
  AOI211_X1 g471(.A(KEYINPUT102), .B(new_n883), .C1(new_n893), .C2(new_n894), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n889), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g474(.A1(new_n850), .A2(new_n634), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n735), .A2(G290), .ZN(new_n901));
  NAND4_X1  g476(.A1(G305), .A2(new_n614), .A3(new_n613), .A4(new_n615), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(G303), .B(G288), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n901), .A3(new_n902), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(KEYINPUT103), .B2(KEYINPUT42), .ZN(new_n909));
  NAND2_X1  g484(.A1(KEYINPUT103), .A2(KEYINPUT42), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT41), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n630), .A2(G299), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT79), .B1(new_n622), .B2(new_n624), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n627), .A2(new_n626), .A3(new_n628), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI22_X1  g491(.A1(new_n916), .A2(new_n620), .B1(new_n585), .B2(new_n587), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n912), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n630), .A2(G299), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n916), .A2(new_n585), .A3(new_n587), .A4(new_n620), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n920), .A3(KEYINPUT41), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n571), .A2(new_n850), .ZN(new_n924));
  INV_X1    g499(.A(new_n853), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n641), .B(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n919), .A2(new_n920), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n928), .B1(new_n929), .B2(new_n927), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n911), .B(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n900), .B1(new_n931), .B2(new_n634), .ZN(G295));
  OAI21_X1  g507(.A(new_n900), .B1(new_n931), .B2(new_n634), .ZN(G331));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n934));
  NAND2_X1  g509(.A1(G301), .A2(KEYINPUT104), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n549), .A2(new_n550), .A3(new_n936), .A4(new_n554), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(G286), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(G168), .A2(G171), .A3(new_n936), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n854), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n939), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n943));
  INV_X1    g518(.A(new_n850), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n944), .B1(new_n569), .B2(new_n570), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n942), .B(new_n943), .C1(new_n945), .C2(new_n853), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n943), .B1(new_n926), .B2(new_n942), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n941), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n923), .ZN(new_n950));
  INV_X1    g525(.A(new_n929), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n942), .B1(new_n945), .B2(new_n853), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n941), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n908), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n942), .A2(new_n945), .A3(new_n853), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT105), .B1(new_n940), .B2(new_n854), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n955), .B1(new_n956), .B2(new_n946), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n908), .B(new_n953), .C1(new_n957), .C2(new_n922), .ZN(new_n958));
  INV_X1    g533(.A(G37), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n934), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n941), .A2(new_n952), .ZN(new_n964));
  OR2_X1    g539(.A1(new_n922), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n951), .B(new_n941), .C1(new_n947), .C2(new_n948), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n908), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT43), .B1(new_n967), .B2(new_n960), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT107), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n970), .B(KEYINPUT43), .C1(new_n967), .C2(new_n960), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n963), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT43), .B1(new_n954), .B2(new_n960), .ZN(new_n973));
  INV_X1    g548(.A(new_n908), .ZN(new_n974));
  AOI211_X1 g549(.A(new_n929), .B(new_n955), .C1(new_n956), .C2(new_n946), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n922), .A2(new_n964), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n977), .A2(new_n962), .A3(new_n959), .A4(new_n958), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT106), .B1(new_n979), .B2(new_n934), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n981));
  AOI211_X1 g556(.A(new_n981), .B(KEYINPUT44), .C1(new_n973), .C2(new_n978), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n972), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(KEYINPUT108), .B(new_n972), .C1(new_n980), .C2(new_n982), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(G397));
  AND2_X1   g562(.A1(new_n476), .A2(KEYINPUT67), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n476), .A2(KEYINPUT67), .ZN(new_n989));
  OAI211_X1 g564(.A(G40), .B(new_n470), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1384), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n497), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G8), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1976), .ZN(new_n997));
  NOR2_X1   g572(.A1(G288), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT52), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT52), .B1(G288), .B2(new_n997), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n995), .B(new_n1000), .C1(new_n997), .C2(G288), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1981), .ZN(new_n1003));
  XOR2_X1   g578(.A(KEYINPUT114), .B(G86), .Z(new_n1004));
  NAND2_X1  g579(.A1(new_n530), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1003), .B1(new_n602), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(G1981), .B2(G305), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(KEYINPUT115), .A3(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(G305), .A2(G1981), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1011), .B2(new_n1006), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n995), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1002), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(G166), .A2(new_n994), .ZN(new_n1019));
  NAND2_X1  g594(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1022), .B1(new_n1019), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1384), .B1(new_n493), .B2(new_n496), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n990), .B1(KEYINPUT45), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1384), .B1(new_n498), .B2(new_n500), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(KEYINPUT45), .B2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT110), .B(G1971), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1034), .A2(KEYINPUT111), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1028), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(G160), .A2(new_n1037), .A3(G40), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1030), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1038), .B1(new_n1039), .B2(KEYINPUT50), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT112), .B(G2090), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(new_n1034), .B2(KEYINPUT111), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1027), .B(G8), .C1(new_n1035), .C2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1034), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n990), .B1(KEYINPUT50), .B2(new_n992), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1030), .A2(new_n1036), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1046), .A2(new_n1047), .A3(new_n1041), .ZN(new_n1048));
  OAI21_X1  g623(.A(G8), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n1026), .ZN(new_n1050));
  AND3_X1   g625(.A1(G160), .A2(new_n1037), .A3(G40), .ZN(new_n1051));
  INV_X1    g626(.A(G2084), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1051), .B(new_n1052), .C1(new_n1036), .C2(new_n1030), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT45), .ZN(new_n1054));
  AOI211_X1 g629(.A(new_n1054), .B(G1384), .C1(new_n498), .C2(new_n500), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n992), .A2(new_n1054), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(G40), .A3(G160), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n815), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  AOI211_X1 g633(.A(new_n994), .B(G286), .C1(new_n1053), .C2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1018), .A2(new_n1044), .A3(new_n1050), .A4(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT63), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1059), .A2(KEYINPUT63), .ZN(new_n1065));
  OAI21_X1  g640(.A(G8), .B1(new_n1035), .B2(new_n1043), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1065), .B1(new_n1066), .B2(new_n1026), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(new_n1044), .A3(new_n1018), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT119), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1060), .A2(KEYINPUT118), .A3(new_n1061), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1067), .A2(new_n1071), .A3(new_n1044), .A4(new_n1018), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1064), .A2(new_n1069), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1011), .B(KEYINPUT116), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1016), .B1(new_n1014), .B2(new_n1010), .ZN(new_n1075));
  NOR2_X1   g650(.A1(G288), .A2(G1976), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1074), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n995), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1044), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1018), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1079), .A2(new_n1081), .A3(KEYINPUT117), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1051), .B1(new_n1036), .B2(new_n1030), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n817), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(G2078), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1030), .A2(KEYINPUT45), .ZN(new_n1094));
  OAI211_X1 g669(.A(G160), .B(G40), .C1(new_n1054), .C2(new_n992), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT53), .B1(new_n1096), .B2(new_n809), .ZN(new_n1097));
  OAI21_X1  g672(.A(G171), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1053), .A2(new_n1058), .A3(G168), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT51), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1100), .A2(new_n1101), .A3(G8), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1053), .A2(new_n1058), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(G286), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1104), .A2(G8), .A3(new_n1100), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1102), .B1(new_n1105), .B2(KEYINPUT51), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1099), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI211_X1 g683(.A(KEYINPUT62), .B(new_n1102), .C1(KEYINPUT51), .C2(new_n1105), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1040), .B2(G1961), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1087), .A2(KEYINPUT124), .A3(new_n817), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1029), .B(new_n809), .C1(KEYINPUT45), .C2(new_n1030), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT125), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n463), .A2(new_n467), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n469), .A2(G101), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(G40), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1117), .B1(new_n1120), .B2(new_n476), .ZN(new_n1121));
  INV_X1    g696(.A(new_n476), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1122), .A2(new_n470), .A3(KEYINPUT125), .A4(G40), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1028), .A2(KEYINPUT45), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1116), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1056), .A2(KEYINPUT126), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g703(.A(new_n1090), .B(G2078), .C1(new_n1028), .C2(KEYINPUT45), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1115), .A2(new_n1090), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1114), .A2(G301), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT54), .B1(new_n1131), .B2(new_n1098), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1114), .A2(new_n1130), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(G171), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1115), .A2(new_n1090), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1135), .A2(G301), .A3(new_n1088), .A4(new_n1092), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1134), .A2(KEYINPUT127), .A3(KEYINPUT54), .A4(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT127), .ZN(new_n1138));
  AOI21_X1  g713(.A(G301), .B1(new_n1114), .B2(new_n1130), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1136), .A2(KEYINPUT54), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI211_X1 g716(.A(new_n1132), .B(new_n1106), .C1(new_n1137), .C2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(KEYINPUT56), .B(G2072), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n1094), .A2(new_n1095), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(G1956), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n1148));
  NAND3_X1  g723(.A1(G299), .A2(new_n1148), .A3(KEYINPUT57), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(KEYINPUT57), .B1(G299), .B2(new_n1148), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1147), .A2(new_n1152), .ZN(new_n1153));
  OAI22_X1  g728(.A1(new_n1145), .A2(new_n1146), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(G2067), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n993), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1040), .B2(G1348), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1158), .A2(new_n631), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1153), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(KEYINPUT58), .B(G1341), .ZN(new_n1161));
  OAI22_X1  g736(.A1(new_n1031), .A2(G1996), .B1(new_n993), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT121), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1163), .A2(KEYINPUT59), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1162), .A2(new_n572), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1162), .B2(new_n572), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1153), .A2(KEYINPUT61), .A3(new_n1154), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1153), .A2(new_n1169), .A3(new_n1154), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1171), .B1(new_n1154), .B2(new_n1169), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1167), .B(new_n1168), .C1(new_n1170), .C2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g748(.A(KEYINPUT60), .B(new_n1157), .C1(new_n1040), .C2(G1348), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(KEYINPUT123), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n631), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1174), .A2(KEYINPUT123), .A3(new_n630), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n1174), .A2(KEYINPUT123), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT60), .ZN(new_n1180));
  AOI22_X1  g755(.A1(new_n1178), .A2(new_n1179), .B1(new_n1180), .B2(new_n1158), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1160), .B1(new_n1173), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1110), .B1(new_n1142), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1018), .A2(new_n1044), .A3(new_n1050), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1073), .B(new_n1086), .C1(new_n1183), .C2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1056), .A2(new_n990), .ZN(new_n1186));
  INV_X1    g761(.A(G1996), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1188), .A2(new_n776), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n805), .B(new_n1156), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1190), .B1(new_n1187), .B2(new_n777), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1186), .B(KEYINPUT109), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1189), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1192), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n713), .B(new_n715), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1193), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g771(.A(G290), .B(G1986), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1196), .B1(new_n1186), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1185), .A2(new_n1198), .ZN(new_n1199));
  XOR2_X1   g774(.A(new_n1188), .B(KEYINPUT46), .Z(new_n1200));
  NAND2_X1  g775(.A1(new_n1190), .A2(new_n777), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1200), .B1(new_n1192), .B2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT47), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n713), .A2(new_n716), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1193), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n806), .A2(new_n1156), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1194), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g782(.A1(G290), .A2(G1986), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1208), .A2(new_n1186), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1209), .B(KEYINPUT48), .Z(new_n1210));
  NOR2_X1   g785(.A1(new_n1196), .A2(new_n1210), .ZN(new_n1211));
  NOR3_X1   g786(.A1(new_n1203), .A2(new_n1207), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1199), .A2(new_n1212), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g788(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1215));
  NAND3_X1  g789(.A1(new_n898), .A2(new_n708), .A3(new_n1215), .ZN(new_n1216));
  INV_X1    g790(.A(new_n979), .ZN(new_n1217));
  NOR2_X1   g791(.A1(new_n1216), .A2(new_n1217), .ZN(G308));
  OR2_X1    g792(.A1(new_n1216), .A2(new_n1217), .ZN(G225));
endmodule


