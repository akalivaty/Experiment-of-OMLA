

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U555 ( .A1(n698), .A2(n809), .ZN(n739) );
  NOR2_X1 U556 ( .A1(G164), .A2(G1384), .ZN(n809) );
  OR2_X1 U557 ( .A1(n941), .A2(n714), .ZN(n715) );
  NOR2_X1 U558 ( .A1(n732), .A2(G168), .ZN(n733) );
  XNOR2_X1 U559 ( .A(KEYINPUT97), .B(KEYINPUT29), .ZN(n722) );
  XNOR2_X1 U560 ( .A(n723), .B(n722), .ZN(n728) );
  AND2_X1 U561 ( .A1(n831), .A2(n830), .ZN(n832) );
  NOR2_X1 U562 ( .A1(G543), .A2(G651), .ZN(n660) );
  NOR2_X1 U563 ( .A1(G651), .A2(n630), .ZN(n653) );
  OR2_X1 U564 ( .A1(n833), .A2(n832), .ZN(n834) );
  INV_X1 U565 ( .A(KEYINPUT89), .ZN(n530) );
  NOR2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  XOR2_X1 U567 ( .A(KEYINPUT17), .B(n521), .Z(n894) );
  NAND2_X1 U568 ( .A1(G138), .A2(n894), .ZN(n524) );
  XNOR2_X1 U569 ( .A(G2104), .B(KEYINPUT64), .ZN(n526) );
  INV_X1 U570 ( .A(G2105), .ZN(n525) );
  AND2_X1 U571 ( .A1(n526), .A2(n525), .ZN(n522) );
  XOR2_X2 U572 ( .A(KEYINPUT65), .B(n522), .Z(n895) );
  NAND2_X1 U573 ( .A1(G102), .A2(n895), .ZN(n523) );
  NAND2_X1 U574 ( .A1(n524), .A2(n523), .ZN(n533) );
  NOR2_X1 U575 ( .A1(n526), .A2(n525), .ZN(n891) );
  NAND2_X1 U576 ( .A1(n891), .A2(G126), .ZN(n529) );
  NAND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  XOR2_X2 U578 ( .A(KEYINPUT66), .B(n527), .Z(n892) );
  NAND2_X1 U579 ( .A1(G114), .A2(n892), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n531) );
  XNOR2_X1 U581 ( .A(n531), .B(n530), .ZN(n532) );
  NOR2_X1 U582 ( .A1(n533), .A2(n532), .ZN(G164) );
  XOR2_X1 U583 ( .A(G543), .B(KEYINPUT0), .Z(n630) );
  NAND2_X1 U584 ( .A1(G51), .A2(n653), .ZN(n537) );
  INV_X1 U585 ( .A(G651), .ZN(n540) );
  NOR2_X1 U586 ( .A1(G543), .A2(n540), .ZN(n535) );
  XNOR2_X1 U587 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n534) );
  XNOR2_X1 U588 ( .A(n535), .B(n534), .ZN(n655) );
  NAND2_X1 U589 ( .A1(G63), .A2(n655), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U591 ( .A(KEYINPUT6), .B(n538), .ZN(n546) );
  NAND2_X1 U592 ( .A1(n660), .A2(G89), .ZN(n539) );
  XNOR2_X1 U593 ( .A(KEYINPUT4), .B(n539), .ZN(n543) );
  NOR2_X1 U594 ( .A1(n630), .A2(n540), .ZN(n661) );
  NAND2_X1 U595 ( .A1(n661), .A2(G76), .ZN(n541) );
  XOR2_X1 U596 ( .A(KEYINPUT73), .B(n541), .Z(n542) );
  NAND2_X1 U597 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U598 ( .A(n544), .B(KEYINPUT5), .Z(n545) );
  NOR2_X1 U599 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U600 ( .A(KEYINPUT7), .B(n547), .Z(n548) );
  XNOR2_X1 U601 ( .A(KEYINPUT74), .B(n548), .ZN(G168) );
  XOR2_X1 U602 ( .A(G2443), .B(G2446), .Z(n550) );
  XNOR2_X1 U603 ( .A(G2427), .B(G2451), .ZN(n549) );
  XNOR2_X1 U604 ( .A(n550), .B(n549), .ZN(n556) );
  XOR2_X1 U605 ( .A(G2430), .B(G2454), .Z(n552) );
  XNOR2_X1 U606 ( .A(G1348), .B(G1341), .ZN(n551) );
  XNOR2_X1 U607 ( .A(n552), .B(n551), .ZN(n554) );
  XOR2_X1 U608 ( .A(G2435), .B(G2438), .Z(n553) );
  XNOR2_X1 U609 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U610 ( .A(n556), .B(n555), .Z(n557) );
  AND2_X1 U611 ( .A1(G14), .A2(n557), .ZN(G401) );
  NAND2_X1 U612 ( .A1(G52), .A2(n653), .ZN(n559) );
  NAND2_X1 U613 ( .A1(G64), .A2(n655), .ZN(n558) );
  NAND2_X1 U614 ( .A1(n559), .A2(n558), .ZN(n565) );
  NAND2_X1 U615 ( .A1(n660), .A2(G90), .ZN(n560) );
  XOR2_X1 U616 ( .A(KEYINPUT71), .B(n560), .Z(n562) );
  NAND2_X1 U617 ( .A1(n661), .A2(G77), .ZN(n561) );
  NAND2_X1 U618 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U619 ( .A(KEYINPUT9), .B(n563), .Z(n564) );
  NOR2_X1 U620 ( .A1(n565), .A2(n564), .ZN(G171) );
  AND2_X1 U621 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U622 ( .A1(G111), .A2(n892), .ZN(n572) );
  NAND2_X1 U623 ( .A1(G135), .A2(n894), .ZN(n567) );
  NAND2_X1 U624 ( .A1(G99), .A2(n895), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n567), .A2(n566), .ZN(n570) );
  NAND2_X1 U626 ( .A1(n891), .A2(G123), .ZN(n568) );
  XOR2_X1 U627 ( .A(KEYINPUT18), .B(n568), .Z(n569) );
  NOR2_X1 U628 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U629 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U630 ( .A(KEYINPUT79), .B(n573), .Z(n1008) );
  XNOR2_X1 U631 ( .A(G2096), .B(n1008), .ZN(n574) );
  OR2_X1 U632 ( .A1(G2100), .A2(n574), .ZN(G156) );
  INV_X1 U633 ( .A(G860), .ZN(n611) );
  NAND2_X1 U634 ( .A1(n660), .A2(G81), .ZN(n575) );
  XNOR2_X1 U635 ( .A(n575), .B(KEYINPUT12), .ZN(n577) );
  NAND2_X1 U636 ( .A1(G68), .A2(n661), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U638 ( .A(n578), .B(KEYINPUT13), .ZN(n580) );
  NAND2_X1 U639 ( .A1(G43), .A2(n653), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U641 ( .A1(n655), .A2(G56), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT14), .B(n581), .Z(n582) );
  NOR2_X1 U643 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U644 ( .A(KEYINPUT72), .B(n584), .Z(n962) );
  OR2_X1 U645 ( .A1(n611), .A2(n962), .ZN(G153) );
  INV_X1 U646 ( .A(G120), .ZN(G236) );
  INV_X1 U647 ( .A(G69), .ZN(G235) );
  INV_X1 U648 ( .A(G108), .ZN(G238) );
  NAND2_X1 U649 ( .A1(G137), .A2(n894), .ZN(n586) );
  NAND2_X1 U650 ( .A1(G113), .A2(n892), .ZN(n585) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n694) );
  NAND2_X1 U652 ( .A1(n895), .A2(G101), .ZN(n587) );
  XOR2_X1 U653 ( .A(KEYINPUT23), .B(n587), .Z(n589) );
  NAND2_X1 U654 ( .A1(n891), .A2(G125), .ZN(n588) );
  AND2_X1 U655 ( .A1(n589), .A2(n588), .ZN(n697) );
  INV_X1 U656 ( .A(n697), .ZN(n590) );
  NOR2_X1 U657 ( .A1(n694), .A2(n590), .ZN(G160) );
  XOR2_X1 U658 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U659 ( .A1(G7), .A2(G661), .ZN(n591) );
  XNOR2_X1 U660 ( .A(n591), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U661 ( .A(G223), .ZN(n838) );
  NAND2_X1 U662 ( .A1(n838), .A2(G567), .ZN(n592) );
  XOR2_X1 U663 ( .A(KEYINPUT11), .B(n592), .Z(G234) );
  INV_X1 U664 ( .A(G171), .ZN(G301) );
  NAND2_X1 U665 ( .A1(G868), .A2(G301), .ZN(n601) );
  NAND2_X1 U666 ( .A1(G92), .A2(n660), .ZN(n594) );
  NAND2_X1 U667 ( .A1(G79), .A2(n661), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U669 ( .A1(G54), .A2(n653), .ZN(n596) );
  NAND2_X1 U670 ( .A1(G66), .A2(n655), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U672 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U673 ( .A(KEYINPUT15), .B(n599), .Z(n941) );
  INV_X1 U674 ( .A(n941), .ZN(n615) );
  INV_X1 U675 ( .A(G868), .ZN(n673) );
  NAND2_X1 U676 ( .A1(n615), .A2(n673), .ZN(n600) );
  NAND2_X1 U677 ( .A1(n601), .A2(n600), .ZN(G284) );
  NAND2_X1 U678 ( .A1(G53), .A2(n653), .ZN(n603) );
  NAND2_X1 U679 ( .A1(G65), .A2(n655), .ZN(n602) );
  NAND2_X1 U680 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U681 ( .A1(G91), .A2(n660), .ZN(n605) );
  NAND2_X1 U682 ( .A1(G78), .A2(n661), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n1029) );
  NAND2_X1 U685 ( .A1(n1029), .A2(n673), .ZN(n608) );
  XNOR2_X1 U686 ( .A(n608), .B(KEYINPUT75), .ZN(n610) );
  NOR2_X1 U687 ( .A1(G286), .A2(n673), .ZN(n609) );
  NOR2_X1 U688 ( .A1(n610), .A2(n609), .ZN(G297) );
  NAND2_X1 U689 ( .A1(n611), .A2(G559), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n612), .A2(n941), .ZN(n613) );
  XNOR2_X1 U691 ( .A(n613), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U692 ( .A1(n962), .A2(G868), .ZN(n614) );
  XNOR2_X1 U693 ( .A(KEYINPUT76), .B(n614), .ZN(n620) );
  NOR2_X1 U694 ( .A1(n615), .A2(n673), .ZN(n616) );
  XNOR2_X1 U695 ( .A(n616), .B(KEYINPUT77), .ZN(n617) );
  NOR2_X1 U696 ( .A1(G559), .A2(n617), .ZN(n618) );
  XNOR2_X1 U697 ( .A(KEYINPUT78), .B(n618), .ZN(n619) );
  NOR2_X1 U698 ( .A1(n620), .A2(n619), .ZN(G282) );
  NAND2_X1 U699 ( .A1(G55), .A2(n653), .ZN(n622) );
  NAND2_X1 U700 ( .A1(G67), .A2(n655), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n660), .A2(G93), .ZN(n623) );
  XOR2_X1 U703 ( .A(KEYINPUT80), .B(n623), .Z(n624) );
  NOR2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n661), .A2(G80), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n674) );
  NAND2_X1 U707 ( .A1(G559), .A2(n941), .ZN(n628) );
  XNOR2_X1 U708 ( .A(n628), .B(n962), .ZN(n671) );
  NOR2_X1 U709 ( .A1(n671), .A2(G860), .ZN(n629) );
  XOR2_X1 U710 ( .A(n674), .B(n629), .Z(G145) );
  NAND2_X1 U711 ( .A1(G87), .A2(n630), .ZN(n632) );
  NAND2_X1 U712 ( .A1(G74), .A2(G651), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U714 ( .A1(n655), .A2(n633), .ZN(n636) );
  NAND2_X1 U715 ( .A1(G49), .A2(n653), .ZN(n634) );
  XOR2_X1 U716 ( .A(KEYINPUT81), .B(n634), .Z(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U718 ( .A1(G50), .A2(n653), .ZN(n638) );
  NAND2_X1 U719 ( .A1(G62), .A2(n655), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U721 ( .A(KEYINPUT84), .B(n639), .Z(n643) );
  NAND2_X1 U722 ( .A1(G88), .A2(n660), .ZN(n641) );
  NAND2_X1 U723 ( .A1(G75), .A2(n661), .ZN(n640) );
  AND2_X1 U724 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U725 ( .A1(n643), .A2(n642), .ZN(G303) );
  INV_X1 U726 ( .A(G303), .ZN(G166) );
  NAND2_X1 U727 ( .A1(G73), .A2(n661), .ZN(n644) );
  XNOR2_X1 U728 ( .A(n644), .B(KEYINPUT82), .ZN(n645) );
  XNOR2_X1 U729 ( .A(n645), .B(KEYINPUT2), .ZN(n647) );
  NAND2_X1 U730 ( .A1(G86), .A2(n660), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U732 ( .A1(G48), .A2(n653), .ZN(n649) );
  NAND2_X1 U733 ( .A1(G61), .A2(n655), .ZN(n648) );
  NAND2_X1 U734 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U735 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U736 ( .A(KEYINPUT83), .B(n652), .ZN(G305) );
  NAND2_X1 U737 ( .A1(n653), .A2(G47), .ZN(n654) );
  XNOR2_X1 U738 ( .A(KEYINPUT69), .B(n654), .ZN(n658) );
  NAND2_X1 U739 ( .A1(n655), .A2(G60), .ZN(n656) );
  XOR2_X1 U740 ( .A(KEYINPUT68), .B(n656), .Z(n657) );
  NOR2_X1 U741 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U742 ( .A(KEYINPUT70), .B(n659), .ZN(n665) );
  NAND2_X1 U743 ( .A1(G85), .A2(n660), .ZN(n663) );
  NAND2_X1 U744 ( .A1(G72), .A2(n661), .ZN(n662) );
  AND2_X1 U745 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U746 ( .A1(n665), .A2(n664), .ZN(G290) );
  XNOR2_X1 U747 ( .A(KEYINPUT19), .B(G288), .ZN(n666) );
  XNOR2_X1 U748 ( .A(n666), .B(n674), .ZN(n667) );
  XNOR2_X1 U749 ( .A(n1029), .B(n667), .ZN(n670) );
  XNOR2_X1 U750 ( .A(G166), .B(G305), .ZN(n668) );
  XNOR2_X1 U751 ( .A(n668), .B(G290), .ZN(n669) );
  XNOR2_X1 U752 ( .A(n670), .B(n669), .ZN(n909) );
  XOR2_X1 U753 ( .A(n909), .B(n671), .Z(n672) );
  NOR2_X1 U754 ( .A1(n673), .A2(n672), .ZN(n676) );
  NOR2_X1 U755 ( .A1(G868), .A2(n674), .ZN(n675) );
  NOR2_X1 U756 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U757 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U758 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U759 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U761 ( .A1(n680), .A2(G2072), .ZN(n681) );
  XOR2_X1 U762 ( .A(KEYINPUT85), .B(n681), .Z(G158) );
  XNOR2_X1 U763 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U764 ( .A1(G132), .A2(G82), .ZN(n682) );
  XNOR2_X1 U765 ( .A(n682), .B(KEYINPUT86), .ZN(n683) );
  XNOR2_X1 U766 ( .A(n683), .B(KEYINPUT22), .ZN(n684) );
  NOR2_X1 U767 ( .A1(G218), .A2(n684), .ZN(n685) );
  NAND2_X1 U768 ( .A1(G96), .A2(n685), .ZN(n843) );
  NAND2_X1 U769 ( .A1(n843), .A2(G2106), .ZN(n691) );
  NOR2_X1 U770 ( .A1(G235), .A2(G236), .ZN(n686) );
  XNOR2_X1 U771 ( .A(n686), .B(KEYINPUT87), .ZN(n687) );
  NOR2_X1 U772 ( .A1(G238), .A2(n687), .ZN(n688) );
  NAND2_X1 U773 ( .A1(G57), .A2(n688), .ZN(n842) );
  NAND2_X1 U774 ( .A1(G567), .A2(n842), .ZN(n689) );
  XNOR2_X1 U775 ( .A(KEYINPUT88), .B(n689), .ZN(n690) );
  NAND2_X1 U776 ( .A1(n691), .A2(n690), .ZN(n921) );
  NAND2_X1 U777 ( .A1(G483), .A2(G661), .ZN(n692) );
  NOR2_X1 U778 ( .A1(n921), .A2(n692), .ZN(n841) );
  NAND2_X1 U779 ( .A1(n841), .A2(G36), .ZN(G176) );
  NOR2_X1 U780 ( .A1(G1971), .A2(G303), .ZN(n693) );
  NOR2_X1 U781 ( .A1(G1976), .A2(G288), .ZN(n952) );
  NOR2_X1 U782 ( .A1(n693), .A2(n952), .ZN(n761) );
  XNOR2_X1 U783 ( .A(KEYINPUT101), .B(KEYINPUT32), .ZN(n750) );
  INV_X1 U784 ( .A(G40), .ZN(n695) );
  NOR2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U786 ( .A1(n697), .A2(n696), .ZN(n808) );
  INV_X1 U787 ( .A(n808), .ZN(n698) );
  NAND2_X1 U788 ( .A1(n739), .A2(G1956), .ZN(n701) );
  INV_X1 U789 ( .A(n739), .ZN(n704) );
  NAND2_X1 U790 ( .A1(n704), .A2(G2072), .ZN(n699) );
  XOR2_X1 U791 ( .A(KEYINPUT27), .B(n699), .Z(n700) );
  NAND2_X1 U792 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U793 ( .A(n702), .B(KEYINPUT95), .ZN(n717) );
  OR2_X1 U794 ( .A1(n1029), .A2(n717), .ZN(n703) );
  XNOR2_X1 U795 ( .A(n703), .B(KEYINPUT28), .ZN(n721) );
  NAND2_X1 U796 ( .A1(n704), .A2(G1996), .ZN(n705) );
  XNOR2_X1 U797 ( .A(n705), .B(KEYINPUT26), .ZN(n707) );
  NAND2_X1 U798 ( .A1(G1341), .A2(n739), .ZN(n706) );
  NAND2_X1 U799 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U800 ( .A(n708), .B(KEYINPUT96), .ZN(n709) );
  NOR2_X1 U801 ( .A1(n709), .A2(n962), .ZN(n714) );
  NAND2_X1 U802 ( .A1(n714), .A2(n941), .ZN(n713) );
  NOR2_X1 U803 ( .A1(G2067), .A2(n739), .ZN(n711) );
  NOR2_X1 U804 ( .A1(n704), .A2(G1348), .ZN(n710) );
  NOR2_X1 U805 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n716) );
  NAND2_X1 U807 ( .A1(n716), .A2(n715), .ZN(n719) );
  NAND2_X1 U808 ( .A1(n1029), .A2(n717), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U810 ( .A1(n721), .A2(n720), .ZN(n723) );
  NOR2_X1 U811 ( .A1(n704), .A2(G1961), .ZN(n724) );
  XOR2_X1 U812 ( .A(KEYINPUT94), .B(n724), .Z(n726) );
  XNOR2_X1 U813 ( .A(KEYINPUT25), .B(G2078), .ZN(n929) );
  NAND2_X1 U814 ( .A1(n704), .A2(n929), .ZN(n725) );
  NAND2_X1 U815 ( .A1(n726), .A2(n725), .ZN(n734) );
  NAND2_X1 U816 ( .A1(G171), .A2(n734), .ZN(n727) );
  NAND2_X1 U817 ( .A1(n728), .A2(n727), .ZN(n751) );
  NAND2_X1 U818 ( .A1(G8), .A2(n739), .ZN(n822) );
  NOR2_X1 U819 ( .A1(G1966), .A2(n822), .ZN(n757) );
  NOR2_X1 U820 ( .A1(G2084), .A2(n739), .ZN(n753) );
  NOR2_X1 U821 ( .A1(n757), .A2(n753), .ZN(n729) );
  XNOR2_X1 U822 ( .A(n729), .B(KEYINPUT98), .ZN(n730) );
  NAND2_X1 U823 ( .A1(n730), .A2(G8), .ZN(n731) );
  XNOR2_X1 U824 ( .A(KEYINPUT30), .B(n731), .ZN(n732) );
  XNOR2_X1 U825 ( .A(n733), .B(KEYINPUT99), .ZN(n737) );
  NOR2_X1 U826 ( .A1(G171), .A2(n734), .ZN(n735) );
  XOR2_X1 U827 ( .A(KEYINPUT100), .B(n735), .Z(n736) );
  NAND2_X1 U828 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U829 ( .A(n738), .B(KEYINPUT31), .ZN(n752) );
  NOR2_X1 U830 ( .A1(G1971), .A2(n822), .ZN(n741) );
  NOR2_X1 U831 ( .A1(G2090), .A2(n739), .ZN(n740) );
  NOR2_X1 U832 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U833 ( .A1(n742), .A2(G303), .ZN(n744) );
  AND2_X1 U834 ( .A1(n752), .A2(n744), .ZN(n743) );
  NAND2_X1 U835 ( .A1(n751), .A2(n743), .ZN(n747) );
  INV_X1 U836 ( .A(n744), .ZN(n745) );
  OR2_X1 U837 ( .A1(n745), .A2(G286), .ZN(n746) );
  AND2_X1 U838 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U839 ( .A1(n748), .A2(G8), .ZN(n749) );
  XNOR2_X1 U840 ( .A(n750), .B(n749), .ZN(n759) );
  NAND2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n755) );
  NAND2_X1 U842 ( .A1(G8), .A2(n753), .ZN(n754) );
  NAND2_X1 U843 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U844 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X2 U845 ( .A1(n759), .A2(n758), .ZN(n825) );
  INV_X1 U846 ( .A(n825), .ZN(n760) );
  NAND2_X1 U847 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n949) );
  NAND2_X1 U849 ( .A1(n762), .A2(n949), .ZN(n764) );
  INV_X1 U850 ( .A(n822), .ZN(n827) );
  NAND2_X1 U851 ( .A1(n827), .A2(KEYINPUT102), .ZN(n763) );
  NOR2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U853 ( .A1(KEYINPUT33), .A2(n765), .ZN(n772) );
  INV_X1 U854 ( .A(KEYINPUT102), .ZN(n766) );
  NAND2_X1 U855 ( .A1(n766), .A2(n952), .ZN(n769) );
  NAND2_X1 U856 ( .A1(n952), .A2(KEYINPUT33), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n767), .A2(KEYINPUT102), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U859 ( .A1(n822), .A2(n770), .ZN(n771) );
  NOR2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n818) );
  XOR2_X1 U861 ( .A(G1981), .B(G305), .Z(n946) );
  XOR2_X1 U862 ( .A(KEYINPUT92), .B(KEYINPUT38), .Z(n774) );
  NAND2_X1 U863 ( .A1(G105), .A2(n895), .ZN(n773) );
  XNOR2_X1 U864 ( .A(n774), .B(n773), .ZN(n778) );
  NAND2_X1 U865 ( .A1(G141), .A2(n894), .ZN(n776) );
  NAND2_X1 U866 ( .A1(G117), .A2(n892), .ZN(n775) );
  NAND2_X1 U867 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n891), .A2(G129), .ZN(n779) );
  NAND2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n873) );
  NOR2_X1 U871 ( .A1(G1996), .A2(n873), .ZN(n1018) );
  NAND2_X1 U872 ( .A1(G1996), .A2(n873), .ZN(n781) );
  XOR2_X1 U873 ( .A(KEYINPUT93), .B(n781), .Z(n790) );
  NAND2_X1 U874 ( .A1(n891), .A2(G119), .ZN(n783) );
  NAND2_X1 U875 ( .A1(G107), .A2(n892), .ZN(n782) );
  NAND2_X1 U876 ( .A1(n783), .A2(n782), .ZN(n787) );
  NAND2_X1 U877 ( .A1(G131), .A2(n894), .ZN(n785) );
  NAND2_X1 U878 ( .A1(G95), .A2(n895), .ZN(n784) );
  NAND2_X1 U879 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U880 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U881 ( .A(n788), .B(KEYINPUT91), .ZN(n872) );
  NAND2_X1 U882 ( .A1(G1991), .A2(n872), .ZN(n789) );
  NAND2_X1 U883 ( .A1(n790), .A2(n789), .ZN(n1005) );
  NOR2_X1 U884 ( .A1(G1986), .A2(G290), .ZN(n791) );
  NOR2_X1 U885 ( .A1(G1991), .A2(n872), .ZN(n1010) );
  NOR2_X1 U886 ( .A1(n791), .A2(n1010), .ZN(n792) );
  NOR2_X1 U887 ( .A1(n1005), .A2(n792), .ZN(n793) );
  NOR2_X1 U888 ( .A1(n1018), .A2(n793), .ZN(n794) );
  XNOR2_X1 U889 ( .A(KEYINPUT39), .B(n794), .ZN(n805) );
  XNOR2_X1 U890 ( .A(G2067), .B(KEYINPUT37), .ZN(n806) );
  XNOR2_X1 U891 ( .A(KEYINPUT90), .B(KEYINPUT34), .ZN(n798) );
  NAND2_X1 U892 ( .A1(G140), .A2(n894), .ZN(n796) );
  NAND2_X1 U893 ( .A1(G104), .A2(n895), .ZN(n795) );
  NAND2_X1 U894 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U895 ( .A(n798), .B(n797), .ZN(n803) );
  NAND2_X1 U896 ( .A1(n891), .A2(G128), .ZN(n800) );
  NAND2_X1 U897 ( .A1(G116), .A2(n892), .ZN(n799) );
  NAND2_X1 U898 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U899 ( .A(KEYINPUT35), .B(n801), .Z(n802) );
  NOR2_X1 U900 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U901 ( .A(KEYINPUT36), .B(n804), .ZN(n889) );
  NOR2_X1 U902 ( .A1(n806), .A2(n889), .ZN(n811) );
  INV_X1 U903 ( .A(n811), .ZN(n1007) );
  NAND2_X1 U904 ( .A1(n805), .A2(n1007), .ZN(n807) );
  NAND2_X1 U905 ( .A1(n806), .A2(n889), .ZN(n1006) );
  NAND2_X1 U906 ( .A1(n807), .A2(n1006), .ZN(n810) );
  NOR2_X1 U907 ( .A1(n809), .A2(n808), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n810), .A2(n813), .ZN(n830) );
  INV_X1 U909 ( .A(n830), .ZN(n816) );
  XOR2_X1 U910 ( .A(G1986), .B(G290), .Z(n957) );
  NOR2_X1 U911 ( .A1(n811), .A2(n1005), .ZN(n812) );
  NAND2_X1 U912 ( .A1(n957), .A2(n812), .ZN(n814) );
  NAND2_X1 U913 ( .A1(n814), .A2(n813), .ZN(n815) );
  OR2_X1 U914 ( .A1(n816), .A2(n815), .ZN(n819) );
  AND2_X1 U915 ( .A1(n946), .A2(n819), .ZN(n817) );
  NAND2_X1 U916 ( .A1(n818), .A2(n817), .ZN(n835) );
  INV_X1 U917 ( .A(n819), .ZN(n833) );
  NOR2_X1 U918 ( .A1(G1981), .A2(G305), .ZN(n820) );
  XOR2_X1 U919 ( .A(n820), .B(KEYINPUT24), .Z(n821) );
  NOR2_X1 U920 ( .A1(n822), .A2(n821), .ZN(n829) );
  NAND2_X1 U921 ( .A1(G166), .A2(G8), .ZN(n823) );
  NOR2_X1 U922 ( .A1(G2090), .A2(n823), .ZN(n824) );
  NOR2_X1 U923 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U924 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U925 ( .A1(n829), .A2(n828), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n835), .A2(n834), .ZN(n837) );
  XOR2_X1 U927 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n836) );
  XNOR2_X1 U928 ( .A(n837), .B(n836), .ZN(G329) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n838), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n839) );
  NAND2_X1 U931 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U933 ( .A1(n841), .A2(n840), .ZN(G188) );
  XOR2_X1 U934 ( .A(G96), .B(KEYINPUT104), .Z(G221) );
  INV_X1 U936 ( .A(G132), .ZN(G219) );
  INV_X1 U937 ( .A(G82), .ZN(G220) );
  NOR2_X1 U938 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  XOR2_X1 U940 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n845) );
  XNOR2_X1 U941 ( .A(G2678), .B(KEYINPUT105), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U943 ( .A(KEYINPUT43), .B(G2090), .Z(n847) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2072), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U946 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U947 ( .A(G2096), .B(G2100), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n853) );
  XOR2_X1 U949 ( .A(G2078), .B(G2084), .Z(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(G227) );
  XOR2_X1 U951 ( .A(G1991), .B(G1976), .Z(n855) );
  XNOR2_X1 U952 ( .A(G1956), .B(G1971), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U954 ( .A(G1986), .B(G1981), .Z(n857) );
  XNOR2_X1 U955 ( .A(G1966), .B(G1961), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U957 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U958 ( .A(KEYINPUT41), .B(G2474), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(n863) );
  XOR2_X1 U960 ( .A(G1996), .B(KEYINPUT107), .Z(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(G229) );
  NAND2_X1 U962 ( .A1(n895), .A2(G100), .ZN(n865) );
  NAND2_X1 U963 ( .A1(G112), .A2(n892), .ZN(n864) );
  NAND2_X1 U964 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U965 ( .A(KEYINPUT108), .B(n866), .ZN(n871) );
  NAND2_X1 U966 ( .A1(G124), .A2(n891), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n867), .B(KEYINPUT44), .ZN(n869) );
  NAND2_X1 U968 ( .A1(n894), .A2(G136), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U970 ( .A1(n871), .A2(n870), .ZN(G162) );
  XNOR2_X1 U971 ( .A(G164), .B(n872), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n874), .B(n873), .ZN(n886) );
  XOR2_X1 U973 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n884) );
  NAND2_X1 U974 ( .A1(n891), .A2(G127), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G115), .A2(n892), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n877), .B(KEYINPUT47), .ZN(n879) );
  NAND2_X1 U978 ( .A1(G103), .A2(n895), .ZN(n878) );
  NAND2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G139), .A2(n894), .ZN(n880) );
  XNOR2_X1 U981 ( .A(KEYINPUT111), .B(n880), .ZN(n881) );
  NOR2_X1 U982 ( .A1(n882), .A2(n881), .ZN(n1000) );
  XNOR2_X1 U983 ( .A(n1000), .B(KEYINPUT112), .ZN(n883) );
  XNOR2_X1 U984 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U985 ( .A(n886), .B(n885), .Z(n888) );
  XNOR2_X1 U986 ( .A(G160), .B(G162), .ZN(n887) );
  XNOR2_X1 U987 ( .A(n888), .B(n887), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n906) );
  NAND2_X1 U989 ( .A1(G130), .A2(n891), .ZN(n903) );
  NAND2_X1 U990 ( .A1(G118), .A2(n892), .ZN(n893) );
  XNOR2_X1 U991 ( .A(KEYINPUT109), .B(n893), .ZN(n901) );
  NAND2_X1 U992 ( .A1(G142), .A2(n894), .ZN(n897) );
  NAND2_X1 U993 ( .A1(G106), .A2(n895), .ZN(n896) );
  NAND2_X1 U994 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U995 ( .A(KEYINPUT110), .B(n898), .Z(n899) );
  XNOR2_X1 U996 ( .A(KEYINPUT45), .B(n899), .ZN(n900) );
  NOR2_X1 U997 ( .A1(n901), .A2(n900), .ZN(n902) );
  NAND2_X1 U998 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n904), .B(n1008), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n907), .ZN(n908) );
  XOR2_X1 U1002 ( .A(KEYINPUT113), .B(n908), .Z(G395) );
  XNOR2_X1 U1003 ( .A(G286), .B(n909), .ZN(n911) );
  XNOR2_X1 U1004 ( .A(n941), .B(G171), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(n912), .B(n962), .ZN(n913) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n913), .ZN(G397) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(n914), .B(KEYINPUT49), .ZN(n917) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n915), .B(KEYINPUT115), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(n920) );
  NOR2_X1 U1013 ( .A1(G401), .A2(n921), .ZN(n918) );
  XNOR2_X1 U1014 ( .A(n918), .B(KEYINPUT114), .ZN(n919) );
  NAND2_X1 U1015 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(n921), .ZN(G319) );
  INV_X1 U1018 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1019 ( .A(G2067), .B(G26), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(G33), .B(G2072), .ZN(n922) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n928) );
  XOR2_X1 U1022 ( .A(G1991), .B(G25), .Z(n924) );
  NAND2_X1 U1023 ( .A1(n924), .A2(G28), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(G32), .B(G1996), .ZN(n925) );
  NOR2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n931) );
  XOR2_X1 U1027 ( .A(G27), .B(n929), .Z(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1029 ( .A(KEYINPUT53), .B(n932), .Z(n936) );
  XNOR2_X1 U1030 ( .A(KEYINPUT54), .B(KEYINPUT117), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(n933), .B(G34), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(G2084), .B(n934), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(G35), .B(G2090), .ZN(n937) );
  NOR2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1036 ( .A(KEYINPUT55), .B(n939), .Z(n940) );
  NOR2_X1 U1037 ( .A1(G29), .A2(n940), .ZN(n998) );
  XNOR2_X1 U1038 ( .A(G16), .B(KEYINPUT56), .ZN(n968) );
  XNOR2_X1 U1039 ( .A(G1348), .B(n941), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(G171), .B(G1961), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(n942), .B(KEYINPUT118), .ZN(n943) );
  NAND2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(n945), .B(KEYINPUT119), .ZN(n966) );
  XNOR2_X1 U1044 ( .A(G1966), .B(G168), .ZN(n947) );
  NAND2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(KEYINPUT57), .B(n948), .ZN(n961) );
  XNOR2_X1 U1047 ( .A(n1029), .B(G1956), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(G166), .B(G1971), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(n953), .B(KEYINPUT120), .ZN(n954) );
  NAND2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1053 ( .A(KEYINPUT121), .B(n956), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1055 ( .A(KEYINPUT122), .B(n959), .Z(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(G1341), .B(n962), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n994) );
  INV_X1 U1061 ( .A(G16), .ZN(n992) );
  XOR2_X1 U1062 ( .A(G1976), .B(G23), .Z(n970) );
  XOR2_X1 U1063 ( .A(G1971), .B(G22), .Z(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(G24), .B(G1986), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1067 ( .A(KEYINPUT58), .B(n973), .Z(n989) );
  XOR2_X1 U1068 ( .A(G1961), .B(G5), .Z(n983) );
  XNOR2_X1 U1069 ( .A(G1348), .B(KEYINPUT59), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(n974), .B(G4), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(G1341), .B(G19), .ZN(n976) );
  XNOR2_X1 U1072 ( .A(G1981), .B(G6), .ZN(n975) );
  NOR2_X1 U1073 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(G20), .B(G1956), .ZN(n979) );
  NOR2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1077 ( .A(KEYINPUT60), .B(n981), .ZN(n982) );
  NAND2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n986) );
  XOR2_X1 U1079 ( .A(KEYINPUT123), .B(G1966), .Z(n984) );
  XNOR2_X1 U1080 ( .A(G21), .B(n984), .ZN(n985) );
  NOR2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1082 ( .A(KEYINPUT124), .B(n987), .Z(n988) );
  NOR2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1084 ( .A(KEYINPUT61), .B(n990), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(KEYINPUT125), .B(n995), .ZN(n996) );
  NAND2_X1 U1088 ( .A1(n996), .A2(G11), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(n999), .B(KEYINPUT126), .ZN(n1027) );
  XOR2_X1 U1091 ( .A(G2072), .B(n1000), .Z(n1002) );
  XOR2_X1 U1092 ( .A(G164), .B(G2078), .Z(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1094 ( .A(KEYINPUT50), .B(n1003), .Z(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1016) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1014) );
  XNOR2_X1 U1097 ( .A(G160), .B(G2084), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1100 ( .A(KEYINPUT116), .B(n1012), .Z(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1021) );
  XOR2_X1 U1103 ( .A(G2090), .B(G162), .Z(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(n1019), .B(KEYINPUT51), .ZN(n1020) );
  NOR2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(KEYINPUT52), .B(n1022), .ZN(n1024) );
  INV_X1 U1108 ( .A(KEYINPUT55), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(G29), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
  INV_X1 U1114 ( .A(n1029), .ZN(G299) );
endmodule

