//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n611, new_n612, new_n615, new_n617, new_n618, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT68), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(KEYINPUT3), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n470), .A2(G137), .A3(new_n461), .A4(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT68), .B(G2104), .ZN(new_n474));
  INV_X1    g049(.A(G101), .ZN(new_n475));
  NOR4_X1   g050(.A1(new_n474), .A2(KEYINPUT69), .A3(new_n475), .A4(G2105), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n467), .B2(new_n469), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G101), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n473), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI211_X1 g057(.A(KEYINPUT70), .B(new_n473), .C1(new_n476), .C2(new_n479), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n465), .B1(new_n482), .B2(new_n483), .ZN(G160));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n470), .A2(new_n472), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n471), .B1(new_n474), .B2(KEYINPUT3), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n488), .A2(KEYINPUT71), .A3(new_n461), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n486), .A2(new_n461), .ZN(new_n492));
  OR2_X1    g067(.A1(new_n461), .A2(G112), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n492), .A2(G124), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n491), .A2(new_n496), .ZN(G162));
  INV_X1    g072(.A(KEYINPUT72), .ZN(new_n498));
  AND2_X1   g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n488), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n470), .A2(new_n472), .A3(new_n499), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT72), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G138), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(G2105), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n470), .A2(new_n472), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  NOR3_X1   g082(.A1(new_n504), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n462), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n511));
  INV_X1    g086(.A(G114), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(G2105), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n503), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n518), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n518), .A2(G543), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n524), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n520), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G50), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n528), .A2(new_n529), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n522), .A2(new_n523), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(G88), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n527), .A2(new_n536), .ZN(G166));
  NAND3_X1  g112(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n530), .A2(G51), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n533), .A2(G89), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(G168));
  AOI22_X1  g119(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n526), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n530), .A2(G52), .ZN(new_n547));
  XNOR2_X1  g122(.A(KEYINPUT74), .B(G90), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n534), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(G171));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n522), .A2(new_n523), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n526), .B1(new_n554), .B2(KEYINPUT75), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n555), .B1(KEYINPUT75), .B2(new_n554), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n533), .A2(G81), .B1(G43), .B2(new_n530), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(new_n530), .A2(G53), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  XOR2_X1   g142(.A(new_n567), .B(KEYINPUT76), .Z(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n552), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G651), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n533), .A2(G91), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n566), .A2(new_n571), .A3(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  INV_X1    g150(.A(G166), .ZN(G303));
  AOI22_X1  g151(.A1(new_n533), .A2(G87), .B1(G49), .B2(new_n530), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(new_n530), .A2(G48), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT77), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n530), .A2(new_n582), .A3(G48), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n581), .A2(new_n583), .B1(new_n533), .B2(G86), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n552), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n526), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n530), .A2(G47), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n534), .B2(new_n593), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n591), .A2(new_n594), .ZN(G290));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NOR2_X1   g171(.A1(G301), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n533), .A2(G92), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  XOR2_X1   g176(.A(KEYINPUT78), .B(G66), .Z(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n552), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(G54), .B2(new_n530), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT79), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n597), .B1(new_n606), .B2(new_n596), .ZN(G284));
  AOI21_X1  g182(.A(new_n597), .B1(new_n606), .B2(new_n596), .ZN(G321));
  NOR2_X1   g183(.A1(G168), .A2(new_n596), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT80), .ZN(new_n610));
  AOI21_X1  g185(.A(G868), .B1(G299), .B2(KEYINPUT81), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(KEYINPUT81), .B2(G299), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n612), .ZN(G297));
  NAND2_X1  g188(.A1(new_n610), .A2(new_n612), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n606), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n606), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g194(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n620));
  XNOR2_X1  g195(.A(G323), .B(new_n620), .ZN(G282));
  NAND2_X1  g196(.A1(new_n478), .A2(new_n462), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT12), .Z(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT13), .Z(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT83), .B(G2100), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT85), .Z(new_n627));
  NOR2_X1   g202(.A1(new_n624), .A2(new_n625), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT84), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n490), .A2(G135), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n461), .A2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  AOI22_X1  g208(.A1(new_n492), .A2(G123), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  AND2_X1   g209(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2096), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n627), .A2(new_n629), .A3(new_n636), .ZN(G156));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n641), .B(new_n647), .Z(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  AND3_X1   g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  NAND3_X1  g231(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT18), .Z(new_n658));
  INV_X1    g233(.A(new_n655), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n656), .B1(new_n659), .B2(new_n653), .ZN(new_n660));
  XOR2_X1   g235(.A(KEYINPUT86), .B(KEYINPUT17), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n653), .B(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n660), .B1(new_n663), .B2(new_n659), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(new_n659), .A3(new_n656), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n658), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2096), .B(G2100), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1961), .B(G1966), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n671), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(KEYINPUT87), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(new_n674), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT20), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G229));
  NAND2_X1  g262(.A1(G162), .A2(G29), .ZN(new_n688));
  OR2_X1    g263(.A1(G29), .A2(G35), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT102), .B(KEYINPUT29), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G2090), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G19), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(new_n559), .B2(new_n694), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n693), .B1(G1341), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n635), .A2(G29), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT100), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT30), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n700), .A2(G28), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n700), .B2(G28), .ZN(new_n703));
  AND2_X1   g278(.A1(KEYINPUT31), .A2(G11), .ZN(new_n704));
  NOR2_X1   g279(.A1(KEYINPUT31), .A2(G11), .ZN(new_n705));
  OAI22_X1  g280(.A1(new_n701), .A2(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n694), .A2(G21), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G168), .B2(new_n694), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n706), .B1(new_n708), .B2(G1966), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n699), .B(new_n709), .C1(G1966), .C2(new_n708), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n694), .A2(G20), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT23), .ZN(new_n712));
  INV_X1    g287(.A(G299), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n694), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(G1956), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n694), .A2(G5), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G171), .B2(new_n694), .ZN(new_n717));
  INV_X1    g292(.A(G1961), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g295(.A1(new_n697), .A2(new_n710), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n492), .A2(G128), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT95), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n490), .A2(G140), .ZN(new_n724));
  OR2_X1    g299(.A1(G104), .A2(G2105), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n725), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n702), .A2(G26), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT28), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT96), .B(G2067), .Z(new_n732));
  AND2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n696), .A2(G1341), .ZN(new_n735));
  NOR3_X1   g310(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n721), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n606), .A2(G16), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT94), .ZN(new_n739));
  OR3_X1    g314(.A1(new_n739), .A2(G4), .A3(G16), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(G4), .B2(G16), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1348), .ZN(new_n743));
  INV_X1    g318(.A(G34), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n744), .A2(KEYINPUT24), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(KEYINPUT24), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n702), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G160), .B2(new_n702), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT98), .ZN(new_n749));
  INV_X1    g324(.A(G2084), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n743), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT25), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n462), .A2(G127), .ZN(new_n756));
  INV_X1    g331(.A(G115), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(new_n466), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n461), .B1(new_n758), .B2(KEYINPUT97), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT97), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n756), .B(new_n760), .C1(new_n757), .C2(new_n466), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n755), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n490), .ZN(new_n763));
  INV_X1    g338(.A(G139), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  MUX2_X1   g340(.A(G33), .B(new_n765), .S(G29), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n490), .A2(G141), .ZN(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT26), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n478), .A2(G105), .ZN(new_n770));
  AOI211_X1 g345(.A(new_n769), .B(new_n770), .C1(new_n492), .C2(G129), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G29), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n702), .A2(G32), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT27), .B(G1996), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT99), .Z(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g353(.A1(G2072), .A2(new_n766), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n775), .A2(new_n778), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n779), .B(new_n780), .C1(G2072), .C2(new_n766), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n702), .A2(G27), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G164), .B2(new_n702), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT101), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n781), .B1(G2078), .B2(new_n784), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(G2078), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n737), .A2(new_n753), .A3(new_n787), .A4(KEYINPUT103), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT103), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n721), .A2(new_n785), .A3(new_n786), .A4(new_n736), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n743), .A2(new_n751), .A3(new_n752), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n694), .A2(G23), .ZN(new_n794));
  INV_X1    g369(.A(G288), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n694), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT91), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT33), .B(G1976), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT92), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n797), .A2(new_n800), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n694), .A2(G22), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G166), .B2(new_n694), .ZN(new_n804));
  INV_X1    g379(.A(G1971), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G6), .B(G305), .S(G16), .Z(new_n807));
  XOR2_X1   g382(.A(KEYINPUT32), .B(G1981), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n801), .A2(new_n802), .A3(new_n806), .A4(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT34), .ZN(new_n811));
  NOR2_X1   g386(.A1(G16), .A2(G24), .ZN(new_n812));
  INV_X1    g387(.A(G290), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(G16), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n814), .A2(G1986), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(G1986), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n815), .A2(KEYINPUT93), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n490), .A2(G131), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT88), .Z(new_n819));
  OR2_X1    g394(.A1(G95), .A2(G2105), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n820), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT89), .Z(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G119), .B2(new_n492), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(new_n702), .ZN(new_n825));
  NOR2_X1   g400(.A1(G25), .A2(G29), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT35), .B(G1991), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT90), .ZN(new_n828));
  OR3_X1    g403(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n825), .B2(new_n826), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n817), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n810), .A2(KEYINPUT34), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n811), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT36), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n793), .A2(new_n834), .ZN(G311));
  INV_X1    g410(.A(KEYINPUT104), .ZN(new_n836));
  AND3_X1   g411(.A1(new_n793), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n836), .B1(new_n793), .B2(new_n834), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(G150));
  AOI22_X1  g414(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n840), .A2(new_n526), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n530), .A2(G55), .ZN(new_n842));
  INV_X1    g417(.A(G93), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n534), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT105), .B(G860), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT37), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n606), .A2(G559), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT38), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n841), .A2(new_n844), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n558), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n845), .A2(new_n556), .A3(new_n557), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n850), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(new_n846), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n855), .A2(new_n856), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n848), .B1(new_n858), .B2(new_n859), .ZN(G145));
  INV_X1    g435(.A(KEYINPUT40), .ZN(new_n861));
  INV_X1    g436(.A(new_n623), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n824), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n765), .B(new_n772), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n513), .B1(new_n500), .B2(new_n502), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT107), .ZN(new_n867));
  AOI221_X4 g442(.A(new_n867), .B1(new_n462), .B2(new_n508), .C1(new_n506), .C2(KEYINPUT4), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT107), .B1(new_n507), .B2(new_n509), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n727), .B(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n492), .A2(G130), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n461), .A2(G118), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(G142), .B2(new_n490), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n871), .B(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n865), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n865), .A2(new_n877), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n635), .B(KEYINPUT106), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(G160), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G162), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n878), .A2(new_n879), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n883), .B1(new_n878), .B2(new_n879), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n861), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n889), .A2(KEYINPUT40), .A3(new_n885), .A4(new_n884), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n888), .A2(new_n890), .ZN(G395));
  XOR2_X1   g466(.A(new_n617), .B(new_n854), .Z(new_n892));
  NAND2_X1  g467(.A1(new_n605), .A2(new_n713), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n600), .A2(G299), .A3(new_n604), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT109), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n897), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT109), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n893), .A2(new_n901), .A3(new_n894), .ZN(new_n902));
  INV_X1    g477(.A(new_n605), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n903), .A2(KEYINPUT108), .A3(G299), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n897), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n898), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n892), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n617), .B(new_n854), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n902), .A2(new_n904), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n911), .A2(KEYINPUT42), .ZN(new_n912));
  XOR2_X1   g487(.A(G290), .B(G305), .Z(new_n913));
  XNOR2_X1  g488(.A(G166), .B(G288), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n913), .B(new_n914), .Z(new_n915));
  NAND2_X1  g490(.A1(new_n911), .A2(KEYINPUT42), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n912), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n915), .B1(new_n912), .B2(new_n916), .ZN(new_n918));
  OAI21_X1  g493(.A(G868), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n851), .A2(new_n596), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(G295));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n920), .ZN(G331));
  AND3_X1   g497(.A1(new_n852), .A2(G301), .A3(new_n853), .ZN(new_n923));
  AOI21_X1  g498(.A(G301), .B1(new_n852), .B2(new_n853), .ZN(new_n924));
  OAI21_X1  g499(.A(G286), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n854), .A2(G171), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n852), .A2(G301), .A3(new_n853), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(G168), .A3(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n893), .A2(KEYINPUT41), .A3(new_n894), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT111), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n925), .A2(new_n928), .A3(KEYINPUT41), .ZN(new_n933));
  INV_X1    g508(.A(new_n909), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI211_X1 g510(.A(KEYINPUT112), .B(new_n915), .C1(new_n932), .C2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT112), .ZN(new_n937));
  AOI22_X1  g512(.A1(new_n929), .A2(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n938));
  INV_X1    g513(.A(new_n915), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT110), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n934), .B1(new_n925), .B2(new_n928), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n943), .B1(new_n906), .B2(new_n929), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n942), .B1(new_n944), .B2(new_n915), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n929), .A2(new_n906), .ZN(new_n946));
  INV_X1    g521(.A(new_n943), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n915), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(G37), .B1(new_n948), .B2(KEYINPUT110), .ZN(new_n949));
  AND4_X1   g524(.A1(KEYINPUT43), .A2(new_n941), .A3(new_n945), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n946), .A2(new_n947), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(KEYINPUT110), .A3(new_n939), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n944), .A2(new_n915), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n945), .A2(new_n952), .A3(new_n885), .A4(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT44), .B1(new_n950), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n941), .A2(new_n955), .A3(new_n945), .A4(new_n949), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n957), .A2(new_n962), .ZN(G397));
  INV_X1    g538(.A(KEYINPUT123), .ZN(new_n964));
  INV_X1    g539(.A(G8), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n966));
  OAI22_X1  g541(.A1(G168), .A2(new_n965), .B1(KEYINPUT122), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1966), .ZN(new_n969));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n870), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G40), .ZN(new_n974));
  AOI211_X1 g549(.A(new_n974), .B(new_n465), .C1(new_n482), .C2(new_n483), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n972), .A2(G1384), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n515), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n870), .A2(new_n979), .A3(new_n970), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n498), .B1(new_n488), .B2(new_n499), .ZN(new_n981));
  AND4_X1   g556(.A1(new_n498), .A2(new_n470), .A3(new_n472), .A4(new_n499), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n514), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n507), .A2(new_n509), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n970), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT50), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n975), .A2(new_n980), .A3(new_n986), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n969), .A2(new_n978), .B1(new_n987), .B2(new_n750), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n968), .B1(new_n988), .B2(new_n965), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n966), .A2(KEYINPUT122), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n988), .ZN(new_n992));
  NOR2_X1   g567(.A1(G168), .A2(new_n965), .ZN(new_n993));
  AOI22_X1  g568(.A1(new_n989), .A2(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n968), .B(new_n990), .C1(new_n988), .C2(new_n965), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n964), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n978), .A2(new_n969), .ZN(new_n997));
  INV_X1    g572(.A(new_n465), .ZN(new_n998));
  INV_X1    g573(.A(new_n483), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n468), .A2(G2104), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n466), .A2(KEYINPUT68), .ZN(new_n1001));
  OAI211_X1 g576(.A(G101), .B(new_n461), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT69), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n478), .A2(new_n477), .A3(G101), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT70), .B1(new_n1005), .B2(new_n473), .ZN(new_n1006));
  OAI211_X1 g581(.A(G40), .B(new_n998), .C1(new_n999), .C2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n979), .B1(new_n515), .B2(new_n970), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1009), .A2(new_n750), .A3(new_n980), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n965), .B1(new_n997), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n991), .B1(new_n1011), .B2(new_n967), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n992), .A2(new_n993), .ZN(new_n1013));
  AND4_X1   g588(.A1(new_n964), .A2(new_n1012), .A3(new_n995), .A4(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT62), .B1(new_n996), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1016));
  INV_X1    g591(.A(new_n995), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT123), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n994), .A2(new_n964), .A3(new_n995), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT62), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n510), .A2(new_n867), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n507), .A2(KEYINPUT107), .A3(new_n509), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1384), .B1(new_n1025), .B2(new_n866), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n975), .B(new_n1022), .C1(new_n1026), .C2(new_n979), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n979), .B1(new_n870), .B2(new_n970), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT116), .B1(new_n1028), .B2(new_n1007), .ZN(new_n1029));
  INV_X1    g604(.A(G2090), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1384), .B1(new_n866), .B2(new_n510), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n979), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .A4(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n985), .A2(new_n972), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n870), .A2(new_n976), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n975), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n805), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1033), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(G8), .ZN(new_n1039));
  NAND2_X1  g614(.A1(G303), .A2(G8), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n1041));
  OR3_X1    g616(.A1(new_n1040), .A2(KEYINPUT115), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT115), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1039), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1037), .A2(KEYINPUT114), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1036), .A2(new_n1049), .A3(new_n805), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n987), .A2(new_n1030), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(G8), .A3(new_n1045), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n975), .A2(new_n1026), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n795), .A2(G1976), .ZN(new_n1055));
  INV_X1    g630(.A(G1976), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT52), .B1(G288), .B2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1054), .A2(G8), .A3(new_n1055), .A4(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1981), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(new_n584), .B2(new_n588), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n584), .A2(new_n1059), .A3(new_n588), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(KEYINPUT49), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT49), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1062), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1064), .B1(new_n1065), .B2(new_n1060), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1054), .A2(G8), .A3(new_n1063), .A4(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(G8), .B(new_n1055), .C1(new_n971), .C2(new_n1007), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT52), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1058), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1058), .A2(new_n1067), .A3(new_n1069), .A4(KEYINPUT117), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1047), .A2(new_n1053), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G2078), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n975), .A2(new_n1034), .A3(new_n1035), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(G160), .B(G40), .C1(new_n979), .C2(new_n1031), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n870), .A2(new_n979), .A3(new_n970), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n718), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1078), .A2(G2078), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n973), .A2(new_n975), .A3(new_n977), .A4(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1079), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1085), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT124), .B1(new_n1085), .B2(G171), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1075), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1015), .A2(new_n1021), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1007), .B1(new_n971), .B2(new_n972), .ZN(new_n1091));
  AOI21_X1  g666(.A(G1966), .B1(new_n1091), .B2(new_n977), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1080), .A2(new_n1081), .A3(G2084), .ZN(new_n1093));
  OAI211_X1 g668(.A(G8), .B(G168), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1047), .A2(new_n1053), .A3(new_n1074), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT63), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1058), .A2(new_n1067), .A3(new_n1069), .A4(KEYINPUT63), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1094), .A2(new_n1099), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1053), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1052), .A2(G8), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1046), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1098), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1053), .A2(new_n1070), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1067), .A2(new_n1056), .A3(new_n795), .ZN(new_n1108));
  OAI211_X1 g683(.A(G8), .B(new_n1054), .C1(new_n1108), .C2(new_n1065), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1105), .A2(new_n1106), .A3(new_n1111), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1096), .A2(new_n1097), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT118), .B1(new_n1113), .B2(new_n1110), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT120), .B(G1996), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n975), .A2(new_n1034), .A3(new_n1035), .A4(new_n1115), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n1117));
  XNOR2_X1  g692(.A(new_n1117), .B(G1341), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n971), .B2(new_n1007), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n558), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1120), .B(KEYINPUT59), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n1122));
  AOI21_X1  g697(.A(G1348), .B1(new_n1009), .B2(new_n980), .ZN(new_n1123));
  INV_X1    g698(.A(G2067), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n975), .A2(new_n1026), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n903), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1125), .B(new_n605), .C1(new_n987), .C2(G1348), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1122), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NOR4_X1   g704(.A1(new_n1123), .A2(new_n1126), .A3(KEYINPUT60), .A4(new_n605), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1121), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n1132));
  XOR2_X1   g707(.A(G299), .B(KEYINPUT57), .Z(new_n1133));
  NAND3_X1  g708(.A1(new_n1027), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT119), .B(G1956), .Z(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT56), .B(G2072), .Z(new_n1138));
  NOR2_X1   g713(.A1(new_n1036), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1133), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1133), .ZN(new_n1142));
  AOI211_X1 g717(.A(new_n1142), .B(new_n1139), .C1(new_n1134), .C2(new_n1136), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1132), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1007), .B1(new_n971), .B2(KEYINPUT50), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1145), .A2(new_n1022), .B1(new_n979), .B2(new_n1031), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1135), .B1(new_n1146), .B2(new_n1029), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1142), .B1(new_n1147), .B2(new_n1139), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1137), .A2(new_n1133), .A3(new_n1140), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(KEYINPUT61), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1131), .A2(new_n1144), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1127), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1149), .B1(new_n1141), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1091), .A2(new_n1035), .A3(new_n1083), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(new_n1079), .A3(new_n1082), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1156), .A2(G171), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT54), .B1(new_n1088), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(G171), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1079), .A2(new_n1082), .A3(new_n1084), .A4(G301), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(KEYINPUT54), .A3(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1047), .A2(new_n1161), .A3(new_n1053), .A4(new_n1074), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1158), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1154), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1090), .A2(new_n1112), .A3(new_n1114), .A4(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n975), .A2(new_n972), .A3(new_n971), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n824), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n827), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n727), .B(new_n1124), .ZN(new_n1172));
  XOR2_X1   g747(.A(new_n772), .B(G1996), .Z(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1169), .A2(new_n827), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1171), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(G290), .A2(G1986), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT113), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(G1986), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1180), .B1(new_n1181), .B2(new_n813), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1168), .B1(new_n1177), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1166), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT48), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(new_n1180), .B2(new_n1167), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1179), .A2(KEYINPUT48), .A3(new_n1168), .ZN(new_n1187));
  OAI211_X1 g762(.A(new_n1186), .B(new_n1187), .C1(new_n1176), .C2(new_n1167), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT46), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1190), .B1(new_n1167), .B2(G1996), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT125), .ZN(new_n1192));
  INV_X1    g767(.A(new_n772), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1172), .B(new_n1193), .C1(new_n1190), .C2(G1996), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1192), .B1(new_n1194), .B2(new_n1168), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1195), .B(KEYINPUT47), .ZN(new_n1196));
  OAI22_X1  g771(.A1(new_n1170), .A2(new_n1174), .B1(G2067), .B2(new_n727), .ZN(new_n1197));
  AOI211_X1 g772(.A(new_n1189), .B(new_n1196), .C1(new_n1168), .C2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1184), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g774(.A1(new_n889), .A2(new_n885), .A3(new_n884), .ZN(new_n1201));
  INV_X1    g775(.A(new_n459), .ZN(new_n1202));
  NOR3_X1   g776(.A1(G401), .A2(new_n1202), .A3(G227), .ZN(new_n1203));
  XOR2_X1   g777(.A(new_n1203), .B(KEYINPUT126), .Z(new_n1204));
  NOR2_X1   g778(.A1(new_n1204), .A2(G229), .ZN(new_n1205));
  AND3_X1   g779(.A1(new_n1201), .A2(new_n960), .A3(new_n1205), .ZN(G308));
  NAND3_X1  g780(.A1(new_n1201), .A2(new_n960), .A3(new_n1205), .ZN(G225));
endmodule


