//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1288, new_n1289, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346, new_n1347;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(KEYINPUT64), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT64), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n215), .A2(G1), .A3(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G20), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n212), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(new_n209), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n220), .B(new_n228), .C1(KEYINPUT1), .C2(new_n226), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XNOR2_X1  g0037(.A(G68), .B(G77), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT66), .B(G50), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  XNOR2_X1  g0045(.A(KEYINPUT3), .B(G33), .ZN(new_n246));
  INV_X1    g0046(.A(G1698), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n246), .A2(G222), .A3(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G77), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n246), .A2(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(G223), .ZN(new_n251));
  OAI221_X1 g0051(.A(new_n248), .B1(new_n249), .B2(new_n246), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  AND2_X1   g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n253), .B1(new_n214), .B2(new_n216), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT67), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT68), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(new_n253), .B2(new_n213), .ZN(new_n262));
  AND2_X1   g0062(.A1(G1), .A2(G13), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(KEYINPUT68), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n260), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n257), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n268), .B1(new_n262), .B2(new_n265), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G226), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n255), .A2(new_n267), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G169), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G20), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n277), .B(KEYINPUT69), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n214), .A2(new_n216), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n280), .A2(new_n282), .B1(new_n202), .B2(new_n284), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n214), .A2(new_n216), .A3(new_n283), .A4(new_n281), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G20), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(G1), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(G50), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n273), .B(new_n292), .C1(G179), .C2(new_n271), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n285), .A2(KEYINPUT9), .A3(new_n291), .ZN(new_n295));
  XOR2_X1   g0095(.A(new_n295), .B(KEYINPUT70), .Z(new_n296));
  INV_X1    g0096(.A(new_n271), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT9), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n297), .A2(G190), .B1(new_n292), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G200), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT71), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  OR3_X1    g0101(.A1(new_n297), .A2(KEYINPUT71), .A3(new_n300), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n296), .A2(new_n299), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n302), .A2(new_n299), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n305), .A2(new_n306), .A3(new_n296), .A4(new_n301), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n294), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT13), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G33), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n310), .A2(new_n312), .A3(G232), .A4(G1698), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n310), .A2(new_n312), .A3(G226), .A4(new_n247), .ZN(new_n314));
  NAND2_X1  g0114(.A1(G33), .A2(G97), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n254), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT72), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT72), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(new_n254), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n266), .A2(new_n259), .B1(new_n269), .B2(G238), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n309), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n316), .A2(new_n254), .A3(new_n319), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n319), .B1(new_n316), .B2(new_n254), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n309), .B(new_n322), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(G169), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT14), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n322), .B1(new_n324), .B2(new_n325), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT13), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(G179), .A3(new_n326), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n326), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT14), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(new_n334), .A3(G169), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n329), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G68), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n274), .A2(G50), .B1(G20), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n278), .B2(new_n249), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n282), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT11), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n339), .A2(KEYINPUT11), .A3(new_n282), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n286), .A2(new_n337), .A3(new_n289), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT12), .B1(new_n283), .B2(G68), .ZN(new_n345));
  OR3_X1    g0145(.A1(new_n283), .A2(KEYINPUT12), .A3(G68), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n342), .A2(new_n343), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT74), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n342), .A2(KEYINPUT74), .A3(new_n343), .A4(new_n347), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n336), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n331), .A2(G190), .A3(new_n326), .ZN(new_n354));
  INV_X1    g0154(.A(new_n348), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT73), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n300), .B1(new_n331), .B2(new_n326), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n354), .A2(new_n355), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT73), .B1(new_n361), .B2(new_n358), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n246), .A2(G232), .A3(new_n247), .ZN(new_n364));
  INV_X1    g0164(.A(G238), .ZN(new_n365));
  OAI221_X1 g0165(.A(new_n364), .B1(new_n206), .B2(new_n246), .C1(new_n250), .C2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n254), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n269), .A2(G244), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n267), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(G200), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(G20), .A2(G77), .ZN(new_n372));
  INV_X1    g0172(.A(new_n274), .ZN(new_n373));
  INV_X1    g0173(.A(new_n277), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT15), .B(G87), .ZN(new_n375));
  OAI221_X1 g0175(.A(new_n372), .B1(new_n279), .B2(new_n373), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n376), .A2(new_n282), .B1(new_n249), .B2(new_n284), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n287), .A2(G77), .A3(new_n290), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n367), .A2(G190), .A3(new_n267), .A4(new_n369), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n371), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n272), .B1(new_n368), .B2(new_n370), .ZN(new_n383));
  INV_X1    g0183(.A(G179), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n367), .A2(new_n384), .A3(new_n267), .A4(new_n369), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n385), .A3(new_n379), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n308), .A2(new_n353), .A3(new_n363), .A4(new_n387), .ZN(new_n388));
  XNOR2_X1  g0188(.A(G58), .B(G68), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n389), .A2(G20), .B1(G159), .B2(new_n274), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  AOI211_X1 g0191(.A(new_n391), .B(G20), .C1(new_n310), .C2(new_n312), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n310), .A2(new_n312), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT75), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n246), .A2(KEYINPUT75), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(new_n396), .A3(new_n288), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n392), .B1(new_n397), .B2(new_n391), .ZN(new_n398));
  OAI211_X1 g0198(.A(KEYINPUT16), .B(new_n390), .C1(new_n398), .C2(new_n337), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT16), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n391), .B1(new_n246), .B2(G20), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n393), .A2(KEYINPUT7), .A3(new_n288), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n337), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n390), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n400), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n399), .A2(new_n405), .A3(new_n282), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n310), .A2(new_n312), .A3(G226), .A4(G1698), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n310), .A2(new_n312), .A3(G223), .A4(new_n247), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G87), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n254), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n269), .A2(G232), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n267), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n300), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(G190), .B2(new_n413), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n286), .A2(new_n279), .A3(new_n289), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n284), .B2(new_n279), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n406), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT17), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n406), .A2(new_n415), .A3(KEYINPUT17), .A4(new_n417), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT18), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n406), .A2(new_n417), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT76), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n413), .A2(new_n384), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n266), .A2(new_n259), .B1(new_n269), .B2(G232), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n272), .B1(new_n427), .B2(new_n411), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n425), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n413), .A2(G169), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n427), .A2(G179), .A3(new_n411), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(KEYINPUT76), .A3(new_n431), .ZN(new_n432));
  AND4_X1   g0232(.A1(new_n423), .A2(new_n424), .A3(new_n429), .A4(new_n432), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n430), .A2(KEYINPUT76), .A3(new_n431), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT76), .B1(new_n430), .B2(new_n431), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n423), .B1(new_n436), .B2(new_n424), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT77), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n433), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n424), .A2(new_n429), .A3(new_n432), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT18), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n436), .A2(new_n423), .A3(new_n424), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT77), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n422), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n388), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n282), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT7), .B1(new_n393), .B2(new_n288), .ZN(new_n447));
  OAI21_X1  g0247(.A(G107), .B1(new_n447), .B2(new_n392), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n373), .A2(new_n249), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT6), .ZN(new_n450));
  AND2_X1   g0250(.A1(G97), .A2(G107), .ZN(new_n451));
  NOR2_X1   g0251(.A1(G97), .A2(G107), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AND2_X1   g0253(.A1(KEYINPUT78), .A2(G97), .ZN(new_n454));
  NOR2_X1   g0254(.A1(KEYINPUT78), .A2(G97), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n453), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n449), .B1(new_n458), .B2(G20), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n446), .B1(new_n448), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n283), .A2(G97), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n276), .A2(G1), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n286), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n461), .B1(new_n463), .B2(G97), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT81), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n455), .ZN(new_n467));
  NAND2_X1  g0267(.A1(KEYINPUT78), .A2(G97), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n457), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G97), .A2(G107), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT6), .B1(new_n207), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(G20), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n449), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n206), .B1(new_n401), .B2(new_n402), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n282), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT81), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(new_n477), .A3(new_n464), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n310), .A2(new_n312), .A3(G244), .A4(new_n247), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT79), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT4), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n481), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n246), .A2(G244), .A3(new_n247), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n246), .A2(G250), .A3(G1698), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G283), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n482), .A2(new_n484), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n254), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n256), .A2(G45), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT5), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(G41), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT80), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(G41), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n494), .B2(KEYINPUT5), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(KEYINPUT5), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n493), .A2(new_n497), .B1(new_n262), .B2(new_n265), .ZN(new_n498));
  INV_X1    g0298(.A(G45), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(G1), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n492), .A2(new_n494), .A3(KEYINPUT5), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT80), .B1(new_n490), .B2(G41), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n500), .B(new_n501), .C1(new_n502), .C2(new_n491), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n498), .A2(G257), .B1(new_n504), .B2(new_n266), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n488), .A2(G179), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n272), .B1(new_n488), .B2(new_n505), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n466), .B(new_n478), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT82), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n488), .A2(new_n505), .A3(G179), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n262), .A2(new_n265), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n511), .A2(G274), .A3(new_n497), .A4(new_n493), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n503), .A3(G257), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(new_n254), .B2(new_n487), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n510), .B1(new_n515), .B2(new_n272), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT82), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(new_n466), .A4(new_n478), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n509), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n476), .A2(new_n464), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n488), .A2(new_n505), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(G200), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n515), .A2(G190), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n310), .A2(new_n312), .A3(G244), .A4(G1698), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n310), .A2(new_n312), .A3(G238), .A4(new_n247), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G116), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n254), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n253), .A2(new_n261), .A3(new_n213), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT68), .B1(new_n263), .B2(new_n264), .ZN(new_n532));
  OAI211_X1 g0332(.A(G274), .B(new_n500), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n489), .A2(G250), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n511), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(G200), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n246), .A2(new_n288), .A3(G68), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT19), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n456), .B2(new_n374), .ZN(new_n540));
  NOR2_X1   g0340(.A1(G87), .A2(G107), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n456), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n543), .A2(new_n288), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n538), .B(new_n540), .C1(new_n542), .C2(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n545), .A2(new_n282), .B1(new_n284), .B2(new_n375), .ZN(new_n546));
  INV_X1    g0346(.A(new_n462), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n287), .A2(G87), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT83), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n463), .A2(KEYINPUT83), .A3(G87), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n266), .A2(new_n500), .B1(new_n511), .B2(new_n534), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n553), .A2(G190), .A3(new_n529), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n537), .A2(new_n546), .A3(new_n552), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n540), .A2(new_n538), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n544), .B1(new_n456), .B2(new_n541), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n282), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n375), .A2(new_n284), .ZN(new_n559));
  INV_X1    g0359(.A(new_n375), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n463), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n272), .B1(new_n530), .B2(new_n536), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n553), .A2(new_n384), .A3(new_n529), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n555), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n310), .A2(new_n312), .A3(new_n288), .A4(G87), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT22), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT22), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n246), .A2(new_n569), .A3(new_n288), .A4(G87), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT24), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n527), .A2(G20), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT23), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n288), .B2(G107), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n571), .A2(new_n572), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n572), .B1(new_n571), .B2(new_n577), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n282), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT25), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n283), .B2(G107), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n284), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n463), .A2(G107), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n246), .A2(G257), .A3(G1698), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n246), .A2(G250), .A3(new_n247), .ZN(new_n587));
  INV_X1    g0387(.A(G294), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n586), .B(new_n587), .C1(new_n276), .C2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n254), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT85), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n498), .B2(G264), .ZN(new_n592));
  AND4_X1   g0392(.A1(new_n591), .A2(new_n511), .A3(new_n503), .A4(G264), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n590), .B(new_n512), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(G190), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n585), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(G200), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n566), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n519), .A2(new_n524), .A3(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n310), .A2(new_n312), .A3(G264), .A4(G1698), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n310), .A2(new_n312), .A3(G257), .A4(new_n247), .ZN(new_n602));
  INV_X1    g0402(.A(G303), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n601), .B(new_n602), .C1(new_n603), .C2(new_n246), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n254), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n511), .A2(new_n503), .A3(G270), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n512), .A3(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n607), .A2(G169), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT20), .ZN(new_n609));
  INV_X1    g0409(.A(G116), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(G20), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n282), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n486), .A2(new_n288), .ZN(new_n613));
  XNOR2_X1  g0413(.A(KEYINPUT78), .B(G97), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n614), .B2(new_n276), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n609), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n613), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n456), .B2(G33), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(KEYINPUT20), .A3(new_n282), .A4(new_n611), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT84), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n283), .A2(G116), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n463), .B2(G116), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n620), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n621), .B1(new_n620), .B2(new_n623), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n608), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT21), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n620), .A2(new_n623), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT84), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n620), .A2(new_n621), .A3(new_n623), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n607), .A2(KEYINPUT21), .A3(G169), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n605), .A2(G179), .A3(new_n512), .A4(new_n606), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n605), .A2(new_n512), .A3(new_n606), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(G190), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n607), .A2(G200), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n630), .A2(new_n638), .A3(new_n631), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n511), .A2(new_n503), .ZN(new_n641));
  INV_X1    g0441(.A(G264), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT85), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n498), .A2(new_n591), .A3(G264), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n645), .A2(new_n384), .A3(new_n512), .A4(new_n590), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n594), .A2(new_n272), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n585), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AND4_X1   g0448(.A1(new_n628), .A2(new_n636), .A3(new_n640), .A4(new_n648), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n445), .A2(new_n600), .A3(new_n649), .ZN(G372));
  NOR2_X1   g0450(.A1(new_n426), .A2(new_n428), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n424), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT18), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n651), .B1(new_n406), .B2(new_n417), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n423), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n386), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n361), .B2(new_n358), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n353), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT87), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n422), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n353), .A2(new_n661), .A3(new_n659), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n657), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n304), .A2(new_n307), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n294), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n516), .A2(new_n520), .A3(new_n555), .A4(new_n565), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n565), .B1(new_n667), .B2(KEYINPUT26), .ZN(new_n668));
  INV_X1    g0468(.A(new_n566), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n509), .A2(new_n518), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n668), .B1(new_n670), .B2(KEYINPUT26), .ZN(new_n671));
  INV_X1    g0471(.A(new_n648), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT86), .ZN(new_n673));
  AOI21_X1  g0473(.A(KEYINPUT21), .B1(new_n632), .B2(new_n608), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n630), .A2(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n628), .A2(KEYINPUT86), .A3(new_n636), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n519), .A2(new_n599), .A3(new_n524), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n671), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n445), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n666), .B1(new_n681), .B2(new_n682), .ZN(G369));
  NAND3_X1  g0483(.A1(new_n256), .A2(new_n288), .A3(G13), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n632), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n690), .B1(new_n676), .B2(new_n677), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n674), .A2(new_n675), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n640), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n691), .B1(new_n693), .B2(new_n690), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT88), .Z(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n648), .A2(new_n689), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n597), .A2(new_n598), .B1(new_n585), .B2(new_n689), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n698), .B1(new_n700), .B2(new_n648), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n692), .A2(new_n689), .ZN(new_n703));
  XOR2_X1   g0503(.A(new_n703), .B(KEYINPUT89), .Z(new_n704));
  AOI21_X1  g0504(.A(new_n698), .B1(new_n704), .B2(new_n701), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n702), .A2(new_n705), .ZN(G399));
  NAND2_X1  g0506(.A1(new_n542), .A2(new_n610), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n210), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n219), .B2(new_n711), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n628), .A2(new_n636), .A3(new_n648), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n519), .A2(new_n715), .A3(new_n599), .A4(new_n524), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT26), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n509), .A2(new_n717), .A3(new_n518), .A4(new_n669), .ZN(new_n718));
  INV_X1    g0518(.A(new_n565), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n667), .B2(KEYINPUT26), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n716), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT90), .ZN(new_n722));
  INV_X1    g0522(.A(new_n689), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n722), .B1(new_n721), .B2(new_n723), .ZN(new_n725));
  OAI21_X1  g0525(.A(KEYINPUT29), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n681), .B2(new_n689), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n637), .A2(G179), .A3(new_n488), .A4(new_n505), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n645), .A2(new_n529), .A3(new_n553), .A4(new_n590), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n521), .A2(new_n634), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n590), .B1(new_n592), .B2(new_n593), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n553), .A2(new_n529), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n733), .A2(new_n736), .A3(KEYINPUT30), .ZN(new_n737));
  AOI21_X1  g0537(.A(G179), .B1(new_n553), .B2(new_n529), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n594), .A2(new_n521), .A3(new_n607), .A4(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n732), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n740), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n741));
  AOI21_X1  g0541(.A(KEYINPUT31), .B1(new_n740), .B2(new_n689), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n509), .A2(new_n518), .B1(new_n523), .B2(new_n522), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(new_n649), .A3(new_n599), .A4(new_n723), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n726), .A2(new_n728), .B1(G330), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT91), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n714), .B1(new_n748), .B2(G1), .ZN(G364));
  INV_X1    g0549(.A(G13), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n256), .B1(new_n751), .B2(G45), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n710), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n697), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G330), .B2(new_n695), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n217), .B1(new_n288), .B2(G169), .ZN(new_n757));
  NAND3_X1  g0557(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n595), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n288), .A2(G190), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n384), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n760), .A2(new_n202), .B1(new_n763), .B2(new_n249), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n288), .A2(new_n595), .ZN(new_n765));
  AND3_X1   g0565(.A1(new_n765), .A2(KEYINPUT94), .A3(new_n762), .ZN(new_n766));
  AOI21_X1  g0566(.A(KEYINPUT94), .B1(new_n765), .B2(new_n762), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n764), .B1(new_n769), .B2(G58), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT95), .Z(new_n771));
  NOR2_X1   g0571(.A1(new_n300), .A2(G179), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n761), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G107), .ZN(new_n775));
  INV_X1    g0575(.A(G87), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n765), .A2(new_n772), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n775), .B(new_n246), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n758), .A2(G190), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G179), .A2(G200), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n288), .B1(new_n781), .B2(G190), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n780), .A2(new_n337), .B1(new_n782), .B2(new_n205), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n761), .A2(new_n781), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G159), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT32), .ZN(new_n787));
  OR4_X1    g0587(.A1(new_n771), .A2(new_n778), .A3(new_n783), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n782), .A2(new_n588), .ZN(new_n789));
  INV_X1    g0589(.A(new_n763), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n246), .B1(new_n790), .B2(G311), .ZN(new_n791));
  INV_X1    g0591(.A(G283), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n791), .B1(new_n792), .B2(new_n773), .C1(new_n603), .C2(new_n777), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n789), .B(new_n793), .C1(G326), .C2(new_n759), .ZN(new_n794));
  XNOR2_X1  g0594(.A(KEYINPUT33), .B(G317), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n780), .B1(KEYINPUT97), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(KEYINPUT97), .B2(new_n796), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n784), .B(KEYINPUT96), .Z(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G329), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n769), .A2(G322), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n794), .A2(new_n798), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n757), .B1(new_n788), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n754), .ZN(new_n804));
  INV_X1    g0604(.A(new_n757), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G13), .A2(G33), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(G20), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n395), .A2(new_n396), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n210), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT93), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n241), .A2(G45), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(G45), .C2(new_n219), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n709), .A2(new_n393), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT92), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n818), .A2(G355), .B1(new_n610), .B2(new_n709), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n810), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n803), .A2(new_n804), .A3(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n808), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n695), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n756), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  NAND2_X1  g0625(.A1(new_n379), .A2(new_n689), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n382), .A2(new_n386), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(KEYINPUT99), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT99), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n382), .A2(new_n386), .A3(new_n829), .A4(new_n826), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n658), .A2(new_n689), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n681), .B2(new_n689), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n689), .B1(new_n828), .B2(new_n830), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n680), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n746), .A2(G330), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n754), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n837), .B2(new_n836), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n805), .A2(new_n806), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n754), .B1(new_n841), .B2(G77), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n790), .A2(G159), .B1(G137), .B2(new_n759), .ZN(new_n843));
  INV_X1    g0643(.A(G150), .ZN(new_n844));
  INV_X1    g0644(.A(G143), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n843), .B1(new_n844), .B2(new_n780), .C1(new_n768), .C2(new_n845), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT34), .Z(new_n847));
  NAND2_X1  g0647(.A1(new_n799), .A2(G132), .ZN(new_n848));
  INV_X1    g0648(.A(new_n782), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(G58), .ZN(new_n850));
  INV_X1    g0650(.A(new_n777), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n851), .A2(G50), .B1(new_n774), .B2(G68), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n848), .A2(new_n811), .A3(new_n850), .A4(new_n852), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n768), .A2(new_n588), .B1(new_n205), .B2(new_n782), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT98), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n799), .A2(G311), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n779), .A2(G283), .B1(new_n759), .B2(G303), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n246), .B1(new_n774), .B2(G87), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n851), .A2(G107), .B1(new_n790), .B2(G116), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n856), .A2(new_n857), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n847), .A2(new_n853), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n842), .B1(new_n861), .B2(new_n805), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n862), .B1(new_n863), .B2(new_n807), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n839), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(G384));
  NOR2_X1   g0666(.A1(new_n751), .A2(new_n256), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n832), .B1(new_n743), .B2(new_n745), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT40), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n350), .A2(new_n351), .A3(new_n689), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n356), .B2(new_n359), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n353), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n336), .B1(new_n362), .B2(new_n360), .ZN(new_n873));
  INV_X1    g0673(.A(new_n870), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n868), .A2(new_n869), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n390), .B1(new_n398), .B2(new_n337), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n400), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n878), .A2(new_n282), .A3(new_n399), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n417), .ZN(new_n880));
  INV_X1    g0680(.A(new_n687), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n444), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n880), .A2(new_n652), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT102), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(new_n886), .A3(new_n418), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n651), .B1(new_n879), .B2(new_n417), .ZN(new_n888));
  INV_X1    g0688(.A(new_n418), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT102), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n887), .A2(new_n890), .A3(new_n882), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n687), .B(KEYINPUT103), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n424), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n440), .A2(new_n894), .A3(new_n895), .A4(new_n418), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n884), .A2(new_n897), .A3(KEYINPUT38), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n438), .B1(new_n433), .B2(new_n437), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n441), .A2(KEYINPUT77), .A3(new_n442), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n882), .B1(new_n902), .B2(new_n422), .ZN(new_n903));
  INV_X1    g0703(.A(new_n893), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n406), .B2(new_n417), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n889), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT37), .B1(new_n436), .B2(new_n424), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n891), .A2(KEYINPUT37), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n899), .B1(new_n903), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n876), .B1(new_n898), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n868), .A2(new_n875), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n654), .A2(new_n420), .A3(new_n656), .A4(new_n421), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n905), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n889), .A2(new_n655), .A3(new_n905), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n896), .B1(new_n915), .B2(new_n895), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT104), .B1(new_n917), .B2(new_n899), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT104), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n919), .B(KEYINPUT38), .C1(new_n914), .C2(new_n916), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n903), .A2(new_n908), .A3(new_n899), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n912), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n910), .B1(new_n923), .B2(KEYINPUT40), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT105), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n445), .A2(new_n746), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(G330), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n657), .A2(new_n893), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n335), .A2(new_n332), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n363), .A2(new_n329), .A3(new_n931), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n932), .A2(new_n870), .B1(new_n353), .B2(new_n871), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT101), .ZN(new_n934));
  INV_X1    g0734(.A(new_n834), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n674), .A2(new_n673), .A3(new_n675), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT86), .B1(new_n628), .B2(new_n636), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n648), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n600), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n935), .B1(new_n939), .B2(new_n671), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n386), .A2(new_n689), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n934), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n941), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n835), .A2(KEYINPUT101), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n933), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n898), .A2(new_n909), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n930), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT39), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n921), .B2(new_n922), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n336), .A2(new_n352), .A3(new_n723), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n898), .A2(new_n909), .A3(KEYINPUT39), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n949), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n947), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n726), .A2(new_n445), .A3(new_n728), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n666), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n954), .B(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n867), .B1(new_n929), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n957), .B2(new_n929), .ZN(new_n959));
  INV_X1    g0759(.A(G58), .ZN(new_n960));
  OAI21_X1  g0760(.A(G77), .B1(new_n960), .B2(new_n337), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n961), .A2(new_n219), .B1(G50), .B2(new_n337), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(G1), .A3(new_n750), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT100), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n610), .B(new_n218), .C1(new_n458), .C2(KEYINPUT35), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(KEYINPUT35), .B2(new_n458), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT36), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n967), .B2(new_n966), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n959), .A2(new_n969), .ZN(G367));
  NAND2_X1  g0770(.A1(new_n520), .A2(new_n689), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n744), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n516), .A2(new_n520), .A3(new_n689), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT107), .Z(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n704), .A2(new_n701), .A3(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT42), .ZN(new_n977));
  INV_X1    g0777(.A(new_n975), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n519), .B1(new_n978), .B2(new_n648), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n977), .B1(new_n723), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n546), .A2(new_n552), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n669), .B1(new_n982), .B2(new_n723), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n719), .A2(new_n981), .A3(new_n689), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n980), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n985), .ZN(new_n988));
  XNOR2_X1  g0788(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  MUX2_X1   g0790(.A(new_n980), .B(new_n987), .S(new_n990), .Z(new_n991));
  NOR2_X1   g0791(.A1(new_n702), .A2(new_n978), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(KEYINPUT108), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n991), .A2(new_n993), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OR3_X1    g0796(.A1(new_n991), .A2(KEYINPUT108), .A3(new_n993), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n710), .B(KEYINPUT41), .Z(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n705), .A2(new_n975), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT45), .Z(new_n1002));
  NOR2_X1   g0802(.A1(new_n705), .A2(new_n975), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT44), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(new_n702), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n704), .B(new_n701), .Z(new_n1008));
  XNOR2_X1  g0808(.A(new_n696), .B(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT109), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n748), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1010), .B1(new_n748), .B2(new_n1009), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(KEYINPUT110), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT110), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1007), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n748), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1000), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n998), .B1(new_n1021), .B2(new_n752), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n777), .A2(new_n610), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT46), .ZN(new_n1024));
  INV_X1    g0824(.A(G311), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n760), .A2(new_n1025), .B1(new_n782), .B2(new_n206), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n769), .A2(G303), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(KEYINPUT111), .B(G317), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n773), .A2(new_n456), .B1(new_n784), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G283), .B2(new_n790), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n811), .B1(G294), .B2(new_n779), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1027), .A2(new_n1028), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n760), .A2(new_n845), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n774), .A2(G77), .B1(new_n785), .B2(G137), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1035), .B(new_n246), .C1(new_n960), .C2(new_n777), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT113), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n790), .A2(G50), .B1(G159), .B2(new_n779), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1034), .B(new_n1036), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n782), .A2(new_n337), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n769), .B2(G150), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT112), .Z(new_n1043));
  OAI21_X1  g0843(.A(new_n1033), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT47), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n805), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n988), .A2(new_n808), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n814), .A2(new_n236), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n810), .B1(new_n709), .B2(new_n560), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n804), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1046), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1022), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(G387));
  OAI21_X1  g0854(.A(new_n710), .B1(new_n748), .B2(new_n1009), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1016), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1009), .A2(new_n753), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n790), .A2(G303), .B1(G322), .B2(new_n759), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n1025), .B2(new_n780), .C1(new_n768), .C2(new_n1029), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT48), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n851), .A2(G294), .B1(new_n849), .B2(G283), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT49), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n773), .A2(new_n610), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1069), .B(new_n811), .C1(G326), .C2(new_n785), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n769), .A2(G50), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n849), .A2(new_n560), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n811), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n279), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1075), .A2(new_n779), .B1(G159), .B2(new_n759), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n777), .A2(new_n249), .B1(new_n763), .B2(new_n337), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n773), .A2(new_n205), .B1(new_n784), .B2(new_n844), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1072), .A2(new_n1074), .A3(new_n1076), .A4(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n757), .B1(new_n1071), .B2(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n818), .A2(new_n707), .B1(new_n206), .B2(new_n709), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT114), .Z(new_n1083));
  NOR2_X1   g0883(.A1(new_n233), .A2(new_n499), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n279), .A2(G50), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT50), .ZN(new_n1086));
  AOI21_X1  g0886(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1086), .A2(new_n708), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n814), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1083), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n804), .B(new_n1081), .C1(new_n809), .C2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n701), .B2(new_n822), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1058), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1057), .A2(new_n1094), .ZN(G393));
  OAI21_X1  g0895(.A(new_n809), .B1(new_n210), .B2(new_n456), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n814), .B2(new_n244), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT115), .Z(new_n1098));
  AOI22_X1  g0898(.A1(new_n769), .A2(G311), .B1(G317), .B2(new_n759), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT52), .Z(new_n1100));
  NAND2_X1  g0900(.A1(new_n851), .A2(G283), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n785), .A2(G322), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1101), .A2(new_n775), .A3(new_n1102), .A4(new_n393), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n1103), .A2(KEYINPUT116), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1103), .A2(KEYINPUT116), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n782), .A2(new_n610), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n780), .A2(new_n603), .B1(new_n763), .B2(new_n588), .ZN(new_n1107));
  NOR4_X1   g0907(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(G159), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n768), .A2(new_n1109), .B1(new_n844), .B2(new_n760), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT51), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n811), .B1(new_n249), .B2(new_n782), .C1(new_n780), .C2(new_n202), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n777), .A2(new_n337), .B1(new_n773), .B2(new_n776), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n763), .A2(new_n279), .B1(new_n784), .B2(new_n845), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1100), .A2(new_n1108), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1098), .B(new_n754), .C1(new_n757), .C2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n808), .B2(new_n978), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n1006), .B2(new_n753), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n710), .B1(new_n1016), .B2(new_n1006), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1120), .B1(new_n1019), .B2(new_n1121), .ZN(G390));
  AND3_X1   g0922(.A1(new_n868), .A2(G330), .A3(new_n875), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT101), .B1(new_n835), .B2(new_n943), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n934), .B(new_n941), .C1(new_n680), .C2(new_n834), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n875), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n949), .A2(new_n952), .B1(new_n1126), .B2(new_n950), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n653), .A2(new_n894), .A3(new_n418), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(KEYINPUT37), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n905), .A2(new_n913), .B1(new_n1129), .B2(new_n896), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n919), .B1(new_n1130), .B2(KEYINPUT38), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n917), .A2(KEYINPUT104), .A3(new_n899), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n898), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n950), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n863), .B1(new_n724), .B2(new_n725), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n933), .B1(new_n1136), .B2(new_n943), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1123), .B1(new_n1127), .B2(new_n1138), .ZN(new_n1139));
  AND4_X1   g0939(.A1(new_n519), .A2(new_n715), .A3(new_n599), .A4(new_n524), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n718), .A2(new_n720), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n723), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(KEYINPUT90), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n941), .B1(new_n1145), .B2(new_n863), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n950), .B(new_n1134), .C1(new_n1146), .C2(new_n933), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n868), .A2(G330), .A3(new_n875), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n898), .A2(new_n909), .A3(KEYINPUT39), .ZN(new_n1149));
  AOI21_X1  g0949(.A(KEYINPUT39), .B1(new_n1133), .B2(new_n898), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n942), .A2(new_n944), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n951), .B1(new_n1152), .B2(new_n875), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1147), .B(new_n1148), .C1(new_n1151), .C2(new_n1153), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1139), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n806), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n754), .B1(new_n841), .B2(new_n1075), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n851), .A2(G150), .ZN(new_n1158));
  INV_X1    g0958(.A(G128), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1158), .A2(KEYINPUT53), .B1(new_n1159), .B2(new_n760), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT54), .B(G143), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n246), .B1(new_n763), .B2(new_n1161), .C1(new_n202), .C2(new_n773), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(G137), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n780), .A2(new_n1164), .B1(new_n782), .B2(new_n1109), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(KEYINPUT53), .B2(new_n1158), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n769), .A2(G132), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n799), .A2(G125), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1163), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n456), .A2(new_n763), .B1(new_n773), .B2(new_n337), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n780), .A2(new_n206), .B1(new_n760), .B2(new_n792), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(G77), .C2(new_n849), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n799), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1172), .B1(new_n610), .B2(new_n768), .C1(new_n588), .C2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n393), .B1(new_n777), .B2(new_n776), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT120), .Z(new_n1176));
  OAI21_X1  g0976(.A(new_n1169), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1157), .B1(new_n1177), .B2(new_n805), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1155), .A2(new_n753), .B1(new_n1156), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n445), .A2(new_n746), .A3(G330), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n955), .A2(new_n666), .A3(new_n1180), .ZN(new_n1181));
  AND4_X1   g0981(.A1(new_n744), .A2(new_n649), .A3(new_n599), .A4(new_n723), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n740), .A2(new_n689), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT31), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n740), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(G330), .B(new_n863), .C1(new_n1182), .C2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n933), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n942), .A2(new_n944), .B1(new_n1189), .B2(new_n1148), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT118), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n875), .B1(new_n868), .B2(G330), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1123), .A2(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1190), .A2(new_n1191), .B1(new_n1146), .B2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1195));
  OAI21_X1  g0995(.A(KEYINPUT118), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1181), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1139), .A2(new_n1197), .A3(new_n1154), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1198), .A2(KEYINPUT119), .A3(new_n710), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n1155), .B2(new_n1197), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT119), .B1(new_n1198), .B2(new_n710), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1179), .B1(new_n1200), .B2(new_n1201), .ZN(G378));
  INV_X1    g1002(.A(new_n1181), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1198), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(G330), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n903), .A2(new_n908), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1206), .A2(KEYINPUT38), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT40), .B1(new_n1207), .B2(new_n911), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n910), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1205), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n954), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n292), .A2(new_n881), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n308), .B(new_n1212), .Z(new_n1213));
  XNOR2_X1  g1013(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1213), .B(new_n1214), .Z(new_n1215));
  OAI211_X1 g1015(.A(new_n953), .B(new_n947), .C1(new_n924), .C2(new_n1205), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1211), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1215), .B1(new_n1211), .B2(new_n1216), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1204), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT57), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n711), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1204), .B(KEYINPUT57), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT122), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1211), .A2(new_n1216), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1215), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1211), .A2(new_n1216), .A3(new_n1215), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1229), .A2(KEYINPUT122), .A3(KEYINPUT57), .A4(new_n1204), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1221), .A2(new_n1224), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1215), .A2(new_n806), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n754), .B1(new_n841), .B2(G50), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n494), .B1(new_n777), .B2(new_n249), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n375), .A2(new_n763), .B1(new_n773), .B2(new_n960), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1234), .B(new_n1235), .C1(new_n769), .C2(G107), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n792), .B2(new_n1173), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n780), .A2(new_n205), .B1(new_n760), .B2(new_n610), .ZN(new_n1238));
  NOR4_X1   g1038(.A1(new_n1237), .A2(new_n811), .A3(new_n1041), .A4(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n494), .B1(new_n812), .B2(new_n276), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1239), .A2(KEYINPUT58), .B1(new_n202), .B2(new_n1240), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n777), .A2(new_n1161), .B1(new_n763), .B2(new_n1164), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G132), .B2(new_n779), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n849), .A2(G150), .B1(G125), .B2(new_n759), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1243), .B(new_n1244), .C1(new_n1159), .C2(new_n768), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1245), .A2(KEYINPUT59), .ZN(new_n1246));
  AOI211_X1 g1046(.A(G33), .B(G41), .C1(new_n774), .C2(G159), .ZN(new_n1247));
  INV_X1    g1047(.A(G124), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1247), .B1(new_n1248), .B2(new_n784), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT121), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1245), .A2(KEYINPUT59), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1241), .B1(KEYINPUT58), .B2(new_n1239), .C1(new_n1246), .C2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1233), .B1(new_n1253), .B2(new_n805), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1229), .A2(new_n753), .B1(new_n1232), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1231), .A2(new_n1255), .ZN(G375));
  NAND2_X1  g1056(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n753), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n841), .A2(G68), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n777), .A2(new_n205), .B1(new_n763), .B2(new_n206), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n246), .B(new_n1260), .C1(G77), .C2(new_n774), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n1261), .B1(new_n792), .B2(new_n768), .C1(new_n603), .C2(new_n1173), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n1073), .B1(new_n760), .B2(new_n588), .C1(new_n610), .C2(new_n780), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n812), .B1(G132), .B2(new_n759), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n1264), .B1(new_n202), .B2(new_n782), .C1(new_n780), .C2(new_n1161), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n777), .A2(new_n1109), .B1(new_n773), .B2(new_n960), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(G150), .B2(new_n790), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n1267), .B1(new_n1164), .B2(new_n768), .C1(new_n1173), .C2(new_n1159), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n1262), .A2(new_n1263), .B1(new_n1265), .B2(new_n1268), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n804), .B(new_n1259), .C1(new_n1269), .C2(new_n805), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n875), .B2(new_n807), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1258), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1197), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1194), .A2(new_n1181), .A3(new_n1196), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n1000), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1273), .A2(new_n1276), .ZN(G381));
  NOR3_X1   g1077(.A1(new_n1056), .A2(G396), .A3(new_n1093), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n865), .ZN(new_n1279));
  XOR2_X1   g1079(.A(new_n1279), .B(KEYINPUT123), .Z(new_n1280));
  OR4_X1    g1080(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G378), .A2(KEYINPUT124), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT124), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1179), .B(new_n1283), .C1(new_n1200), .C2(new_n1201), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(new_n1255), .A3(new_n1231), .ZN(new_n1286));
  OR2_X1    g1086(.A1(new_n1281), .A2(new_n1286), .ZN(G407));
  NAND2_X1  g1087(.A1(new_n688), .A2(G213), .ZN(new_n1288));
  OR2_X1    g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G213), .B(new_n1289), .C1(new_n1281), .C2(new_n1286), .ZN(G409));
  AOI21_X1  g1090(.A(new_n824), .B1(new_n1057), .B2(new_n1094), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1291), .A2(new_n1278), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(G390), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(G390), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1053), .A2(new_n1293), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1293), .ZN(new_n1297));
  OAI22_X1  g1097(.A1(new_n1297), .A2(new_n1294), .B1(new_n1022), .B2(new_n1052), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT61), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1288), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(G2897), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT60), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1275), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1274), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT126), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT126), .B1(new_n1304), .B2(new_n1274), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n710), .B1(new_n1275), .B2(new_n1303), .ZN(new_n1309));
  NOR3_X1   g1109(.A1(new_n1307), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n865), .B1(new_n1310), .B2(new_n1272), .ZN(new_n1311));
  OR2_X1    g1111(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1312));
  OAI211_X1 g1112(.A(G384), .B(new_n1273), .C1(new_n1312), .C2(new_n1307), .ZN(new_n1313));
  AOI211_X1 g1113(.A(KEYINPUT127), .B(new_n1302), .C1(new_n1311), .C2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT127), .ZN(new_n1316));
  OAI211_X1 g1116(.A(G2897), .B(new_n1301), .C1(new_n1315), .C2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1314), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1255), .B1(new_n999), .B2(new_n1219), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1282), .A2(new_n1320), .A3(new_n1284), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1231), .A2(G378), .A3(new_n1255), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT125), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1231), .A2(KEYINPUT125), .A3(G378), .A4(new_n1255), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1321), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1319), .B1(new_n1326), .B2(new_n1301), .ZN(new_n1327));
  NOR3_X1   g1127(.A1(new_n1326), .A2(new_n1301), .A3(new_n1315), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT62), .ZN(new_n1329));
  OAI211_X1 g1129(.A(new_n1300), .B(new_n1327), .C1(new_n1328), .C2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1321), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1315), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1333), .A2(new_n1288), .A3(new_n1334), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1335), .A2(KEYINPUT62), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1299), .B1(new_n1330), .B2(new_n1336), .ZN(new_n1337));
  AND2_X1   g1137(.A1(new_n1327), .A2(new_n1300), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1299), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT63), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1335), .A2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1328), .A2(KEYINPUT63), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1338), .A2(new_n1339), .A3(new_n1341), .A4(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1337), .A2(new_n1343), .ZN(G405));
  NAND2_X1  g1144(.A1(new_n1285), .A2(G375), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1331), .A2(new_n1345), .ZN(new_n1346));
  XNOR2_X1  g1146(.A(new_n1346), .B(new_n1334), .ZN(new_n1347));
  XNOR2_X1  g1147(.A(new_n1347), .B(new_n1299), .ZN(G402));
endmodule


