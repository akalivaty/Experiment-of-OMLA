//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024;
  INV_X1    g000(.A(G1gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT16), .ZN(new_n203));
  INV_X1    g002(.A(G15gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(G22gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G15gat), .ZN(new_n207));
  AND3_X1   g006(.A1(new_n203), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(G1gat), .B1(new_n205), .B2(new_n207), .ZN(new_n209));
  OAI21_X1  g008(.A(G8gat), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n203), .A2(new_n205), .A3(new_n207), .ZN(new_n211));
  INV_X1    g010(.A(G8gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(G15gat), .B(G22gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n211), .B(new_n212), .C1(G1gat), .C2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT86), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n210), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n215), .B1(new_n210), .B2(new_n214), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G43gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G50gat), .ZN(new_n220));
  INV_X1    g019(.A(G50gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G43gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n222), .A3(KEYINPUT15), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(KEYINPUT85), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT85), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G50gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n226), .A3(new_n219), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT15), .B1(new_n227), .B2(new_n222), .ZN(new_n228));
  INV_X1    g027(.A(G29gat), .ZN(new_n229));
  INV_X1    g028(.A(G36gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(new_n230), .A3(KEYINPUT14), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT14), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G29gat), .B2(G36gat), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n231), .B(new_n233), .C1(new_n229), .C2(new_n230), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n223), .B1(new_n228), .B2(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n234), .A2(new_n223), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT17), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT17), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n235), .A2(new_n239), .A3(new_n236), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n218), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n210), .A2(new_n214), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n237), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G229gat), .A2(G233gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n241), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT18), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n237), .B(new_n243), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n246), .B(KEYINPUT13), .Z(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n241), .A2(KEYINPUT18), .A3(new_n245), .A4(new_n246), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n249), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G141gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G169gat), .B(G197gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(new_n259), .B(KEYINPUT12), .Z(new_n260));
  NAND2_X1  g059(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n260), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n262), .A2(new_n249), .A3(new_n252), .A4(new_n253), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n261), .A2(KEYINPUT87), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT87), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n254), .A2(new_n265), .A3(new_n260), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G78gat), .B(G106gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT31), .B(G50gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  AND2_X1   g069(.A1(G228gat), .A2(G233gat), .ZN(new_n271));
  XOR2_X1   g070(.A(G141gat), .B(G148gat), .Z(new_n272));
  INV_X1    g071(.A(G155gat), .ZN(new_n273));
  INV_X1    g072(.A(G162gat), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT2), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G155gat), .B(G162gat), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT3), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n272), .A2(new_n277), .A3(new_n275), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT29), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n285));
  OR2_X1    g084(.A1(G197gat), .A2(G204gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(G197gat), .A2(G204gat), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(G211gat), .B(G218gat), .Z(new_n289));
  OR3_X1    g088(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT73), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n288), .B2(KEYINPUT73), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n284), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n292), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT3), .B1(new_n294), .B2(new_n283), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n279), .A2(new_n281), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n271), .B(new_n293), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n289), .A2(KEYINPUT77), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n298), .A2(new_n288), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n289), .A2(KEYINPUT77), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(new_n288), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n283), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT78), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n299), .A2(KEYINPUT78), .A3(new_n283), .A4(new_n301), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n305), .A3(new_n280), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n279), .A2(new_n281), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n306), .A2(new_n307), .B1(new_n292), .B2(new_n284), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n206), .B(new_n297), .C1(new_n308), .C2(new_n271), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n270), .B1(new_n310), .B2(KEYINPUT79), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n297), .B1(new_n308), .B2(new_n271), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G22gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n309), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n313), .A2(KEYINPUT79), .A3(new_n309), .A4(new_n270), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT66), .ZN(new_n319));
  NAND2_X1  g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G183gat), .A2(G190gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT24), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n322), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n329), .B1(G169gat), .B2(G176gat), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n325), .A2(new_n328), .A3(KEYINPUT25), .A4(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT23), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n319), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n330), .B(new_n320), .C1(KEYINPUT24), .C2(new_n322), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n323), .A2(new_n326), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n338), .A2(KEYINPUT66), .A3(KEYINPUT25), .A4(new_n333), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT64), .B(G169gat), .ZN(new_n341));
  INV_X1    g140(.A(G176gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(KEYINPUT23), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT65), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT65), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n341), .A2(new_n345), .A3(KEYINPUT23), .A4(new_n342), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n338), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT25), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n340), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT27), .B(G183gat), .ZN(new_n351));
  INV_X1    g150(.A(G190gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  XOR2_X1   g152(.A(new_n353), .B(KEYINPUT28), .Z(new_n354));
  INV_X1    g153(.A(KEYINPUT26), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n321), .B1(new_n355), .B2(new_n332), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n356), .B1(new_n355), .B2(new_n332), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(new_n322), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n350), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT67), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n340), .A2(new_n362), .A3(new_n349), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n362), .B1(new_n340), .B2(new_n349), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n358), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n294), .B(new_n361), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n359), .A2(new_n366), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(new_n365), .B2(new_n360), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n367), .B1(new_n369), .B2(new_n294), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT30), .ZN(new_n371));
  XNOR2_X1  g170(.A(G64gat), .B(G92gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(G36gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(KEYINPUT74), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(new_n212), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n370), .A2(new_n371), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n370), .A2(new_n376), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n367), .B(new_n375), .C1(new_n369), .C2(new_n294), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(KEYINPUT30), .A3(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT0), .B(G57gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(G85gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(G1gat), .B(G29gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  XOR2_X1   g183(.A(G127gat), .B(G134gat), .Z(new_n385));
  XOR2_X1   g184(.A(G113gat), .B(G120gat), .Z(new_n386));
  AOI21_X1  g185(.A(new_n385), .B1(KEYINPUT68), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT1), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n388), .B(new_n386), .C1(new_n385), .C2(KEYINPUT68), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n296), .ZN(new_n393));
  NAND2_X1  g192(.A1(G225gat), .A2(G233gat), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n280), .B1(new_n279), .B2(new_n281), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n398), .A2(new_n391), .A3(new_n390), .A4(new_n282), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n392), .A2(new_n296), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n400), .B1(new_n392), .B2(new_n296), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n396), .B(new_n399), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT5), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n307), .A2(new_n391), .A3(new_n390), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n393), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n407), .B2(new_n395), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n393), .A2(KEYINPUT4), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n392), .A2(new_n397), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n410), .A2(new_n401), .B1(new_n282), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n395), .A2(KEYINPUT5), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n384), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT76), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT6), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n416), .B1(new_n415), .B2(KEYINPUT6), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n409), .A2(new_n414), .ZN(new_n420));
  INV_X1    g219(.A(new_n384), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT75), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n404), .A2(new_n408), .B1(new_n412), .B2(new_n413), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT6), .B1(new_n424), .B2(new_n384), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT75), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n415), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n423), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n377), .A2(new_n380), .B1(new_n419), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n318), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n425), .A2(new_n422), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n419), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n292), .B(new_n361), .C1(new_n365), .C2(new_n366), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n433), .A2(KEYINPUT81), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(KEYINPUT81), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n434), .B(new_n435), .C1(new_n292), .C2(new_n369), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT38), .B1(new_n436), .B2(KEYINPUT37), .ZN(new_n437));
  XOR2_X1   g236(.A(KEYINPUT82), .B(KEYINPUT37), .Z(new_n438));
  AOI21_X1  g237(.A(new_n376), .B1(new_n370), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n432), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT37), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n439), .B1(new_n441), .B2(new_n370), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n442), .A2(KEYINPUT38), .B1(new_n370), .B2(new_n376), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n380), .A2(new_n377), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT80), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT39), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n407), .A2(new_n395), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n399), .B1(new_n402), .B2(new_n403), .ZN(new_n448));
  AOI211_X1 g247(.A(new_n446), .B(new_n447), .C1(new_n448), .C2(new_n395), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n446), .A3(new_n395), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n384), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n445), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n452), .A2(KEYINPUT40), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n444), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n415), .B1(new_n452), .B2(KEYINPUT40), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n440), .A2(new_n443), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n430), .B1(new_n456), .B2(new_n318), .ZN(new_n457));
  XNOR2_X1  g256(.A(G15gat), .B(G43gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(G71gat), .B(G99gat), .ZN(new_n459));
  XOR2_X1   g258(.A(new_n458), .B(new_n459), .Z(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT69), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n392), .B(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n463), .B(new_n358), .C1(new_n363), .C2(new_n364), .ZN(new_n464));
  NAND2_X1  g263(.A1(G227gat), .A2(G233gat), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n358), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n350), .A2(KEYINPUT67), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n340), .A2(new_n362), .A3(new_n349), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n392), .A2(KEYINPUT69), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n464), .B(new_n466), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT70), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n365), .A2(KEYINPUT69), .A3(new_n392), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT70), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n474), .A2(new_n475), .A3(new_n466), .A4(new_n464), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT33), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n461), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n477), .A2(KEYINPUT32), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT34), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT71), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n483), .B1(new_n465), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n482), .A2(new_n465), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n486), .B1(new_n482), .B2(new_n465), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n481), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n482), .A2(new_n465), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n485), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n482), .A2(new_n465), .A3(new_n486), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT32), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(new_n473), .B2(new_n476), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n480), .B1(new_n490), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n489), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n494), .A2(new_n496), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n479), .A3(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n498), .A2(KEYINPUT72), .A3(new_n499), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n499), .A2(KEYINPUT72), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n499), .A2(KEYINPUT72), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n500), .A2(new_n479), .A3(new_n501), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n479), .B1(new_n500), .B2(new_n501), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n504), .B(new_n505), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n457), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n506), .A2(new_n507), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT83), .B(KEYINPUT35), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n432), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n510), .A2(new_n317), .A3(new_n444), .A4(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n498), .A2(new_n429), .A3(new_n502), .A4(new_n317), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT35), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n267), .B1(new_n509), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G71gat), .B(G78gat), .ZN(new_n519));
  INV_X1    g318(.A(G57gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(G64gat), .ZN(new_n521));
  INV_X1    g320(.A(G64gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(G57gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT88), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n524), .B1(new_n521), .B2(new_n523), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT9), .ZN(new_n528));
  INV_X1    g327(.A(G71gat), .ZN(new_n529));
  INV_X1    g328(.A(G78gat), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n519), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n519), .A2(new_n531), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n522), .A2(KEYINPUT89), .A3(G57gat), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT89), .B1(new_n522), .B2(G57gat), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n521), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT21), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n243), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(G183gat), .ZN(new_n542));
  INV_X1    g341(.A(G183gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n540), .A2(new_n243), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n545), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n543), .B1(new_n540), .B2(new_n243), .ZN(new_n548));
  AOI211_X1 g347(.A(G183gat), .B(new_n242), .C1(new_n539), .C2(KEYINPUT21), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G127gat), .B(G155gat), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n552), .B(G211gat), .Z(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n539), .A2(KEYINPUT21), .ZN(new_n555));
  NAND2_X1  g354(.A1(G231gat), .A2(G233gat), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n556), .B(KEYINPUT90), .Z(new_n557));
  XNOR2_X1  g356(.A(new_n555), .B(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n553), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n546), .A2(new_n550), .A3(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n554), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n558), .B1(new_n554), .B2(new_n560), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G134gat), .B(G162gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  INV_X1    g367(.A(G92gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(KEYINPUT8), .A2(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT7), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(new_n568), .B2(new_n569), .ZN(new_n572));
  NAND3_X1  g371(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(new_n567), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n567), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n570), .A2(new_n577), .A3(new_n572), .A4(new_n573), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT92), .ZN(new_n580));
  XOR2_X1   g379(.A(G190gat), .B(G218gat), .Z(new_n581));
  OAI22_X1  g380(.A1(new_n237), .A2(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n235), .A2(new_n239), .A3(new_n236), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n239), .B1(new_n235), .B2(new_n236), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT91), .B1(new_n586), .B2(new_n579), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n238), .A2(KEYINPUT91), .A3(new_n240), .A4(new_n579), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n566), .B(new_n583), .C1(new_n587), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT93), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n581), .A2(new_n580), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n592), .B(new_n593), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n238), .A2(new_n240), .A3(new_n579), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT91), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n582), .B1(new_n598), .B2(new_n588), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT93), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(new_n566), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n591), .A2(new_n595), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n595), .B1(new_n591), .B2(new_n601), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n565), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n598), .A2(new_n588), .ZN(new_n605));
  AND4_X1   g404(.A1(new_n600), .A2(new_n605), .A3(new_n566), .A4(new_n583), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n600), .B1(new_n599), .B2(new_n566), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n594), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n595), .A3(new_n601), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n608), .A2(new_n564), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n563), .A2(new_n604), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT94), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT94), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n563), .A2(new_n604), .A3(new_n614), .A4(new_n610), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(G230gat), .ZN(new_n617));
  INV_X1    g416(.A(G233gat), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n579), .B1(new_n532), .B2(new_n538), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT10), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n521), .A2(new_n523), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT88), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(new_n531), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n519), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n627), .A2(new_n537), .A3(new_n578), .A4(new_n576), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n620), .A2(new_n621), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n579), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n539), .A2(KEYINPUT10), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n619), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n620), .A2(new_n628), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n619), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(G204gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT95), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(new_n342), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n633), .A2(new_n635), .A3(new_n640), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n613), .A2(new_n616), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n518), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT96), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n518), .A2(KEYINPUT96), .A3(new_n645), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n419), .A2(new_n428), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g453(.A(KEYINPUT16), .B(G8gat), .Z(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  AOI211_X1 g455(.A(new_n444), .B(new_n656), .C1(new_n648), .C2(new_n649), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT42), .B1(new_n657), .B2(KEYINPUT97), .ZN(new_n658));
  INV_X1    g457(.A(new_n444), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n650), .A2(new_n659), .A3(new_n655), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT97), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n650), .ZN(new_n664));
  OAI21_X1  g463(.A(G8gat), .B1(new_n664), .B2(new_n444), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n658), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT98), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n658), .A2(new_n663), .A3(KEYINPUT98), .A4(new_n665), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(G1325gat));
  AOI21_X1  g469(.A(G15gat), .B1(new_n650), .B2(new_n510), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n508), .A2(new_n503), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT99), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n508), .A2(KEYINPUT99), .A3(new_n503), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n664), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n671), .B1(new_n677), .B2(G15gat), .ZN(G1326gat));
  NAND2_X1  g477(.A1(new_n650), .A2(new_n318), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n608), .A2(new_n564), .A3(new_n609), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n564), .B1(new_n608), .B2(new_n609), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI211_X1 g484(.A(new_n682), .B(new_n685), .C1(new_n509), .C2(new_n517), .ZN(new_n686));
  INV_X1    g485(.A(new_n685), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n514), .A2(new_n688), .A3(new_n516), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n688), .B1(new_n514), .B2(new_n516), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n674), .A2(new_n457), .A3(new_n675), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n687), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n686), .B1(new_n694), .B2(new_n682), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n264), .A2(KEYINPUT100), .A3(new_n266), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT100), .B1(new_n264), .B2(new_n266), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n563), .A2(new_n644), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n695), .A2(new_n696), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n509), .A2(new_n517), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n703), .A2(KEYINPUT44), .A3(new_n687), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n515), .A2(KEYINPUT35), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n498), .A2(new_n502), .A3(new_n317), .A4(new_n444), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n512), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT101), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n689), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n674), .A2(new_n457), .A3(new_n675), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n685), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n701), .B(new_n704), .C1(new_n711), .C2(KEYINPUT44), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT102), .B1(new_n712), .B2(new_n699), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n702), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(G29gat), .B1(new_n715), .B2(new_n651), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n685), .A2(new_n563), .A3(new_n644), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n518), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(new_n229), .A3(new_n652), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT45), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n716), .A2(new_n721), .ZN(G1328gat));
  OAI21_X1  g521(.A(G36gat), .B1(new_n715), .B2(new_n444), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n718), .A2(G36gat), .A3(new_n444), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT46), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(G1329gat));
  NAND3_X1  g525(.A1(new_n695), .A2(new_n700), .A3(new_n701), .ZN(new_n727));
  OAI21_X1  g526(.A(G43gat), .B1(new_n727), .B2(new_n676), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n719), .A2(new_n219), .A3(new_n510), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n728), .A2(KEYINPUT47), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT103), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT103), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n728), .A2(new_n732), .A3(KEYINPUT47), .A4(new_n729), .ZN(new_n733));
  INV_X1    g532(.A(new_n729), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n674), .A2(new_n675), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n714), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n734), .B1(new_n736), .B2(G43gat), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n731), .B(new_n733), .C1(new_n737), .C2(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g537(.A1(new_n224), .A2(new_n226), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(new_n727), .B2(new_n317), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n719), .A2(new_n318), .A3(new_n739), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n741), .A2(KEYINPUT48), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT104), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n741), .A2(new_n745), .A3(KEYINPUT48), .A4(new_n742), .ZN(new_n746));
  INV_X1    g545(.A(new_n742), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n714), .A2(new_n318), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n740), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n744), .B(new_n746), .C1(new_n749), .C2(KEYINPUT48), .ZN(G1331gat));
  AOI211_X1 g549(.A(new_n613), .B(new_n616), .C1(new_n709), .C2(new_n710), .ZN(new_n751));
  INV_X1    g550(.A(new_n644), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n700), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n651), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(new_n520), .ZN(G1332gat));
  NOR2_X1   g555(.A1(new_n754), .A2(new_n444), .ZN(new_n757));
  NOR2_X1   g556(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n758));
  AND2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n757), .B2(new_n758), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n754), .B2(new_n676), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n751), .A2(new_n529), .A3(new_n510), .A4(new_n753), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n763), .B1(new_n762), .B2(new_n764), .ZN(new_n768));
  OR3_X1    g567(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n766), .B2(new_n768), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1334gat));
  NOR2_X1   g570(.A1(new_n754), .A2(new_n317), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(new_n530), .ZN(G1335gat));
  INV_X1    g572(.A(new_n563), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n695), .A2(new_n774), .A3(new_n753), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n775), .A2(new_n568), .A3(new_n651), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n711), .A2(new_n774), .A3(new_n699), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n644), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n781), .A2(new_n651), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n776), .B1(new_n782), .B2(new_n568), .ZN(G1336gat));
  INV_X1    g582(.A(new_n775), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n569), .B1(new_n784), .B2(new_n659), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n777), .A2(KEYINPUT106), .A3(KEYINPUT51), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT51), .B1(new_n777), .B2(KEYINPUT106), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n444), .A2(G92gat), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NOR4_X1   g588(.A1(new_n786), .A2(new_n787), .A3(new_n752), .A4(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT52), .B1(new_n785), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n781), .B2(new_n789), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n785), .B2(new_n793), .ZN(G1337gat));
  OAI21_X1  g593(.A(G99gat), .B1(new_n775), .B2(new_n676), .ZN(new_n795));
  INV_X1    g594(.A(new_n510), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n796), .A2(G99gat), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n795), .B1(new_n781), .B2(new_n797), .ZN(G1338gat));
  NAND4_X1  g597(.A1(new_n695), .A2(new_n318), .A3(new_n774), .A4(new_n753), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n799), .A2(G106gat), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n317), .A2(G106gat), .A3(new_n752), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n786), .A2(new_n787), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT53), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT53), .B1(new_n799), .B2(G106gat), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n801), .B1(new_n779), .B2(new_n780), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n805), .A2(KEYINPUT107), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT107), .B1(new_n805), .B2(new_n806), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(G1339gat));
  NAND2_X1  g608(.A1(new_n629), .A2(new_n631), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  INV_X1    g610(.A(new_n619), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n629), .A2(new_n631), .A3(new_n619), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT54), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n641), .B(new_n813), .C1(new_n815), .C2(new_n632), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n643), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n633), .A2(KEYINPUT54), .A3(new_n814), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n640), .B1(new_n632), .B2(new_n811), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT55), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT108), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n816), .A2(new_n817), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n819), .A2(new_n820), .A3(KEYINPUT55), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT108), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n823), .A2(new_n824), .A3(new_n825), .A4(new_n643), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT100), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n267), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n264), .A2(KEYINPUT100), .A3(new_n266), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n827), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n246), .B1(new_n241), .B2(new_n245), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n250), .A2(new_n251), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n259), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n263), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n752), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT110), .B1(new_n831), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT110), .ZN(new_n838));
  INV_X1    g637(.A(new_n836), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n838), .B(new_n839), .C1(new_n699), .C2(new_n827), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n837), .A2(new_n685), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n835), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n842), .B1(new_n683), .B2(new_n684), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT109), .B1(new_n843), .B2(new_n827), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n835), .B1(new_n604), .B2(new_n610), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT109), .ZN(new_n846));
  INV_X1    g645(.A(new_n827), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n563), .B1(new_n841), .B2(new_n849), .ZN(new_n850));
  AND4_X1   g649(.A1(new_n612), .A2(new_n615), .A3(new_n752), .A4(new_n699), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(new_n318), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT111), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n796), .A2(new_n659), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(new_n652), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(G113gat), .B1(new_n857), .B2(new_n267), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n853), .A2(new_n510), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n659), .A2(new_n651), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n863), .A2(G113gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n858), .B1(new_n699), .B2(new_n864), .ZN(G1340gat));
  OAI21_X1  g664(.A(G120gat), .B1(new_n857), .B2(new_n752), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n863), .A2(G120gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n752), .B2(new_n867), .ZN(G1341gat));
  AOI21_X1  g667(.A(G127gat), .B1(new_n862), .B2(new_n563), .ZN(new_n869));
  INV_X1    g668(.A(G127gat), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n857), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n869), .B1(new_n871), .B2(new_n563), .ZN(G1342gat));
  OAI21_X1  g671(.A(G134gat), .B1(new_n857), .B2(new_n685), .ZN(new_n873));
  INV_X1    g672(.A(G134gat), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n862), .A2(new_n874), .A3(new_n687), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n875), .A2(KEYINPUT56), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(KEYINPUT56), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n873), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT112), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n873), .A2(new_n876), .A3(KEYINPUT112), .A4(new_n877), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1343gat));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n735), .A2(new_n861), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n841), .A2(new_n849), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n774), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n612), .A2(new_n615), .A3(new_n752), .A4(new_n699), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n884), .A2(new_n888), .A3(new_n318), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n889), .A2(G141gat), .A3(new_n267), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n890), .B(new_n891), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n823), .A2(KEYINPUT113), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n823), .A2(KEYINPUT113), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n893), .A2(new_n266), .A3(new_n264), .A4(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n839), .B1(new_n895), .B2(new_n818), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n685), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n843), .A2(KEYINPUT109), .A3(new_n827), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n846), .B1(new_n845), .B2(new_n847), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n851), .B1(new_n900), .B2(new_n774), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT114), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n317), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n901), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  AOI22_X1  g705(.A1(new_n844), .A2(new_n848), .B1(new_n685), .B2(new_n896), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n887), .B1(new_n907), .B2(new_n563), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT114), .B1(new_n908), .B2(new_n904), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n318), .B1(new_n850), .B2(new_n851), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n903), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n267), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(new_n914), .A3(new_n884), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT58), .B1(new_n915), .B2(G141gat), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n883), .B1(new_n892), .B2(new_n916), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n892), .A2(new_n883), .A3(new_n916), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT57), .B1(new_n888), .B2(new_n318), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n902), .B1(new_n901), .B2(new_n905), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n908), .A2(KEYINPUT114), .A3(new_n904), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n884), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT115), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n913), .A2(KEYINPUT115), .A3(new_n884), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n700), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n890), .B1(new_n928), .B2(G141gat), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT58), .ZN(new_n930));
  OAI22_X1  g729(.A1(new_n917), .A2(new_n918), .B1(new_n929), .B2(new_n930), .ZN(G1344gat));
  AOI21_X1  g730(.A(new_n752), .B1(new_n925), .B2(new_n926), .ZN(new_n932));
  INV_X1    g731(.A(G148gat), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n933), .A2(KEYINPUT59), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n932), .A2(KEYINPUT118), .A3(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT118), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT115), .B1(new_n913), .B2(new_n884), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n676), .A2(new_n860), .ZN(new_n939));
  AOI211_X1 g738(.A(new_n924), .B(new_n939), .C1(new_n910), .C2(new_n912), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n644), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n937), .B1(new_n941), .B2(new_n934), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT119), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n888), .A2(new_n943), .A3(new_n904), .ZN(new_n944));
  OAI21_X1  g743(.A(KEYINPUT119), .B1(new_n852), .B2(new_n905), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n645), .A2(new_n267), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n845), .A2(new_n643), .A3(new_n824), .A4(new_n823), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n563), .B1(new_n897), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n318), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(new_n903), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n944), .A2(new_n945), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(new_n644), .A3(new_n884), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G148gat), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT120), .B1(new_n953), .B2(KEYINPUT59), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT120), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT59), .ZN(new_n956));
  AOI211_X1 g755(.A(new_n955), .B(new_n956), .C1(new_n952), .C2(G148gat), .ZN(new_n957));
  OAI22_X1  g756(.A1(new_n936), .A2(new_n942), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n889), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n959), .A2(new_n933), .A3(new_n644), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(G1345gat));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n563), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT121), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n563), .A2(G155gat), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT122), .ZN(new_n965));
  AOI22_X1  g764(.A1(new_n963), .A2(new_n273), .B1(new_n927), .B2(new_n965), .ZN(G1346gat));
  AOI21_X1  g765(.A(G162gat), .B1(new_n959), .B2(new_n687), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n685), .B1(new_n925), .B2(new_n926), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n967), .B1(new_n968), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g768(.A1(new_n652), .A2(new_n444), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n855), .A2(new_n510), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g770(.A(G169gat), .B1(new_n971), .B2(new_n267), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n859), .A2(new_n652), .A3(new_n444), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n973), .A2(new_n341), .A3(new_n700), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n974), .ZN(G1348gat));
  AOI21_X1  g774(.A(G176gat), .B1(new_n973), .B2(new_n644), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n971), .A2(new_n752), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n976), .B1(new_n977), .B2(G176gat), .ZN(G1349gat));
  OAI21_X1  g777(.A(G183gat), .B1(new_n971), .B2(new_n774), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT123), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n563), .A2(new_n351), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n980), .B1(new_n973), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(KEYINPUT60), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT60), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n979), .A2(new_n985), .A3(new_n982), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n984), .A2(new_n986), .ZN(G1350gat));
  NAND3_X1  g786(.A1(new_n973), .A2(new_n352), .A3(new_n687), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n855), .A2(new_n510), .A3(new_n687), .A4(new_n970), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT61), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n989), .A2(new_n990), .A3(G190gat), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n990), .B1(new_n989), .B2(G190gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(G1351gat));
  XOR2_X1   g792(.A(KEYINPUT124), .B(G197gat), .Z(new_n994));
  NOR4_X1   g793(.A1(new_n735), .A2(KEYINPUT125), .A3(new_n652), .A4(new_n444), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT125), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n996), .B1(new_n676), .B2(new_n970), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n951), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n994), .B1(new_n999), .B2(new_n267), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n676), .A2(new_n970), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n1001), .A2(new_n911), .ZN(new_n1002));
  INV_X1    g801(.A(new_n1002), .ZN(new_n1003));
  OR2_X1    g802(.A1(new_n699), .A2(new_n994), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1000), .B1(new_n1003), .B2(new_n1004), .ZN(G1352gat));
  NAND3_X1  g804(.A1(new_n951), .A2(new_n998), .A3(new_n644), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1006), .A2(KEYINPUT126), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT126), .ZN(new_n1008));
  NAND4_X1  g807(.A1(new_n951), .A2(new_n998), .A3(new_n1008), .A4(new_n644), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n1007), .A2(G204gat), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g809(.A(G204gat), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n1002), .A2(new_n1011), .A3(new_n644), .ZN(new_n1012));
  XOR2_X1   g811(.A(new_n1012), .B(KEYINPUT62), .Z(new_n1013));
  NAND2_X1  g812(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1015));
  XNOR2_X1  g814(.A(new_n1014), .B(new_n1015), .ZN(G1353gat));
  OR3_X1    g815(.A1(new_n1003), .A2(G211gat), .A3(new_n774), .ZN(new_n1017));
  OAI21_X1  g816(.A(G211gat), .B1(new_n999), .B2(new_n774), .ZN(new_n1018));
  INV_X1    g817(.A(KEYINPUT63), .ZN(new_n1019));
  AND2_X1   g818(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1021));
  OAI21_X1  g820(.A(new_n1017), .B1(new_n1020), .B2(new_n1021), .ZN(G1354gat));
  OAI21_X1  g821(.A(G218gat), .B1(new_n999), .B2(new_n685), .ZN(new_n1023));
  OR2_X1    g822(.A1(new_n685), .A2(G218gat), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1023), .B1(new_n1003), .B2(new_n1024), .ZN(G1355gat));
endmodule


