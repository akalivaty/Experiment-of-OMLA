//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989;
  INV_X1    g000(.A(KEYINPUT96), .ZN(new_n202));
  NAND2_X1  g001(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(G1gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT92), .ZN(new_n206));
  INV_X1    g005(.A(G1gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n206), .B1(KEYINPUT16), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n209));
  NOR3_X1   g008(.A1(new_n209), .A2(KEYINPUT92), .A3(G1gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n204), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT95), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G8gat), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n205), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT93), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n204), .A2(G1gat), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n216), .A2(new_n211), .B1(new_n217), .B2(KEYINPUT94), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n211), .A2(new_n216), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n214), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n202), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n205), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n211), .B(KEYINPUT95), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(G8gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n218), .A2(new_n219), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G8gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n226), .A3(KEYINPUT96), .ZN(new_n227));
  XOR2_X1   g026(.A(G43gat), .B(G50gat), .Z(new_n228));
  XOR2_X1   g027(.A(KEYINPUT91), .B(KEYINPUT15), .Z(new_n229));
  OR3_X1    g028(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n228), .A2(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT15), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G36gat), .ZN(new_n235));
  XOR2_X1   g034(.A(KEYINPUT90), .B(G29gat), .Z(new_n236));
  OAI211_X1 g035(.A(new_n232), .B(new_n234), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n235), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT89), .ZN(new_n239));
  OR2_X1    g038(.A1(new_n230), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n231), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n241), .B1(new_n230), .B2(new_n239), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n238), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n237), .B1(new_n243), .B2(new_n234), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n221), .A2(new_n227), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G229gat), .A2(G233gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT17), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n237), .B(KEYINPUT17), .C1(new_n243), .C2(new_n234), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n248), .A2(new_n226), .A3(new_n224), .A4(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n245), .A2(new_n246), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT18), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT97), .ZN(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G141gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G169gat), .B(G197gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(new_n259), .B(KEYINPUT12), .Z(new_n260));
  NAND2_X1  g059(.A1(new_n221), .A2(new_n227), .ZN(new_n261));
  INV_X1    g060(.A(new_n244), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n245), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n246), .B(KEYINPUT13), .Z(new_n265));
  AOI21_X1  g064(.A(new_n260), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n245), .A2(KEYINPUT18), .A3(new_n246), .A4(new_n250), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT97), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n268), .A3(new_n252), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n254), .A2(new_n266), .A3(new_n267), .A4(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n245), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n244), .B1(new_n221), .B2(new_n227), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n265), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n253), .A2(new_n273), .A3(new_n267), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(new_n260), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(G8gat), .B(G36gat), .Z(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT79), .ZN(new_n279));
  XNOR2_X1  g078(.A(G64gat), .B(G92gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  XNOR2_X1  g080(.A(G197gat), .B(G204gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT22), .ZN(new_n283));
  INV_X1    g082(.A(G211gat), .ZN(new_n284));
  INV_X1    g083(.A(G218gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G211gat), .B(G218gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G169gat), .ZN(new_n290));
  INV_X1    g089(.A(G176gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT23), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT23), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(G169gat), .B2(G176gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n292), .A2(new_n294), .A3(KEYINPUT25), .A4(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G183gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT64), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT64), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(G190gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n298), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT24), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT24), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n302), .A2(KEYINPUT65), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT64), .B(G183gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT65), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n309), .A3(new_n301), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n296), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT25), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n304), .A2(new_n306), .B1(new_n297), .B2(new_n301), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n292), .A2(new_n294), .A3(new_n295), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT66), .B1(new_n311), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT65), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n304), .A2(new_n306), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(new_n310), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n296), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT66), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(new_n323), .A3(new_n315), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT68), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n298), .A2(new_n300), .A3(KEYINPUT67), .A4(KEYINPUT27), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n297), .A2(KEYINPUT27), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(G190gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT67), .B1(new_n308), .B2(KEYINPUT27), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n326), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT28), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n298), .A2(new_n300), .A3(KEYINPUT27), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT67), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n336), .A2(KEYINPUT68), .A3(new_n329), .A4(new_n327), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n332), .A2(new_n333), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT27), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n329), .B(KEYINPUT28), .C1(new_n339), .C2(G183gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NOR3_X1   g140(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT69), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n290), .A2(new_n291), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT26), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n295), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n303), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n341), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G226gat), .A2(G233gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n325), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT29), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n347), .B1(new_n338), .B2(new_n340), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n311), .A2(new_n316), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n353), .B(new_n350), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n289), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT77), .B(KEYINPUT29), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n317), .A2(new_n324), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n359), .B1(new_n360), .B2(new_n354), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n350), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n363), .B(new_n351), .C1(new_n354), .C2(new_n355), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n351), .B1(new_n354), .B2(new_n355), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT78), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n362), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n357), .B1(new_n367), .B2(new_n289), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT37), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n281), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n289), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n350), .A2(new_n361), .B1(new_n365), .B2(KEYINPUT78), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(new_n364), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT37), .B1(new_n373), .B2(new_n357), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT38), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT72), .ZN(new_n377));
  INV_X1    g176(.A(G134gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(G127gat), .ZN(new_n379));
  INV_X1    g178(.A(G127gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(G134gat), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n377), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT71), .ZN(new_n383));
  INV_X1    g182(.A(G120gat), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n383), .B1(new_n384), .B2(G113gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(G113gat), .ZN(new_n386));
  INV_X1    g185(.A(G113gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(KEYINPUT71), .A3(G120gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT1), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n380), .A2(G134gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n378), .A2(G127gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT72), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n382), .A2(new_n389), .A3(new_n390), .A4(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT70), .ZN(new_n395));
  OR3_X1    g194(.A1(new_n378), .A2(KEYINPUT70), .A3(G127gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(G113gat), .B(G120gat), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n395), .B(new_n396), .C1(KEYINPUT1), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(G141gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(G148gat), .ZN(new_n401));
  INV_X1    g200(.A(G148gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(G141gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G155gat), .ZN(new_n405));
  INV_X1    g204(.A(G162gat), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT2), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G155gat), .B(G162gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n404), .A2(new_n409), .A3(new_n407), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n399), .B(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(G225gat), .A2(G233gat), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(KEYINPUT5), .A3(new_n416), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n399), .A2(new_n413), .A3(KEYINPUT4), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT4), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n394), .A2(new_n398), .ZN(new_n420));
  INV_X1    g219(.A(new_n413), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n412), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n409), .B1(new_n407), .B2(new_n404), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT3), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT3), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n411), .A2(new_n426), .A3(new_n412), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n425), .A2(new_n399), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n418), .B1(new_n422), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n429), .A2(new_n416), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n420), .A2(new_n421), .A3(new_n419), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n425), .A2(new_n399), .A3(new_n427), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT4), .B1(new_n399), .B2(new_n413), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n430), .B1(new_n436), .B2(new_n415), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n417), .B1(new_n432), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(G1gat), .B(G29gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(KEYINPUT0), .ZN(new_n440));
  XNOR2_X1  g239(.A(G57gat), .B(G85gat), .ZN(new_n441));
  XOR2_X1   g240(.A(new_n440), .B(new_n441), .Z(new_n442));
  AOI21_X1  g241(.A(KEYINPUT6), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n442), .ZN(new_n444));
  INV_X1    g243(.A(new_n417), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n431), .B1(new_n429), .B2(new_n416), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n436), .A2(new_n415), .A3(new_n430), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n444), .B1(new_n448), .B2(KEYINPUT86), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT86), .ZN(new_n450));
  AOI211_X1 g249(.A(new_n450), .B(new_n445), .C1(new_n446), .C2(new_n447), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n443), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n368), .A2(new_n281), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n438), .A2(new_n454), .A3(new_n442), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n452), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n367), .A2(new_n371), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n352), .A2(new_n356), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n369), .B1(new_n459), .B2(new_n289), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT38), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n370), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n376), .A2(new_n457), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT40), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT39), .B1(new_n414), .B2(new_n416), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n465), .B1(new_n416), .B2(new_n429), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT39), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n429), .A2(new_n467), .A3(new_n416), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n442), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n464), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n465), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n429), .A2(new_n416), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n473), .A2(KEYINPUT40), .A3(new_n442), .A4(new_n468), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n451), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n442), .B1(new_n438), .B2(new_n450), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n281), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n479), .B1(new_n373), .B2(new_n357), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n367), .A2(new_n289), .ZN(new_n481));
  INV_X1    g280(.A(new_n357), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n481), .A2(KEYINPUT30), .A3(new_n482), .A4(new_n281), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  XOR2_X1   g283(.A(KEYINPUT80), .B(KEYINPUT30), .Z(new_n485));
  AOI21_X1  g284(.A(new_n485), .B1(new_n368), .B2(new_n281), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n478), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT87), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n373), .A2(new_n357), .A3(new_n479), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n483), .B(new_n480), .C1(new_n490), .C2(new_n485), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n491), .A2(KEYINPUT87), .A3(new_n478), .ZN(new_n492));
  XOR2_X1   g291(.A(G78gat), .B(G106gat), .Z(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT31), .B(G50gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT84), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT83), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n289), .A2(new_n499), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n288), .A2(new_n282), .A3(new_n286), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n358), .B1(new_n501), .B2(KEYINPUT83), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n498), .B(new_n413), .C1(new_n503), .C2(KEYINPUT3), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT3), .B1(new_n500), .B2(new_n502), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT84), .B1(new_n505), .B2(new_n421), .ZN(new_n506));
  NAND2_X1  g305(.A1(G228gat), .A2(G233gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n427), .A2(new_n359), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(new_n289), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n504), .A2(new_n506), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G22gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n371), .A2(new_n353), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n421), .B1(new_n512), .B2(new_n426), .ZN(new_n513));
  INV_X1    g312(.A(new_n509), .ZN(new_n514));
  OAI211_X1 g313(.A(G228gat), .B(G233gat), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n510), .A2(new_n511), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n511), .B1(new_n510), .B2(new_n515), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n497), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n518), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n495), .B(new_n496), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n516), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n463), .A2(new_n489), .A3(new_n492), .A4(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n491), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n454), .B1(new_n448), .B2(new_n444), .ZN(new_n526));
  OAI22_X1  g325(.A1(new_n526), .A2(KEYINPUT82), .B1(new_n438), .B2(new_n442), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n526), .A2(KEYINPUT82), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n456), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n523), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n325), .A2(new_n349), .A3(new_n399), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n420), .B1(new_n360), .B2(new_n354), .ZN(new_n535));
  NAND2_X1  g334(.A1(G227gat), .A2(G233gat), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G15gat), .B(G43gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(G71gat), .B(G99gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT33), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT73), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n538), .A2(KEYINPUT32), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n534), .A2(new_n535), .A3(new_n537), .A4(new_n542), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n544), .B1(new_n548), .B2(new_n543), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n538), .A2(KEYINPUT32), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n547), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT34), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n534), .A2(new_n535), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(new_n554), .B2(new_n536), .ZN(new_n555));
  AOI211_X1 g354(.A(KEYINPUT34), .B(new_n537), .C1(new_n534), .C2(new_n535), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n533), .B1(new_n552), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT74), .B1(new_n555), .B2(new_n556), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n399), .B1(new_n325), .B2(new_n349), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n360), .A2(new_n354), .A3(new_n420), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n536), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT34), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT74), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n554), .A2(new_n553), .A3(new_n536), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n559), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT75), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n548), .A2(new_n543), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT73), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n546), .B1(new_n570), .B2(new_n550), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n567), .A2(new_n568), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n568), .B1(new_n567), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n558), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n552), .A2(new_n557), .ZN(new_n575));
  INV_X1    g374(.A(new_n557), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n524), .A2(new_n532), .A3(new_n581), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n552), .A2(new_n557), .B1(new_n519), .B2(new_n522), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n583), .B1(new_n572), .B2(new_n573), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT35), .B1(new_n584), .B2(new_n530), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n578), .A2(new_n531), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT35), .B1(new_n452), .B2(new_n456), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n525), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n277), .B1(new_n582), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n529), .ZN(new_n591));
  AND2_X1   g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n592), .A2(KEYINPUT41), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT103), .ZN(new_n594));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G99gat), .B(G106gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(G85gat), .A2(G92gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT7), .ZN(new_n600));
  NOR2_X1   g399(.A1(G85gat), .A2(G92gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n601), .B1(KEYINPUT8), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n598), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT104), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n600), .A2(new_n603), .ZN(new_n607));
  INV_X1    g406(.A(new_n598), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n600), .A2(new_n598), .A3(new_n603), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(KEYINPUT104), .A3(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n248), .A2(new_n249), .A3(new_n606), .A4(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G190gat), .B(G218gat), .Z(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n606), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n244), .A2(new_n615), .B1(KEYINPUT41), .B2(new_n592), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n612), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n614), .B1(new_n612), .B2(new_n616), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n597), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n619), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n621), .A2(new_n596), .A3(new_n617), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G183gat), .B(G211gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT102), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(new_n405), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n625), .B(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT21), .ZN(new_n630));
  XNOR2_X1  g429(.A(G71gat), .B(G78gat), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G57gat), .B(G64gat), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n631), .B(new_n634), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(G71gat), .ZN(new_n640));
  INV_X1    g439(.A(G78gat), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n640), .A2(new_n641), .A3(KEYINPUT98), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT98), .B1(new_n640), .B2(new_n641), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n640), .A2(new_n641), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n632), .B(KEYINPUT99), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n645), .B1(new_n646), .B2(new_n635), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n639), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n261), .B1(new_n630), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT101), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n630), .ZN(new_n651));
  NAND2_X1  g450(.A1(G231gat), .A2(G233gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G127gat), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n650), .A2(new_n655), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n629), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n658), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n660), .A2(new_n656), .A3(new_n628), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n623), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT105), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT10), .ZN(new_n664));
  AOI22_X1  g463(.A1(new_n611), .A2(new_n606), .B1(new_n639), .B2(new_n647), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n600), .A2(new_n598), .A3(new_n603), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n604), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n648), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n664), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n639), .A2(new_n647), .A3(KEYINPUT10), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n670), .B1(new_n606), .B2(new_n611), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(G230gat), .A2(G233gat), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n663), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n674), .ZN(new_n676));
  AOI211_X1 g475(.A(KEYINPUT105), .B(new_n676), .C1(new_n669), .C2(new_n672), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n648), .A2(new_n667), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n666), .A2(new_n604), .A3(new_n605), .ZN(new_n680));
  INV_X1    g479(.A(new_n606), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n648), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n679), .A2(new_n682), .A3(new_n676), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G120gat), .B(G148gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(G176gat), .B(G204gat), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n685), .B(new_n686), .Z(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n678), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n679), .A2(new_n682), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n671), .B1(new_n691), .B2(new_n664), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n676), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n688), .B1(new_n693), .B2(new_n684), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n662), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n590), .A2(new_n591), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(G1gat), .ZN(G1324gat));
  AND3_X1   g499(.A1(new_n590), .A2(new_n491), .A3(new_n698), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT16), .B(G8gat), .Z(new_n702));
  AND2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n701), .A2(new_n214), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT42), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n705), .B1(KEYINPUT42), .B2(new_n703), .ZN(G1325gat));
  NAND2_X1  g505(.A1(new_n590), .A2(new_n698), .ZN(new_n707));
  OAI21_X1  g506(.A(G15gat), .B1(new_n707), .B2(new_n581), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n697), .A2(G15gat), .A3(new_n578), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n590), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(G1326gat));
  NOR2_X1   g510(.A1(new_n707), .A2(new_n523), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT43), .B(G22gat), .Z(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1327gat));
  NAND2_X1  g513(.A1(new_n659), .A2(new_n661), .ZN(new_n715));
  INV_X1    g514(.A(new_n623), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n715), .A2(new_n716), .A3(new_n695), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n590), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(new_n591), .A3(new_n236), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT45), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n582), .A2(new_n589), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT107), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n582), .A2(new_n589), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n716), .A2(KEYINPUT44), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n723), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n722), .A2(new_n623), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT44), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n695), .B(KEYINPUT106), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n732), .A2(new_n715), .A3(new_n277), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n529), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n721), .B1(new_n236), .B2(new_n735), .ZN(G1328gat));
  NOR3_X1   g535(.A1(new_n718), .A2(G36gat), .A3(new_n525), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT46), .ZN(new_n738));
  OAI21_X1  g537(.A(G36gat), .B1(new_n734), .B2(new_n525), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1329gat));
  OAI21_X1  g539(.A(G43gat), .B1(new_n734), .B2(new_n581), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT108), .ZN(new_n742));
  OR3_X1    g541(.A1(new_n718), .A2(G43gat), .A3(new_n578), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n742), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n741), .B(new_n743), .C1(KEYINPUT108), .C2(KEYINPUT47), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(G1330gat));
  AND3_X1   g547(.A1(new_n582), .A2(new_n589), .A3(new_n724), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n724), .B1(new_n582), .B2(new_n589), .ZN(new_n750));
  INV_X1    g549(.A(new_n726), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n716), .B1(new_n582), .B2(new_n589), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT44), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n531), .B(new_n733), .C1(new_n752), .C2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n730), .A2(KEYINPUT110), .A3(new_n531), .A4(new_n733), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n758), .A2(G50gat), .A3(new_n759), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n718), .A2(G50gat), .A3(new_n523), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(KEYINPUT48), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n733), .ZN(new_n764));
  AOI211_X1 g563(.A(new_n523), .B(new_n764), .C1(new_n727), .C2(new_n729), .ZN(new_n765));
  INV_X1    g564(.A(G50gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n762), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT48), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT109), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n761), .B1(new_n756), .B2(G50gat), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n770), .A2(new_n771), .A3(KEYINPUT48), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n763), .B1(new_n769), .B2(new_n772), .ZN(G1331gat));
  NOR2_X1   g572(.A1(new_n749), .A2(new_n750), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n662), .A2(new_n277), .A3(new_n732), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n591), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g577(.A1(new_n774), .A2(new_n775), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(new_n525), .ZN(new_n780));
  NOR2_X1   g579(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n781));
  AND2_X1   g580(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(new_n780), .B2(new_n781), .ZN(G1333gat));
  INV_X1    g583(.A(new_n578), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n776), .A2(new_n640), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G71gat), .B1(new_n779), .B2(new_n581), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n788), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g588(.A1(new_n779), .A2(new_n523), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(new_n641), .ZN(G1335gat));
  NOR2_X1   g590(.A1(new_n715), .A2(new_n276), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n695), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n727), .B2(new_n729), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G85gat), .B1(new_n795), .B2(new_n529), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n753), .A2(new_n792), .ZN(new_n797));
  NOR2_X1   g596(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n797), .B1(new_n800), .B2(new_n798), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(KEYINPUT112), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT112), .B1(new_n799), .B2(new_n801), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n695), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n529), .A2(G85gat), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n796), .B1(new_n805), .B2(new_n806), .ZN(G1336gat));
  NAND2_X1  g606(.A1(new_n799), .A2(new_n801), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n731), .A2(new_n525), .A3(G92gat), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT52), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n491), .ZN(new_n811));
  OAI21_X1  g610(.A(G92gat), .B1(new_n811), .B2(KEYINPUT115), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n794), .B2(new_n491), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n810), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n722), .A2(KEYINPUT113), .A3(new_n623), .A4(new_n792), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT51), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(KEYINPUT51), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n753), .A2(new_n792), .B1(KEYINPUT113), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n811), .A2(G92gat), .B1(new_n821), .B2(new_n809), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n815), .B1(new_n822), .B2(new_n823), .ZN(G1337gat));
  OAI21_X1  g623(.A(G99gat), .B1(new_n795), .B2(new_n581), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n578), .A2(G99gat), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n805), .B2(new_n826), .ZN(G1338gat));
  NOR3_X1   g626(.A1(new_n731), .A2(G106gat), .A3(new_n523), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT116), .B1(new_n821), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(G106gat), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(new_n794), .B2(new_n531), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832));
  INV_X1    g631(.A(new_n828), .ZN(new_n833));
  NOR4_X1   g632(.A1(new_n818), .A2(new_n820), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n829), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n836));
  INV_X1    g635(.A(new_n808), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n833), .ZN(new_n838));
  OAI22_X1  g637(.A1(new_n835), .A2(new_n836), .B1(new_n838), .B2(new_n831), .ZN(G1339gat));
  INV_X1    g638(.A(new_n715), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n669), .A2(new_n672), .A3(new_n676), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT54), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n675), .A2(new_n677), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n673), .A2(new_n674), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n688), .B1(new_n845), .B2(KEYINPUT54), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n841), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(KEYINPUT105), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n673), .A2(new_n663), .A3(new_n674), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n850), .B1(new_n692), .B2(new_n676), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n687), .B1(new_n693), .B2(new_n850), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n853), .A3(KEYINPUT55), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n847), .A2(new_n690), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n264), .A2(new_n265), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n246), .B1(new_n245), .B2(new_n250), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n259), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n270), .A2(new_n623), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n855), .A2(new_n859), .A3(KEYINPUT117), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n847), .A2(new_n690), .A3(new_n854), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n270), .A2(new_n623), .A3(new_n858), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n846), .B1(new_n678), .B2(new_n851), .ZN(new_n866));
  AOI22_X1  g665(.A1(new_n866), .A2(KEYINPUT55), .B1(new_n678), .B2(new_n689), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n276), .A3(new_n847), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n270), .A2(new_n695), .A3(new_n858), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n623), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n840), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n662), .A2(new_n277), .A3(new_n696), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n586), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n529), .A2(new_n491), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(G113gat), .B1(new_n878), .B2(new_n277), .ZN(new_n879));
  AOI211_X1 g678(.A(new_n529), .B(new_n584), .C1(new_n871), .C2(new_n872), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n525), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT118), .Z(new_n882));
  NAND2_X1  g681(.A1(new_n276), .A2(new_n387), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n879), .B1(new_n882), .B2(new_n883), .ZN(G1340gat));
  OAI21_X1  g683(.A(G120gat), .B1(new_n878), .B2(new_n731), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n695), .A2(new_n384), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n882), .B2(new_n886), .ZN(G1341gat));
  NOR3_X1   g686(.A1(new_n881), .A2(G127gat), .A3(new_n840), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n380), .B1(new_n877), .B2(new_n715), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT119), .ZN(G1342gat));
  NAND4_X1  g690(.A1(new_n880), .A2(new_n378), .A3(new_n525), .A4(new_n623), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n892), .A2(KEYINPUT56), .ZN(new_n893));
  OAI21_X1  g692(.A(G134gat), .B1(new_n878), .B2(new_n716), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(KEYINPUT56), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(G1343gat));
  NAND2_X1  g695(.A1(new_n873), .A2(new_n531), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(KEYINPUT57), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT57), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT120), .B1(new_n844), .B2(new_n846), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n852), .A2(new_n853), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n900), .A2(new_n841), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n276), .A3(new_n867), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n623), .B1(new_n904), .B2(new_n869), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n840), .B1(new_n865), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n872), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n899), .B1(new_n907), .B2(new_n531), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n581), .A2(new_n875), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n898), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n400), .B1(new_n910), .B2(new_n276), .ZN(new_n911));
  AND4_X1   g710(.A1(new_n531), .A2(new_n873), .A3(new_n591), .A4(new_n581), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NOR4_X1   g712(.A1(new_n913), .A2(G141gat), .A3(new_n491), .A4(new_n277), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n915), .B(new_n916), .ZN(G1344gat));
  NAND4_X1  g716(.A1(new_n912), .A2(new_n402), .A3(new_n525), .A4(new_n695), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n909), .A2(new_n696), .ZN(new_n920));
  AOI211_X1 g719(.A(new_n899), .B(new_n523), .C1(new_n871), .C2(new_n872), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n862), .A2(new_n863), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n840), .B1(new_n905), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n523), .B1(new_n924), .B2(new_n872), .ZN(new_n925));
  OAI22_X1  g724(.A1(new_n921), .A2(new_n922), .B1(KEYINPUT57), .B2(new_n925), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n897), .A2(KEYINPUT121), .A3(new_n899), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n920), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n919), .B1(new_n928), .B2(G148gat), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n919), .A2(G148gat), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n930), .B1(new_n910), .B2(new_n695), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n918), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT122), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n934), .B(new_n918), .C1(new_n929), .C2(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1345gat));
  NAND4_X1  g735(.A1(new_n912), .A2(new_n405), .A3(new_n525), .A4(new_n715), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n910), .A2(new_n715), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(new_n405), .ZN(G1346gat));
  NAND2_X1  g738(.A1(new_n910), .A2(new_n623), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n406), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n942), .B1(new_n941), .B2(new_n940), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n525), .A2(new_n406), .A3(new_n623), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n913), .B2(new_n944), .ZN(G1347gat));
  NOR2_X1   g744(.A1(new_n591), .A2(new_n525), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n873), .A2(new_n586), .A3(new_n946), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n947), .A2(new_n290), .A3(new_n277), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n591), .B1(new_n871), .B2(new_n872), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n584), .A2(new_n525), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n276), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n948), .B1(new_n954), .B2(new_n290), .ZN(G1348gat));
  OAI21_X1  g754(.A(G176gat), .B1(new_n947), .B2(new_n731), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n695), .A2(new_n291), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n952), .B2(new_n957), .ZN(G1349gat));
  NOR2_X1   g757(.A1(new_n339), .A2(G183gat), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n840), .A2(new_n328), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n953), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n947), .A2(new_n840), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n308), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n964));
  XOR2_X1   g763(.A(new_n963), .B(new_n964), .Z(G1350gat));
  OAI21_X1  g764(.A(G190gat), .B1(new_n947), .B2(new_n716), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT61), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n953), .A2(new_n301), .A3(new_n623), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(G1351gat));
  OR2_X1    g768(.A1(new_n926), .A2(new_n927), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n581), .A2(new_n946), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(G197gat), .B1(new_n972), .B2(new_n277), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n949), .A2(new_n491), .A3(new_n531), .A4(new_n581), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n974), .A2(G197gat), .A3(new_n277), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT125), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n973), .A2(new_n976), .ZN(G1352gat));
  XOR2_X1   g776(.A(KEYINPUT126), .B(G204gat), .Z(new_n978));
  OAI21_X1  g777(.A(new_n978), .B1(new_n972), .B2(new_n731), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n974), .A2(new_n696), .A3(new_n978), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT62), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n979), .A2(new_n981), .ZN(G1353gat));
  NAND3_X1  g781(.A1(new_n970), .A2(new_n715), .A3(new_n971), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n983), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n984));
  AOI21_X1  g783(.A(KEYINPUT63), .B1(new_n983), .B2(G211gat), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n715), .A2(new_n284), .ZN(new_n986));
  OAI22_X1  g785(.A1(new_n984), .A2(new_n985), .B1(new_n974), .B2(new_n986), .ZN(G1354gat));
  OAI21_X1  g786(.A(G218gat), .B1(new_n972), .B2(new_n716), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n623), .A2(new_n285), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n988), .B1(new_n974), .B2(new_n989), .ZN(G1355gat));
endmodule


