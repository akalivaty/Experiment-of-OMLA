//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT75), .B(G902), .Z(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G234), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT68), .B(G128), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT23), .A3(G119), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  AOI21_X1  g007(.A(KEYINPUT23), .B1(new_n193), .B2(G119), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(G119), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n195), .B1(new_n191), .B2(G119), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT24), .B(G110), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n197), .A2(G110), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G125), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G140), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT77), .ZN(new_n206));
  OR3_X1    g020(.A1(new_n204), .A2(KEYINPUT77), .A3(G140), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT16), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n203), .A2(new_n210), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n208), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n209), .B1(new_n208), .B2(new_n211), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n201), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OAI22_X1  g028(.A1(new_n197), .A2(G110), .B1(new_n198), .B2(new_n200), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n208), .A2(new_n211), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G146), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n203), .A2(new_n205), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n215), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT22), .B(G137), .ZN(new_n222));
  INV_X1    g036(.A(G953), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n223), .A2(G221), .A3(G234), .ZN(new_n224));
  XOR2_X1   g038(.A(new_n222), .B(new_n224), .Z(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n214), .A2(new_n220), .A3(new_n225), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n188), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OR2_X1    g045(.A1(new_n231), .A2(KEYINPUT25), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(KEYINPUT25), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n190), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n189), .A2(G902), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n235), .B(KEYINPUT78), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n229), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G116), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n240), .A2(G119), .ZN(new_n241));
  INV_X1    g055(.A(G119), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT69), .B1(new_n242), .B2(G116), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(new_n240), .A3(G119), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n241), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT2), .B(G113), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n248), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G137), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT11), .A3(G134), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G137), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT67), .A2(G131), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT67), .A2(G131), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT11), .ZN(new_n262));
  OAI211_X1 g076(.A(KEYINPUT66), .B(new_n262), .C1(new_n256), .C2(G137), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n254), .A2(G134), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT66), .B1(new_n265), .B2(new_n262), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n258), .B(new_n261), .C1(new_n264), .C2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G131), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n255), .A2(new_n257), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n262), .B1(new_n256), .B2(G137), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT66), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n269), .B1(new_n272), .B2(new_n263), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n267), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(G143), .B(G146), .ZN(new_n275));
  NAND2_X1  g089(.A1(KEYINPUT0), .A2(G128), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G143), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT64), .B1(new_n279), .B2(G146), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT64), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(new_n209), .A3(G143), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT65), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n284), .B1(new_n209), .B2(G143), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n279), .A2(KEYINPUT65), .A3(G146), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(KEYINPUT0), .A2(G128), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n277), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n278), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n274), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT1), .B1(new_n279), .B2(G146), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n193), .A2(KEYINPUT68), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n193), .A2(KEYINPUT68), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n280), .A2(new_n282), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n285), .A2(new_n286), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n279), .A2(G146), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n209), .A2(G143), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n268), .B1(new_n265), .B2(new_n257), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n304), .B1(new_n273), .B2(new_n261), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n303), .B1(new_n305), .B2(KEYINPUT70), .ZN(new_n306));
  INV_X1    g120(.A(new_n304), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n267), .A2(KEYINPUT70), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n253), .B(new_n291), .C1(new_n306), .C2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n267), .A2(new_n307), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT70), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n303), .A3(new_n308), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n316), .A2(KEYINPUT71), .A3(new_n253), .A4(new_n291), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n291), .B1(new_n306), .B2(new_n309), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n252), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n312), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT28), .ZN(new_n321));
  NOR2_X1   g135(.A1(G237), .A2(G953), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G210), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(KEYINPUT27), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT26), .B(G101), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n324), .B(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT28), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n327), .B1(new_n310), .B2(new_n328), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n329), .A2(KEYINPUT29), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n321), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT74), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n321), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n310), .A2(new_n328), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n326), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n303), .A2(new_n305), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n291), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n252), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n312), .A2(new_n340), .A3(new_n317), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n337), .B1(new_n341), .B2(KEYINPUT28), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT72), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n318), .A2(KEYINPUT30), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT30), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n291), .A2(new_n338), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n253), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n312), .A2(new_n317), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n327), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT73), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI211_X1 g165(.A(KEYINPUT73), .B(new_n327), .C1(new_n347), .C2(new_n348), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n343), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT29), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n342), .B2(KEYINPUT72), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n335), .B(new_n188), .C1(new_n353), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G472), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT76), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(KEYINPUT76), .A3(G472), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT32), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n345), .B1(new_n316), .B2(new_n291), .ZN(new_n363));
  INV_X1    g177(.A(new_n346), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n252), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n365), .A2(new_n312), .A3(new_n317), .A4(new_n326), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT31), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n348), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n369), .A2(KEYINPUT31), .A3(new_n326), .A4(new_n365), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n341), .A2(KEYINPUT28), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n336), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n368), .A2(new_n370), .B1(new_n372), .B2(new_n327), .ZN(new_n373));
  NOR2_X1   g187(.A1(G472), .A2(G902), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n362), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n368), .A2(new_n370), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n372), .A2(new_n327), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(KEYINPUT32), .A3(new_n374), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n239), .B1(new_n361), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT86), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT9), .B(G234), .ZN(new_n384));
  OAI21_X1  g198(.A(G221), .B1(new_n384), .B2(G902), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G107), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n387), .B1(new_n388), .B2(G104), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(G104), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n392), .A2(KEYINPUT3), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n387), .A2(KEYINPUT79), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT79), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G107), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G101), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n391), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(G104), .B2(G107), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n394), .A2(new_n396), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n400), .B1(new_n401), .B2(G104), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n298), .A3(new_n302), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT84), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n193), .B1(new_n301), .B2(KEYINPUT1), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n302), .B1(new_n406), .B2(new_n275), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(new_n399), .A3(new_n402), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n287), .A2(new_n295), .B1(new_n275), .B2(new_n299), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT84), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(new_n403), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n405), .A2(new_n408), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(KEYINPUT12), .A3(new_n274), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT85), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT85), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n412), .A2(new_n415), .A3(KEYINPUT12), .A4(new_n274), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n274), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT12), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n414), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n408), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT82), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT82), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n408), .A2(new_n424), .A3(new_n421), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n274), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n391), .A2(new_n397), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT80), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n391), .A2(new_n397), .A3(KEYINPUT80), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n430), .A2(new_n431), .A3(G101), .A4(new_n432), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n391), .A2(new_n397), .A3(KEYINPUT80), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT80), .B1(new_n391), .B2(new_n397), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n434), .A2(new_n435), .A3(new_n398), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n399), .A2(KEYINPUT4), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n433), .B(new_n290), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n399), .A2(new_n402), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n303), .A2(new_n439), .A3(KEYINPUT10), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n426), .A2(new_n427), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n303), .A2(new_n439), .A3(KEYINPUT10), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(new_n423), .B2(new_n425), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n445), .A2(KEYINPUT83), .A3(new_n427), .A4(new_n438), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n420), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(G110), .B(G140), .ZN(new_n449));
  INV_X1    g263(.A(G227), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(G953), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n449), .B(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n445), .A2(new_n438), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n274), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n452), .B1(new_n443), .B2(new_n446), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n448), .A2(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G469), .B1(new_n456), .B2(G902), .ZN(new_n457));
  INV_X1    g271(.A(G469), .ZN(new_n458));
  INV_X1    g272(.A(new_n452), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n420), .A2(new_n447), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n459), .B1(new_n447), .B2(new_n454), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n458), .B(new_n188), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  AOI211_X1 g276(.A(new_n383), .B(new_n386), .C1(new_n457), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(G469), .A2(G902), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n448), .A2(new_n452), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n455), .A2(new_n454), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(G469), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n462), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT86), .B1(new_n468), .B2(new_n385), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT88), .B1(new_n290), .B2(new_n204), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT88), .ZN(new_n471));
  INV_X1    g285(.A(new_n289), .ZN(new_n472));
  INV_X1    g286(.A(new_n297), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n472), .B1(new_n473), .B2(new_n283), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n471), .B(G125), .C1(new_n474), .C2(new_n278), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n409), .A2(new_n204), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n470), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G224), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(G953), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n477), .B(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n433), .B(new_n252), .C1(new_n436), .C2(new_n437), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n242), .A2(G116), .ZN(new_n482));
  OAI21_X1  g296(.A(G113), .B1(new_n482), .B2(KEYINPUT5), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n483), .B1(new_n246), .B2(KEYINPUT5), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n439), .A2(new_n485), .A3(new_n251), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(G110), .B(G122), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n481), .A2(new_n488), .A3(new_n486), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(KEYINPUT6), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n488), .B1(new_n481), .B2(new_n486), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT87), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT6), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n494), .B1(new_n493), .B2(new_n495), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n480), .B(new_n492), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  XOR2_X1   g312(.A(new_n488), .B(KEYINPUT8), .Z(new_n499));
  INV_X1    g313(.A(new_n251), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n403), .B1(new_n500), .B2(new_n484), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n486), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT89), .B1(new_n303), .B2(G125), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT89), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n409), .A2(new_n504), .A3(new_n204), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n503), .A2(new_n470), .A3(new_n475), .A4(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n479), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT7), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n502), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n470), .A2(new_n475), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n510), .A2(KEYINPUT7), .A3(new_n476), .A4(new_n507), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n511), .A3(new_n491), .ZN(new_n512));
  INV_X1    g326(.A(G902), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n498), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(G210), .B1(G237), .B2(G902), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n516), .B(KEYINPUT90), .Z(new_n517));
  XOR2_X1   g331(.A(new_n517), .B(KEYINPUT91), .Z(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n517), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n498), .A2(new_n514), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n223), .A2(G952), .ZN(new_n524));
  INV_X1    g338(.A(G234), .ZN(new_n525));
  INV_X1    g339(.A(G237), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  AOI211_X1 g342(.A(new_n223), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT21), .B(G898), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(G214), .B1(G237), .B2(G902), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n523), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n463), .A2(new_n469), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n526), .A2(new_n223), .A3(G214), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n279), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n322), .A2(G143), .A3(G214), .ZN(new_n538));
  NAND2_X1  g352(.A1(KEYINPUT18), .A2(G131), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n539), .B1(new_n537), .B2(new_n538), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n206), .A2(new_n207), .A3(G146), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT92), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n543), .A2(new_n219), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n544), .B1(new_n543), .B2(new_n219), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n208), .A2(new_n209), .A3(new_n211), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n259), .A2(new_n260), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n322), .A2(G143), .A3(G214), .ZN(new_n551));
  AOI21_X1  g365(.A(G143), .B1(new_n322), .B2(G214), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n550), .B(KEYINPUT17), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n217), .A2(new_n549), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n537), .A2(new_n261), .A3(new_n538), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT93), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT93), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n537), .A2(new_n558), .A3(new_n261), .A4(new_n538), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT17), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n554), .A2(KEYINPUT95), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n553), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n212), .A2(new_n213), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT95), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n548), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(G113), .B(G122), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(new_n392), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n569), .ZN(new_n571));
  AOI211_X1 g385(.A(new_n571), .B(new_n548), .C1(new_n562), .C2(new_n566), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n513), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(G475), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT19), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(new_n206), .B2(new_n207), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n218), .A2(KEYINPUT19), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n209), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(new_n217), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n547), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n571), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT94), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT94), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(new_n584), .A3(new_n571), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n583), .A2(new_n585), .B1(new_n567), .B2(new_n569), .ZN(new_n586));
  NOR2_X1   g400(.A1(G475), .A2(G902), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(KEYINPUT96), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT20), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  OAI22_X1  g403(.A1(new_n564), .A2(new_n565), .B1(KEYINPUT17), .B2(new_n575), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n554), .A2(KEYINPUT95), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n569), .B(new_n547), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n584), .B1(new_n581), .B2(new_n571), .ZN(new_n593));
  AOI211_X1 g407(.A(KEYINPUT94), .B(new_n569), .C1(new_n580), .C2(new_n547), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT20), .ZN(new_n596));
  INV_X1    g410(.A(new_n588), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n595), .A2(KEYINPUT97), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n589), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n583), .A2(new_n585), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n588), .B1(new_n600), .B2(new_n592), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT97), .B1(new_n601), .B2(new_n596), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n574), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT98), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n593), .A2(new_n594), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n596), .B(new_n597), .C1(new_n605), .C2(new_n572), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(new_n598), .A3(new_n589), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n610), .A3(new_n574), .ZN(new_n611));
  INV_X1    g425(.A(G478), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(KEYINPUT15), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n191), .A2(G143), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT13), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n279), .A2(G128), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT13), .B1(new_n279), .B2(G128), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT99), .ZN(new_n620));
  OAI21_X1  g434(.A(G134), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n615), .A2(new_n617), .ZN(new_n622));
  INV_X1    g436(.A(G122), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(G116), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n240), .A2(G122), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n401), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n401), .A2(new_n626), .ZN(new_n628));
  OAI221_X1 g442(.A(new_n621), .B1(G134), .B2(new_n622), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n622), .B(G134), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n625), .A2(KEYINPUT14), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n240), .A2(G122), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n625), .B1(new_n632), .B2(KEYINPUT14), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n631), .B1(new_n633), .B2(KEYINPUT100), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n634), .B1(KEYINPUT100), .B2(new_n633), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(G107), .ZN(new_n636));
  INV_X1    g450(.A(new_n628), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n630), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n629), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n384), .A2(new_n187), .A3(G953), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n614), .B1(new_n642), .B2(new_n188), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n641), .A2(new_n230), .A3(new_n613), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n604), .A2(new_n611), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n382), .A2(new_n535), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G101), .ZN(G3));
  NAND2_X1  g463(.A1(new_n468), .A2(new_n385), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n383), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n386), .B1(new_n457), .B2(new_n462), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT86), .ZN(new_n653));
  OAI21_X1  g467(.A(G472), .B1(new_n373), .B2(new_n230), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n379), .A2(new_n374), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n654), .A2(new_n238), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n651), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT101), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n651), .A2(new_n653), .A3(KEYINPUT101), .A4(new_n656), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n533), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n515), .A2(new_n517), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n662), .B1(new_n663), .B2(new_n522), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n604), .A2(new_n611), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n642), .A2(new_n188), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n612), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT33), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n669), .B1(new_n639), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n641), .B(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n230), .A2(new_n612), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n668), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n666), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n661), .A2(new_n532), .A3(new_n664), .A4(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT34), .B(G104), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G6));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n595), .A2(new_n681), .A3(new_n596), .A4(new_n597), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n574), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n589), .A2(KEYINPUT103), .A3(new_n606), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n645), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n522), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n521), .B1(new_n498), .B2(new_n514), .ZN(new_n689));
  OAI211_X1 g503(.A(new_n532), .B(new_n533), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n661), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT35), .B(G107), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G9));
  NAND2_X1  g508(.A1(new_n654), .A2(new_n655), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n226), .A2(KEYINPUT36), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n221), .B(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n236), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n234), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n535), .A2(new_n647), .A3(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT37), .B(G110), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G12));
  INV_X1    g518(.A(G472), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n371), .A2(new_n329), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT72), .ZN(new_n707));
  AOI21_X1  g521(.A(KEYINPUT29), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n708), .A2(new_n343), .A3(new_n351), .A4(new_n352), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n230), .B1(new_n332), .B2(new_n334), .ZN(new_n710));
  AOI211_X1 g524(.A(new_n358), .B(new_n705), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT76), .B1(new_n356), .B2(G472), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n381), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n463), .A2(new_n469), .ZN(new_n714));
  INV_X1    g528(.A(new_n700), .ZN(new_n715));
  AND4_X1   g529(.A1(new_n713), .A2(new_n714), .A3(new_n664), .A4(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(G900), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n528), .B1(new_n529), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n687), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G128), .ZN(G30));
  XNOR2_X1  g535(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n523), .B(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n366), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n320), .A2(new_n327), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n513), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(G472), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n376), .A2(new_n380), .A3(new_n727), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n609), .A2(new_n610), .A3(new_n574), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n610), .B1(new_n609), .B2(new_n574), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n686), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n731), .A2(new_n662), .A3(new_n715), .ZN(new_n732));
  AOI211_X1 g546(.A(new_n723), .B(new_n728), .C1(new_n732), .C2(KEYINPUT105), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n718), .B(KEYINPUT39), .Z(new_n734));
  NAND2_X1  g548(.A1(new_n714), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n736), .A2(KEYINPUT40), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(KEYINPUT40), .ZN(new_n738));
  OAI221_X1 g552(.A(new_n733), .B1(KEYINPUT105), .B2(new_n732), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G143), .ZN(G45));
  INV_X1    g554(.A(new_n718), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n675), .B(new_n741), .C1(new_n729), .C2(new_n730), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT106), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n665), .A2(new_n744), .A3(new_n675), .A4(new_n741), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n716), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G146), .ZN(G48));
  AOI211_X1 g562(.A(new_n676), .B(new_n690), .C1(new_n604), .C2(new_n611), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n447), .A2(new_n454), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n750), .A2(new_n452), .B1(new_n455), .B2(new_n420), .ZN(new_n751));
  OAI21_X1  g565(.A(G469), .B1(new_n751), .B2(new_n230), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n462), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n386), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n713), .A2(new_n749), .A3(new_n238), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT41), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G113), .ZN(G15));
  NAND4_X1  g571(.A1(new_n713), .A2(new_n238), .A3(new_n691), .A4(new_n754), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G116), .ZN(G18));
  NAND4_X1  g573(.A1(new_n664), .A2(new_n385), .A3(new_n462), .A4(new_n752), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n646), .A2(new_n760), .A3(new_n531), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n713), .A3(new_n715), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G119), .ZN(G21));
  NAND2_X1  g577(.A1(new_n731), .A2(KEYINPUT107), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n665), .A2(new_n765), .A3(new_n686), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n760), .A2(new_n531), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n321), .A2(new_n336), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n377), .B1(new_n326), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n374), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n770), .A2(new_n654), .A3(new_n238), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n764), .A2(new_n766), .A3(new_n767), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G122), .ZN(G24));
  NAND3_X1  g587(.A1(new_n715), .A2(new_n770), .A3(new_n654), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n760), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n743), .A2(new_n745), .A3(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n743), .A2(new_n745), .A3(new_n775), .A4(KEYINPUT108), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G125), .ZN(G27));
  AND3_X1   g595(.A1(new_n520), .A2(new_n522), .A3(new_n533), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n468), .A3(new_n385), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT42), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n711), .A2(new_n712), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n380), .A2(KEYINPUT109), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT109), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n379), .A2(new_n788), .A3(KEYINPUT32), .A4(new_n374), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n787), .A2(new_n789), .A3(new_n376), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n238), .B(new_n785), .C1(new_n786), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n743), .A2(new_n745), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n746), .A2(new_n382), .A3(new_n652), .A4(new_n782), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n793), .B1(new_n794), .B2(new_n784), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(new_n268), .ZN(G33));
  NAND4_X1  g610(.A1(new_n382), .A2(new_n652), .A3(new_n719), .A4(new_n782), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G134), .ZN(G36));
  NOR2_X1   g612(.A1(new_n665), .A2(new_n676), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT43), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n695), .A2(new_n715), .ZN(new_n801));
  XOR2_X1   g615(.A(new_n801), .B(KEYINPUT110), .Z(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT44), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n800), .A2(new_n802), .A3(KEYINPUT44), .ZN(new_n806));
  INV_X1    g620(.A(new_n462), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n456), .A2(KEYINPUT45), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n456), .A2(KEYINPUT45), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(G469), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n464), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT46), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n807), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n810), .A2(KEYINPUT46), .A3(new_n464), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n386), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n815), .A2(new_n734), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n805), .A2(new_n782), .A3(new_n806), .A4(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G137), .ZN(G39));
  OR2_X1    g632(.A1(new_n815), .A2(KEYINPUT47), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n815), .A2(KEYINPUT47), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n520), .A2(new_n522), .A3(new_n533), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n713), .A2(new_n238), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n821), .A2(new_n746), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G140), .ZN(G42));
  NAND4_X1  g639(.A1(new_n468), .A2(new_n385), .A3(new_n700), .A4(new_n741), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n728), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n764), .A3(new_n766), .A4(new_n664), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n828), .A2(KEYINPUT116), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(KEYINPUT116), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n747), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n780), .A2(new_n720), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n831), .A2(new_n832), .A3(KEYINPUT52), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n713), .A2(new_n714), .A3(new_n664), .A4(new_n715), .ZN(new_n835));
  OAI22_X1  g649(.A1(new_n835), .A2(new_n792), .B1(new_n828), .B2(KEYINPUT116), .ZN(new_n836));
  INV_X1    g650(.A(new_n830), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n778), .A2(new_n779), .B1(new_n716), .B2(new_n719), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n834), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n833), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n665), .A2(new_n645), .A3(new_n534), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n659), .A2(new_n660), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT112), .B1(new_n843), .B2(new_n702), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n534), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n659), .A2(new_n846), .A3(new_n660), .A4(new_n677), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n648), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n843), .A2(KEYINPUT112), .A3(new_n702), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n845), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n762), .A2(new_n772), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT111), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n852), .A2(new_n853), .A3(new_n755), .A4(new_n758), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n755), .A2(new_n758), .A3(new_n762), .A4(new_n772), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT111), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n783), .A2(new_n774), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n743), .A2(new_n745), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT115), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n743), .A2(new_n745), .A3(new_n859), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT113), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n643), .A2(new_n644), .A3(new_n718), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n685), .A2(new_n782), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n683), .A3(new_n684), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT113), .B1(new_n868), .B2(new_n822), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n713), .A2(new_n714), .A3(new_n715), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n797), .B(new_n864), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n795), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n841), .A2(KEYINPUT53), .A3(new_n858), .A4(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n843), .A2(KEYINPUT112), .A3(new_n702), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n879), .A2(new_n844), .A3(new_n848), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n855), .B(new_n853), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n876), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT52), .B1(new_n831), .B2(new_n832), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n838), .A2(new_n834), .A3(new_n839), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n878), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n877), .A2(new_n886), .A3(KEYINPUT117), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n888), .B(new_n878), .C1(new_n882), .C2(new_n885), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n887), .A2(KEYINPUT54), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n800), .A2(new_n528), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n771), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n723), .A2(new_n662), .A3(new_n754), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT50), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n893), .A2(new_n822), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n819), .B(new_n820), .C1(new_n385), .C2(new_n753), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n891), .B(KEYINPUT50), .C1(new_n893), .C2(new_n894), .ZN(new_n901));
  INV_X1    g715(.A(new_n774), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n753), .A2(new_n386), .A3(new_n822), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n892), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n728), .A3(new_n238), .A4(new_n528), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT120), .Z(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n666), .A3(new_n676), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n897), .A2(new_n900), .A3(new_n901), .A4(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT51), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n906), .A2(new_n677), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n524), .B(new_n913), .C1(new_n893), .C2(new_n760), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n786), .A2(new_n790), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(new_n239), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n892), .A2(new_n916), .A3(new_n903), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n917), .A2(KEYINPUT48), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(KEYINPUT48), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n914), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n908), .B1(new_n899), .B2(new_n898), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n921), .A2(KEYINPUT51), .A3(new_n897), .A4(new_n901), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n912), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n855), .A2(new_n878), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n851), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n841), .A2(new_n876), .A3(new_n925), .ZN(new_n926));
  XOR2_X1   g740(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n927));
  NAND3_X1  g741(.A1(new_n886), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n890), .A2(new_n923), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(G952), .A2(G953), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n753), .B(KEYINPUT49), .Z(new_n931));
  NOR4_X1   g745(.A1(new_n239), .A2(new_n676), .A3(new_n386), .A4(new_n662), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n931), .A2(new_n723), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n666), .A2(new_n728), .ZN(new_n934));
  OAI22_X1  g748(.A1(new_n929), .A2(new_n930), .B1(new_n933), .B2(new_n934), .ZN(G75));
  NOR2_X1   g749(.A1(new_n223), .A2(G952), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n886), .A2(new_n926), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n230), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n939), .A2(new_n518), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n492), .B1(new_n496), .B2(new_n497), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(new_n480), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT55), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT56), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n937), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n188), .B1(new_n886), .B2(new_n926), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n517), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n943), .B1(new_n948), .B2(new_n944), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n946), .A2(new_n949), .ZN(G51));
  AND3_X1   g764(.A1(new_n886), .A2(new_n926), .A3(new_n927), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n927), .B1(new_n886), .B2(new_n926), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n464), .B(KEYINPUT57), .ZN(new_n954));
  OAI22_X1  g768(.A1(new_n953), .A2(new_n954), .B1(new_n461), .B2(new_n460), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n939), .A2(new_n810), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n936), .B1(new_n955), .B2(new_n956), .ZN(G54));
  NAND2_X1  g771(.A1(KEYINPUT58), .A2(G475), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n586), .B1(new_n939), .B2(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n947), .A2(KEYINPUT58), .A3(G475), .A4(new_n595), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n959), .A2(new_n937), .A3(new_n960), .ZN(G60));
  NAND2_X1  g775(.A1(G478), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT59), .Z(new_n963));
  NOR2_X1   g777(.A1(new_n672), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n951), .B2(new_n952), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n937), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n890), .A2(new_n928), .ZN(new_n967));
  INV_X1    g781(.A(new_n963), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n966), .B1(new_n969), .B2(new_n672), .ZN(G63));
  XNOR2_X1  g784(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  XNOR2_X1  g786(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n187), .A2(new_n513), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n886), .B2(new_n926), .ZN(new_n977));
  INV_X1    g791(.A(new_n229), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n937), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AOI211_X1 g793(.A(new_n698), .B(new_n976), .C1(new_n886), .C2(new_n926), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n972), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n938), .A2(new_n975), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n229), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n977), .A2(new_n697), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n983), .A2(new_n937), .A3(new_n984), .A4(new_n971), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n981), .A2(new_n985), .ZN(G66));
  OAI21_X1  g800(.A(G953), .B1(new_n530), .B2(new_n478), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n858), .B2(G953), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n941), .B1(G898), .B2(new_n223), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n988), .B(new_n989), .ZN(G69));
  NAND2_X1  g804(.A1(new_n382), .A2(new_n782), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n677), .B1(new_n666), .B2(new_n686), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n735), .B1(new_n992), .B2(KEYINPUT123), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(KEYINPUT123), .B2(new_n992), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n824), .B(new_n817), .C1(new_n991), .C2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n739), .A2(new_n747), .A3(new_n839), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n995), .B1(KEYINPUT62), .B2(new_n996), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n998));
  AOI21_X1  g812(.A(G953), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n363), .A2(new_n364), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n577), .A2(new_n578), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n795), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n824), .A2(new_n817), .A3(new_n1003), .A4(new_n797), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT126), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n916), .A2(new_n734), .A3(new_n815), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n764), .A2(new_n766), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n664), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1005), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1008), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n816), .A2(KEYINPUT126), .A3(new_n1010), .A4(new_n916), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n839), .A2(new_n747), .ZN(new_n1013));
  NOR4_X1   g827(.A1(new_n1004), .A2(new_n1012), .A3(G953), .A4(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1002), .B1(new_n717), .B2(new_n223), .ZN(new_n1015));
  OAI22_X1  g829(.A1(new_n999), .A2(new_n1002), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(G953), .B1(new_n450), .B2(new_n717), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(KEYINPUT125), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1018), .B1(new_n1019), .B2(KEYINPUT124), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1016), .B(new_n1020), .ZN(G72));
  NOR2_X1   g835(.A1(new_n347), .A2(new_n348), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1022), .B(KEYINPUT127), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n997), .A2(new_n858), .A3(new_n998), .ZN(new_n1024));
  NAND2_X1  g838(.A1(G472), .A2(G902), .ZN(new_n1025));
  XOR2_X1   g839(.A(new_n1025), .B(KEYINPUT63), .Z(new_n1026));
  AOI211_X1 g840(.A(new_n327), .B(new_n1023), .C1(new_n1024), .C2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n351), .A2(new_n352), .A3(new_n366), .ZN(new_n1028));
  AND4_X1   g842(.A1(new_n889), .A2(new_n887), .A3(new_n1028), .A4(new_n1026), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1026), .ZN(new_n1030));
  NOR3_X1   g844(.A1(new_n1004), .A2(new_n1013), .A3(new_n1012), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1030), .B1(new_n1031), .B2(new_n858), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1023), .A2(new_n327), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n937), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n1027), .A2(new_n1029), .A3(new_n1034), .ZN(G57));
endmodule


