//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1314, new_n1315,
    new_n1316, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n206), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n206), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT65), .Z(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n214), .A2(new_n217), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n213), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XOR2_X1   g0027(.A(KEYINPUT2), .B(G226), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n229), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(G107), .B(G116), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  AND2_X1   g0041(.A1(G33), .A2(G41), .ZN(new_n242));
  NOR2_X1   g0042(.A1(new_n242), .A2(new_n220), .ZN(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(G33), .A2(G97), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT3), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  AOI21_X1  g0050(.A(G1698), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n246), .B1(new_n251), .B2(G226), .ZN(new_n252));
  AND2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  OAI211_X1 g0054(.A(G232), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n244), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT67), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(new_n242), .B2(new_n220), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n262), .A2(KEYINPUT67), .A3(G1), .A4(G13), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n258), .A2(new_n261), .A3(G274), .A4(new_n263), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n258), .A2(G238), .A3(new_n260), .A4(new_n263), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT13), .B1(new_n256), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  OAI211_X1 g0068(.A(G226), .B(new_n268), .C1(new_n253), .C2(new_n254), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n255), .A2(new_n269), .A3(new_n245), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n243), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT13), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n271), .A2(new_n272), .A3(new_n264), .A4(new_n265), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n267), .A2(KEYINPUT75), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n266), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT75), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n275), .A2(new_n276), .A3(new_n272), .A4(new_n271), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n274), .A2(G169), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT14), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n273), .A2(G179), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n267), .A2(KEYINPUT76), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT76), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n282), .B(KEYINPUT13), .C1(new_n256), .C2(new_n266), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT79), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT14), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n274), .A2(new_n286), .A3(G169), .A4(new_n277), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT79), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n280), .A2(new_n281), .A3(new_n283), .A4(new_n288), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n279), .A2(new_n285), .A3(new_n287), .A4(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT77), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n221), .A2(G68), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT68), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(new_n248), .B2(G20), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n221), .A2(KEYINPUT68), .A3(G33), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G77), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n291), .B(new_n293), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n298), .B1(new_n295), .B2(new_n296), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT77), .B1(new_n300), .B2(new_n292), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G20), .A2(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G50), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n299), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n305), .A2(new_n220), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(KEYINPUT11), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT12), .B1(new_n309), .B2(G68), .ZN(new_n310));
  OR3_X1    g0110(.A1(new_n309), .A2(KEYINPUT12), .A3(G68), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n220), .A3(new_n305), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G68), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n259), .B2(G20), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n310), .A2(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n308), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT11), .B1(new_n304), .B2(new_n307), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n290), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n274), .A2(G200), .A3(new_n277), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n281), .A2(G190), .A3(new_n273), .A4(new_n283), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(new_n323), .A3(new_n319), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT78), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n322), .A2(new_n323), .A3(new_n319), .A4(KEYINPUT78), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n321), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n249), .A2(KEYINPUT7), .A3(new_n221), .A4(new_n250), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n253), .A2(new_n254), .A3(G20), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT7), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT80), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT80), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT7), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n330), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G68), .ZN(new_n338));
  AND2_X1   g0138(.A1(G58), .A2(G68), .ZN(new_n339));
  OAI21_X1  g0139(.A(G20), .B1(new_n339), .B2(new_n202), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n302), .A2(G159), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT16), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT81), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n249), .A2(new_n221), .A3(new_n250), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n314), .B1(new_n348), .B2(KEYINPUT7), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT80), .B(KEYINPUT7), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n331), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  AND4_X1   g0152(.A1(new_n347), .A2(new_n352), .A3(KEYINPUT16), .A4(new_n343), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n342), .B1(new_n349), .B2(new_n351), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n347), .B1(new_n354), .B2(KEYINPUT16), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n346), .B(new_n307), .C1(new_n353), .C2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G58), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT8), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT8), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G58), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n259), .A2(G20), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n363), .A2(new_n312), .B1(new_n361), .B2(new_n309), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G200), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n268), .B1(new_n249), .B2(new_n250), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n368));
  OAI211_X1 g0168(.A(G223), .B(new_n268), .C1(new_n253), .C2(new_n254), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n244), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n258), .A2(G232), .A3(new_n260), .A4(new_n263), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n264), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n366), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n264), .A2(new_n371), .ZN(new_n374));
  OAI211_X1 g0174(.A(G226), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n375));
  INV_X1    g0175(.A(G87), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n369), .B(new_n375), .C1(new_n248), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n243), .ZN(new_n378));
  INV_X1    g0178(.A(G190), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n374), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n373), .A2(new_n380), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n356), .A2(new_n365), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT17), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT82), .ZN(new_n384));
  INV_X1    g0184(.A(G179), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n374), .A2(new_n378), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n374), .A2(new_n378), .A3(new_n385), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT82), .ZN(new_n388));
  AOI21_X1  g0188(.A(G169), .B1(new_n374), .B2(new_n378), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n386), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n342), .B1(new_n337), .B2(G68), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n307), .B1(new_n391), .B2(KEYINPUT16), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n354), .A2(new_n347), .A3(KEYINPUT16), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n352), .A2(KEYINPUT16), .A3(new_n343), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT81), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n392), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n390), .B1(new_n396), .B2(new_n364), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT18), .ZN(new_n398));
  INV_X1    g0198(.A(G169), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n370), .B2(new_n372), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n400), .A2(KEYINPUT82), .A3(new_n387), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n356), .A2(new_n365), .B1(new_n401), .B2(new_n386), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT18), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n356), .A2(new_n365), .A3(new_n381), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT17), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n383), .A2(new_n398), .A3(new_n404), .A4(new_n407), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n258), .A2(new_n263), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(G226), .A3(new_n260), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n253), .A2(new_n254), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n367), .A2(G223), .B1(new_n411), .B2(G77), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n251), .A2(G222), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n264), .B(new_n410), .C1(new_n414), .C2(new_n244), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n399), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(G179), .B2(new_n415), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n295), .A2(new_n296), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n418), .A2(new_n361), .B1(G150), .B2(new_n302), .ZN(new_n419));
  OR2_X1    g0219(.A1(new_n419), .A2(KEYINPUT69), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n419), .A2(KEYINPUT69), .B1(G20), .B2(new_n203), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n306), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n362), .A2(G50), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n312), .A2(new_n423), .B1(G50), .B2(new_n309), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n362), .A2(G77), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n312), .A2(new_n427), .B1(G77), .B2(new_n309), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n221), .A2(new_n248), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n429), .A2(KEYINPUT70), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(KEYINPUT70), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(new_n361), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT71), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT15), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(G87), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n376), .A2(KEYINPUT15), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n433), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n376), .A2(KEYINPUT15), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(G87), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT71), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  OAI221_X1 g0241(.A(new_n432), .B1(new_n221), .B2(new_n298), .C1(new_n441), .C2(new_n297), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n428), .B1(new_n442), .B2(new_n307), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT72), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n409), .A2(G244), .A3(new_n260), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n264), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n367), .A2(G238), .B1(new_n411), .B2(G107), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n249), .A2(new_n250), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(G232), .A3(new_n268), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n244), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n399), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n444), .A2(new_n445), .A3(new_n452), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n446), .A2(new_n264), .ZN(new_n454));
  INV_X1    g0254(.A(new_n451), .ZN(new_n455));
  AOI21_X1  g0255(.A(G169), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT72), .B1(new_n456), .B2(new_n443), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n447), .A2(new_n451), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n385), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n453), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(G190), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n461), .B(new_n443), .C1(new_n366), .C2(new_n458), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n426), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n329), .A2(new_n408), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT10), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n425), .A2(KEYINPUT73), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT73), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n422), .B2(new_n424), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(KEYINPUT9), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT74), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT74), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n466), .A2(new_n471), .A3(KEYINPUT9), .A4(new_n468), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n415), .A2(G200), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n379), .B2(new_n415), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n466), .A2(new_n468), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT9), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n465), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n473), .A2(new_n478), .A3(new_n465), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n464), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G116), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n305), .A2(new_n220), .B1(G20), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  INV_X1    g0285(.A(G97), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n485), .B(new_n221), .C1(G33), .C2(new_n486), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n484), .A2(KEYINPUT20), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT20), .B1(new_n484), .B2(new_n487), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n309), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(G116), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT84), .B1(new_n248), .B2(G1), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT84), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(new_n259), .A3(G33), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(new_n306), .A3(new_n309), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n492), .B1(new_n497), .B2(G116), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT92), .B1(new_n490), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n493), .A2(new_n495), .ZN(new_n500));
  OAI21_X1  g0300(.A(G116), .B1(new_n500), .B2(new_n312), .ZN(new_n501));
  INV_X1    g0301(.A(new_n492), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT92), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n484), .A2(new_n487), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT20), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n484), .A2(KEYINPUT20), .A3(new_n487), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n503), .A2(new_n504), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n499), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT91), .ZN(new_n512));
  INV_X1    g0312(.A(G45), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(G1), .ZN(new_n514));
  NAND2_X1  g0314(.A1(KEYINPUT5), .A2(G41), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(KEYINPUT5), .A2(G41), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n409), .A2(new_n512), .A3(G270), .A4(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(G264), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n520));
  OAI211_X1 g0320(.A(G257), .B(new_n268), .C1(new_n253), .C2(new_n254), .ZN(new_n521));
  INV_X1    g0321(.A(G303), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n520), .B(new_n521), .C1(new_n522), .C2(new_n449), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n243), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n259), .A2(G45), .ZN(new_n525));
  OR2_X1    g0325(.A1(KEYINPUT5), .A2(G41), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n525), .B1(new_n526), .B2(new_n515), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n527), .A2(G274), .A3(new_n258), .A4(new_n263), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n518), .A2(new_n258), .A3(G270), .A4(new_n263), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT91), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n519), .A2(new_n524), .A3(new_n528), .A4(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n511), .A2(KEYINPUT21), .A3(G169), .A4(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n531), .A2(new_n385), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n511), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n531), .A2(G169), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT21), .B1(new_n537), .B2(new_n511), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n518), .A2(new_n258), .A3(new_n263), .ZN(new_n540));
  OAI211_X1 g0340(.A(G257), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n541));
  OAI211_X1 g0341(.A(G250), .B(new_n268), .C1(new_n253), .C2(new_n254), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G294), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n540), .A2(G264), .B1(new_n544), .B2(new_n243), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n545), .A2(G179), .A3(new_n528), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n243), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n518), .A2(new_n258), .A3(G264), .A4(new_n263), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n528), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G169), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n221), .B(G87), .C1(new_n253), .C2(new_n254), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT22), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT22), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n449), .A2(new_n554), .A3(new_n221), .A4(G87), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT24), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G116), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(G20), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT23), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n221), .B2(G107), .ZN(new_n561));
  INV_X1    g0361(.A(G107), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n562), .A2(KEYINPUT23), .A3(G20), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n559), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n556), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n557), .B1(new_n556), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n307), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n309), .A2(G107), .ZN(new_n568));
  XOR2_X1   g0368(.A(new_n568), .B(KEYINPUT25), .Z(new_n569));
  INV_X1    g0369(.A(new_n497), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n569), .B1(G107), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n551), .A2(KEYINPUT94), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT94), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n546), .A2(new_n550), .A3(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n567), .A2(new_n571), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n545), .A2(KEYINPUT95), .A3(new_n379), .A4(new_n528), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT95), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(new_n549), .B2(new_n366), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n549), .A2(G190), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n572), .A2(new_n574), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(G244), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n582));
  OAI211_X1 g0382(.A(G238), .B(new_n268), .C1(new_n253), .C2(new_n254), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n558), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n243), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT89), .ZN(new_n586));
  AOI21_X1  g0386(.A(G250), .B1(new_n259), .B2(G45), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(G274), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n514), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n258), .A2(new_n588), .A3(new_n590), .A4(new_n263), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n585), .A2(new_n586), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n586), .B1(new_n585), .B2(new_n591), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n385), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n585), .A2(new_n591), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT89), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n585), .A2(new_n586), .A3(new_n591), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n399), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n309), .B1(new_n437), .B2(new_n440), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n221), .B(G68), .C1(new_n253), .C2(new_n254), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT19), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n221), .B1(new_n245), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n376), .A2(new_n486), .A3(new_n562), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n486), .B1(new_n295), .B2(new_n296), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n600), .B(new_n604), .C1(new_n605), .C2(KEYINPUT19), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n599), .B1(new_n606), .B2(new_n307), .ZN(new_n607));
  INV_X1    g0407(.A(new_n441), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n570), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT90), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT90), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n607), .A2(new_n612), .A3(new_n609), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n594), .A2(new_n598), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(G190), .B1(new_n592), .B2(new_n593), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n596), .A2(G200), .A3(new_n597), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n570), .A2(G87), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n607), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n615), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT93), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n531), .A2(G200), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n621), .B1(new_n623), .B2(new_n511), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n499), .A2(new_n510), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(KEYINPUT93), .A3(new_n622), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n531), .A2(new_n379), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n539), .A2(new_n581), .A3(new_n620), .A4(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(KEYINPUT4), .A2(G244), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n268), .B(new_n630), .C1(new_n253), .C2(new_n254), .ZN(new_n631));
  INV_X1    g0431(.A(G244), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n249), .B2(new_n250), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n631), .B(new_n485), .C1(new_n633), .C2(KEYINPUT4), .ZN(new_n634));
  OAI21_X1  g0434(.A(G250), .B1(new_n253), .B2(new_n254), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n268), .B1(new_n635), .B2(KEYINPUT4), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n243), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n518), .A2(new_n258), .A3(G257), .A4(new_n263), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n528), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n399), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT85), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n528), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n642), .B1(new_n528), .B2(new_n638), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n385), .B(new_n637), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n302), .A2(G77), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT6), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n647), .A2(new_n486), .A3(G107), .ZN(new_n648));
  XNOR2_X1  g0448(.A(G97), .B(G107), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n646), .B1(new_n650), .B2(new_n221), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n348), .A2(new_n350), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n562), .B1(new_n652), .B2(new_n330), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n307), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT83), .B1(new_n309), .B2(G97), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT83), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n491), .A2(new_n656), .A3(new_n486), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n570), .A2(G97), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n641), .A2(new_n645), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT87), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n637), .B1(new_n643), .B2(new_n644), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G200), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT86), .B1(new_n640), .B2(new_n379), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n654), .A2(new_n658), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT86), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n637), .A2(new_n639), .A3(new_n666), .A4(G190), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n663), .A2(new_n664), .A3(new_n665), .A4(new_n667), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n399), .A2(new_n640), .B1(new_n654), .B2(new_n658), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT87), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(new_n670), .A3(new_n645), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n661), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT88), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n661), .A2(new_n668), .A3(new_n671), .A4(KEYINPUT88), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n482), .A2(new_n629), .A3(new_n676), .ZN(G372));
  INV_X1    g0477(.A(new_n426), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT97), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n481), .B2(new_n479), .ZN(new_n680));
  INV_X1    g0480(.A(new_n479), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n681), .A2(KEYINPUT97), .A3(new_n480), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n356), .A2(new_n365), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n684), .A2(new_n403), .A3(new_n390), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n403), .B1(new_n684), .B2(new_n390), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n460), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n328), .A2(new_n688), .B1(new_n320), .B2(new_n290), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n405), .B(KEYINPUT17), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n687), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n678), .B1(new_n683), .B2(new_n692), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n641), .A2(new_n645), .A3(new_n659), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT96), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n591), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n587), .B1(new_n589), .B2(new_n514), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n697), .A2(KEYINPUT96), .A3(new_n258), .A4(new_n263), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n585), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G200), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n615), .A2(new_n618), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT26), .ZN(new_n702));
  AOI22_X1  g0502(.A1(new_n399), .A2(new_n699), .B1(new_n607), .B2(new_n609), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n594), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n694), .A2(new_n701), .A3(new_n702), .A4(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n704), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n660), .A2(KEYINPUT87), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n670), .B1(new_n669), .B2(new_n645), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n619), .B(new_n614), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n706), .B1(KEYINPUT26), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n672), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n575), .A2(new_n580), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT21), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n625), .B2(new_n536), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n567), .A2(new_n571), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n551), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n714), .A2(new_n716), .A3(new_n534), .A4(new_n532), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n701), .A2(new_n704), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n711), .A2(new_n712), .A3(new_n717), .A4(new_n719), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n710), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n693), .B1(new_n482), .B2(new_n721), .ZN(G369));
  NAND3_X1  g0522(.A1(new_n714), .A2(new_n534), .A3(new_n532), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n259), .A2(new_n221), .A3(G13), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(KEYINPUT27), .ZN(new_n725));
  XOR2_X1   g0525(.A(new_n725), .B(KEYINPUT98), .Z(new_n726));
  INV_X1    g0526(.A(G213), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(new_n724), .B2(KEYINPUT27), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(G343), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n723), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n581), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n715), .A2(new_n551), .A3(new_n732), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT99), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n732), .A2(new_n625), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n539), .A2(new_n628), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(new_n539), .B2(new_n741), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G330), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n581), .B1(new_n575), .B2(new_n732), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n572), .A2(new_n574), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n746), .B1(new_n747), .B2(new_n732), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n739), .A2(new_n749), .ZN(G399));
  INV_X1    g0550(.A(new_n215), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G41), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n603), .A2(G116), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n753), .A2(G1), .A3(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n219), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n755), .B1(new_n756), .B2(new_n753), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT28), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n721), .A2(KEYINPUT29), .A3(new_n731), .ZN(new_n759));
  INV_X1    g0559(.A(new_n712), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n672), .A2(new_n760), .A3(new_n718), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT103), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(new_n539), .B2(new_n747), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n399), .B1(new_n545), .B2(new_n528), .ZN(new_n764));
  AND4_X1   g0564(.A1(G179), .A2(new_n547), .A3(new_n528), .A4(new_n548), .ZN(new_n765));
  OAI21_X1  g0565(.A(KEYINPUT94), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AND3_X1   g0566(.A1(new_n766), .A2(new_n715), .A3(new_n574), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n723), .A2(new_n767), .A3(KEYINPUT103), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n761), .B1(new_n763), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(KEYINPUT104), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT104), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n761), .B(new_n771), .C1(new_n763), .C2(new_n768), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n661), .A2(new_n671), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n620), .A2(new_n702), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(KEYINPUT26), .B1(new_n718), .B2(new_n660), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n774), .A2(new_n704), .A3(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT102), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n774), .A2(KEYINPUT102), .A3(new_n704), .A4(new_n775), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n770), .A2(new_n772), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n732), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n759), .B1(new_n781), .B2(KEYINPUT29), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n674), .A2(new_n675), .ZN(new_n783));
  AND4_X1   g0583(.A1(new_n581), .A2(new_n539), .A3(new_n620), .A4(new_n628), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n783), .A2(new_n784), .A3(new_n732), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n596), .A2(new_n597), .ZN(new_n786));
  AND3_X1   g0586(.A1(new_n545), .A2(new_n637), .A3(new_n639), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n533), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT30), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n533), .A2(new_n786), .A3(new_n787), .A4(KEYINPUT30), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT100), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n662), .A2(new_n792), .A3(new_n549), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n792), .B1(new_n662), .B2(new_n549), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n531), .A2(new_n385), .A3(new_n699), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n790), .B(new_n791), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n798), .A2(KEYINPUT101), .A3(KEYINPUT31), .A4(new_n731), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n790), .A2(new_n791), .ZN(new_n800));
  INV_X1    g0600(.A(new_n795), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n797), .B1(new_n801), .B2(new_n793), .ZN(new_n802));
  OAI211_X1 g0602(.A(KEYINPUT31), .B(new_n731), .C1(new_n800), .C2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT101), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n731), .B1(new_n800), .B2(new_n802), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT31), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n785), .A2(new_n799), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G330), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n782), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n758), .B1(new_n811), .B2(G1), .ZN(G364));
  OAI21_X1  g0612(.A(G20), .B1(KEYINPUT107), .B2(G169), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(KEYINPUT107), .A2(G169), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n220), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n221), .A2(G179), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n818), .A2(G190), .A3(G200), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n376), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G190), .A2(G200), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G159), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(KEYINPUT32), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n221), .A2(new_n385), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(G200), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(G190), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n820), .B(new_n825), .C1(G68), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n826), .A2(new_n821), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n449), .B1(new_n830), .B2(new_n298), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n826), .A2(G190), .A3(new_n366), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n831), .B1(G58), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n818), .A2(new_n379), .A3(G200), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n562), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n824), .B2(KEYINPUT32), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n379), .A2(G179), .A3(G200), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(new_n221), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n827), .A2(new_n379), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G97), .A2(new_n840), .B1(new_n841), .B2(G50), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n829), .A2(new_n834), .A3(new_n837), .A4(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(G322), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n832), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(G311), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n411), .B1(new_n830), .B2(new_n846), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n845), .B(new_n847), .C1(G329), .C2(new_n823), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n841), .A2(G326), .ZN(new_n849));
  XNOR2_X1  g0649(.A(KEYINPUT33), .B(G317), .ZN(new_n850));
  INV_X1    g0650(.A(new_n819), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n828), .A2(new_n850), .B1(new_n851), .B2(G303), .ZN(new_n852));
  INV_X1    g0652(.A(new_n835), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n840), .A2(G294), .B1(new_n853), .B2(G283), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n848), .A2(new_n849), .A3(new_n852), .A4(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n817), .B1(new_n843), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(G13), .A2(G33), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n221), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT106), .Z(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n817), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n411), .A2(new_n215), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT105), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n219), .A2(new_n513), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n862), .B(new_n863), .C1(new_n513), .C2(new_n240), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n751), .A2(new_n411), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n865), .A2(G355), .B1(new_n483), .B2(new_n751), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n860), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(G13), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n868), .A2(G20), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n259), .B1(new_n869), .B2(G45), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n752), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n856), .A2(new_n867), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n743), .B2(new_n859), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n744), .A2(new_n873), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n743), .A2(G330), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT108), .Z(G396));
  AOI21_X1  g0679(.A(new_n731), .B1(new_n710), .B2(new_n720), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT109), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n732), .A2(new_n443), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n460), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n457), .A2(new_n459), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n462), .B1(new_n885), .B2(new_n453), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n882), .B1(new_n460), .B2(new_n881), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n880), .B(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n872), .B1(new_n889), .B2(new_n810), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n810), .B2(new_n889), .ZN(new_n891));
  INV_X1    g0691(.A(new_n841), .ZN(new_n892));
  OAI22_X1  g0692(.A1(new_n892), .A2(new_n522), .B1(new_n819), .B2(new_n562), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(G87), .B2(new_n853), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n449), .B1(new_n833), .B2(G294), .ZN(new_n895));
  INV_X1    g0695(.A(new_n830), .ZN(new_n896));
  AOI22_X1  g0696(.A1(G116), .A2(new_n896), .B1(new_n823), .B2(G311), .ZN(new_n897));
  AOI22_X1  g0697(.A1(G97), .A2(new_n840), .B1(new_n828), .B2(G283), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n894), .A2(new_n895), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n833), .A2(G143), .B1(new_n896), .B2(G159), .ZN(new_n900));
  INV_X1    g0700(.A(new_n828), .ZN(new_n901));
  INV_X1    g0701(.A(G150), .ZN(new_n902));
  INV_X1    g0702(.A(G137), .ZN(new_n903));
  OAI221_X1 g0703(.A(new_n900), .B1(new_n901), .B2(new_n902), .C1(new_n903), .C2(new_n892), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT34), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n835), .A2(new_n314), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n411), .B(new_n907), .C1(G132), .C2(new_n823), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n840), .A2(G58), .B1(new_n851), .B2(G50), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n904), .A2(new_n905), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n899), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n816), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n816), .A2(new_n857), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n873), .B1(new_n914), .B2(new_n298), .ZN(new_n915));
  INV_X1    g0715(.A(new_n857), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n913), .B(new_n915), .C1(new_n888), .C2(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n891), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(G384));
  INV_X1    g0719(.A(new_n650), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n920), .A2(KEYINPUT35), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(KEYINPUT35), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n921), .A2(G116), .A3(new_n222), .A4(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT36), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n756), .A2(new_n298), .A3(new_n339), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n925), .A2(KEYINPUT110), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(KEYINPUT110), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n201), .A2(G68), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT111), .ZN(new_n929));
  NOR3_X1   g0729(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n868), .A2(G1), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n676), .A2(new_n629), .A3(new_n731), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n808), .A2(new_n803), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n320), .A2(new_n731), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n321), .A2(new_n328), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n935), .B1(new_n321), .B2(new_n328), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n888), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT113), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n460), .A2(new_n881), .ZN(new_n940));
  INV_X1    g0740(.A(new_n882), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n942), .B(new_n883), .C1(new_n688), .C2(new_n462), .ZN(new_n943));
  INV_X1    g0743(.A(new_n935), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n329), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n321), .A2(new_n328), .A3(new_n935), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n785), .A2(new_n803), .A3(new_n808), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT40), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT113), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n947), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n729), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n353), .A2(new_n355), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n307), .B1(new_n354), .B2(KEYINPUT16), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n365), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n408), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n952), .B1(new_n396), .B2(new_n364), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT37), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n397), .A2(new_n957), .A3(new_n958), .A4(new_n405), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT112), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n395), .A2(new_n393), .ZN(new_n961));
  INV_X1    g0761(.A(new_n392), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n364), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n955), .A2(new_n952), .B1(new_n963), .B2(new_n381), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n955), .A2(new_n390), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n958), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI211_X1 g0766(.A(KEYINPUT38), .B(new_n956), .C1(new_n960), .C2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT38), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n382), .A2(new_n402), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n969), .A2(KEYINPUT112), .A3(new_n958), .A4(new_n957), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT112), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n959), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n966), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n955), .A2(new_n952), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n687), .B2(new_n690), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n968), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n967), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n939), .A2(new_n951), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n934), .A2(new_n938), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n969), .A2(new_n957), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n970), .A2(new_n972), .B1(new_n980), .B2(KEYINPUT37), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n957), .B1(new_n687), .B2(new_n690), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n968), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n967), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n978), .B1(new_n985), .B2(new_n949), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n482), .A2(new_n934), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n986), .A2(new_n987), .ZN(new_n989));
  INV_X1    g0789(.A(G330), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n693), .B1(new_n782), .B2(new_n482), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT39), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n980), .A2(KEYINPUT37), .ZN(new_n994));
  INV_X1    g0794(.A(new_n972), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n959), .A2(new_n971), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n982), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT38), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n973), .A2(new_n968), .A3(new_n975), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n993), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n290), .A2(new_n320), .A3(new_n732), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n967), .A2(new_n976), .A3(KEYINPUT39), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1001), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n687), .A2(new_n952), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n936), .A2(new_n937), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n880), .A2(new_n888), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n460), .A2(new_n731), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1007), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1006), .B1(new_n1011), .B2(new_n977), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n1005), .A2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n992), .B(new_n1013), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n991), .A2(new_n1014), .B1(new_n259), .B2(new_n869), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n991), .A2(new_n1014), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n924), .B1(new_n930), .B2(new_n931), .C1(new_n1015), .C2(new_n1016), .ZN(G367));
  INV_X1    g0817(.A(new_n862), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n233), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n860), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n215), .B2(new_n441), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n872), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G143), .A2(new_n841), .B1(new_n828), .B2(G159), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n411), .B1(new_n833), .B2(G150), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n201), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n1025), .A2(new_n896), .B1(new_n823), .B2(G137), .ZN(new_n1026));
  AND3_X1   g0826(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n851), .A2(G58), .B1(new_n853), .B2(G77), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(new_n314), .C2(new_n839), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n828), .A2(G294), .B1(new_n853), .B2(G97), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n562), .B2(new_n839), .C1(new_n846), .C2(new_n892), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n833), .A2(G303), .B1(new_n823), .B2(G317), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT46), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n819), .B2(new_n483), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n851), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n449), .B1(new_n896), .B2(G283), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1029), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT47), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1022), .B1(new_n1039), .B2(new_n816), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n732), .A2(new_n618), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1041), .A2(new_n594), .A3(new_n703), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n718), .B2(new_n1041), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1040), .B1(new_n1043), .B2(new_n859), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n749), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n737), .B(KEYINPUT99), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n711), .B1(new_n665), .B2(new_n732), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n694), .A2(new_n731), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT44), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1049), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n739), .A2(new_n1052), .ZN(new_n1053));
  XOR2_X1   g0853(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1053), .B(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1045), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n735), .B1(new_n748), .B2(new_n734), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n744), .B2(KEYINPUT116), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n744), .A2(KEYINPUT116), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1059), .B(new_n1060), .Z(new_n1061));
  AND2_X1   g0861(.A1(new_n811), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT44), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1050), .B(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1053), .B(new_n1054), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1064), .A2(new_n1065), .A3(new_n749), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1057), .A2(new_n1062), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n811), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n752), .B(KEYINPUT41), .Z(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n871), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1049), .A2(new_n735), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT42), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1049), .A2(new_n747), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n732), .B1(new_n1074), .B2(new_n773), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  OR3_X1    g0876(.A1(new_n1076), .A2(KEYINPUT43), .A3(new_n1043), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1043), .B(KEYINPUT43), .Z(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT114), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1076), .A2(KEYINPUT114), .A3(new_n1078), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1077), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1045), .A2(new_n1052), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1083), .B(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1044), .B1(new_n1071), .B2(new_n1085), .ZN(G387));
  OR2_X1    g0886(.A1(new_n748), .A2(new_n859), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n754), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n865), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(G107), .B2(new_n215), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n229), .A2(new_n513), .ZN(new_n1091));
  INV_X1    g0891(.A(G50), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n361), .A2(new_n1092), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT50), .Z(new_n1094));
  AOI211_X1 g0894(.A(G45), .B(new_n1088), .C1(G68), .C2(G77), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1018), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1090), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n872), .B1(new_n1097), .B2(new_n860), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n832), .A2(new_n1092), .B1(new_n822), .B2(new_n902), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n411), .B(new_n1099), .C1(G68), .C2(new_n896), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n819), .A2(new_n298), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G97), .B2(new_n853), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G159), .A2(new_n841), .B1(new_n828), .B2(new_n361), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n608), .A2(new_n840), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1100), .A2(new_n1102), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n449), .B1(new_n823), .B2(G326), .ZN(new_n1106));
  INV_X1    g0906(.A(G283), .ZN(new_n1107));
  INV_X1    g0907(.A(G294), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n839), .A2(new_n1107), .B1(new_n819), .B2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n833), .A2(G317), .B1(new_n896), .B2(G303), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1110), .B1(new_n901), .B2(new_n846), .C1(new_n844), .C2(new_n892), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT48), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1109), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1112), .B2(new_n1111), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT49), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1106), .B1(new_n483), .B2(new_n835), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1105), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1098), .B1(new_n1118), .B2(new_n816), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1061), .A2(new_n871), .B1(new_n1087), .B2(new_n1119), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1062), .A2(new_n753), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n811), .A2(new_n1061), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(G393));
  NAND3_X1  g0923(.A1(new_n1057), .A2(new_n871), .A3(new_n1066), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1020), .B1(new_n486), .B2(new_n215), .C1(new_n1018), .C2(new_n237), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n872), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G150), .A2(new_n841), .B1(new_n833), .B2(G159), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1127), .B(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n411), .B1(new_n823), .B2(G143), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n361), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n830), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n828), .A2(new_n1025), .B1(new_n853), .B2(G87), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n839), .A2(new_n298), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G68), .B2(new_n851), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1129), .A2(new_n1133), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G317), .A2(new_n841), .B1(new_n833), .B2(G311), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT52), .Z(new_n1139));
  OAI21_X1  g0939(.A(new_n411), .B1(new_n822), .B2(new_n844), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n836), .B(new_n1140), .C1(G283), .C2(new_n851), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n840), .A2(G116), .B1(new_n896), .B2(G294), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n522), .B2(new_n901), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT118), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1137), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1126), .B1(new_n1146), .B2(new_n816), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n1052), .B2(new_n859), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1067), .A2(new_n752), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1062), .B1(new_n1057), .B2(new_n1066), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1124), .B(new_n1148), .C1(new_n1149), .C2(new_n1150), .ZN(G390));
  NAND2_X1  g0951(.A1(new_n984), .A2(new_n1002), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n780), .A2(new_n732), .A3(new_n888), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1010), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1007), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1152), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1009), .B1(new_n880), .B2(new_n888), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1002), .B1(new_n1157), .B2(new_n1007), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n967), .A2(new_n976), .A3(KEYINPUT39), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT39), .B1(new_n983), .B2(new_n967), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n809), .A2(new_n947), .A3(G330), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT119), .B1(new_n1156), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1162), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n1158), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT119), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1007), .B1(new_n1153), .B2(new_n1010), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1167), .B(new_n1168), .C1(new_n1169), .C2(new_n1152), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1164), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1161), .B1(new_n1169), .B2(new_n1152), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n979), .A2(G330), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1171), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n948), .A2(G330), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1177), .A2(new_n482), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n693), .B(new_n1178), .C1(new_n782), .C2(new_n482), .ZN(new_n1179));
  OAI211_X1 g0979(.A(G330), .B(new_n888), .C1(new_n932), .C2(new_n933), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n1007), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n1162), .ZN(new_n1182));
  OAI21_X1  g0982(.A(KEYINPUT120), .B1(new_n1154), .B2(new_n1182), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n805), .A2(new_n799), .A3(new_n808), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n990), .B1(new_n1184), .B2(new_n785), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1185), .A2(new_n947), .B1(new_n1180), .B2(new_n1007), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT120), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1186), .A2(new_n1187), .A3(new_n1010), .A4(new_n1153), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1183), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1007), .B1(new_n810), .B2(new_n943), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n1173), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1157), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1179), .B1(new_n1189), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n753), .B1(new_n1176), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1171), .A2(new_n1194), .A3(new_n1175), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1164), .A2(new_n1170), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n871), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1166), .A2(new_n857), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n873), .B1(new_n914), .B2(new_n1131), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G159), .A2(new_n840), .B1(new_n841), .B2(G128), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n903), .B2(new_n901), .C1(new_n201), .C2(new_n835), .ZN(new_n1204));
  INV_X1    g1004(.A(G125), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n449), .B1(new_n822), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(G132), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(KEYINPUT54), .B(G143), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n832), .A2(new_n1207), .B1(new_n830), .B2(new_n1208), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1204), .A2(new_n1206), .A3(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n819), .A2(new_n902), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT53), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n901), .A2(new_n562), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1135), .B(new_n1213), .C1(G283), .C2(new_n841), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n411), .B1(new_n832), .B2(new_n483), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n830), .A2(new_n486), .B1(new_n822), .B2(new_n1108), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1215), .A2(new_n1216), .A3(new_n820), .A4(new_n907), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1210), .A2(new_n1212), .B1(new_n1214), .B2(new_n1217), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1201), .B(new_n1202), .C1(new_n817), .C2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1198), .A2(new_n1200), .A3(new_n1219), .ZN(G378));
  INV_X1    g1020(.A(KEYINPUT57), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1179), .B1(new_n1199), .B2(new_n1194), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n939), .A2(new_n977), .A3(new_n951), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n949), .B1(new_n979), .B2(new_n984), .ZN(new_n1224));
  OAI21_X1  g1024(.A(G330), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n1013), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n680), .A2(new_n682), .A3(new_n426), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n476), .A2(new_n952), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n680), .A2(new_n682), .A3(new_n426), .A4(new_n1228), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1232), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT121), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1005), .A2(new_n1012), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n986), .A2(new_n1237), .A3(G330), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1226), .A2(new_n1236), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1236), .B1(new_n1226), .B2(new_n1238), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1221), .B1(new_n1222), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1179), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1197), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1226), .A2(new_n1238), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1236), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1226), .A2(new_n1236), .A3(new_n1238), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1244), .A2(KEYINPUT57), .A3(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1242), .A2(new_n1250), .A3(new_n752), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n1233), .A2(new_n1234), .A3(new_n916), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n449), .A2(G41), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1253), .B1(new_n1107), .B2(new_n822), .C1(new_n562), .C2(new_n832), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1101), .B(new_n1254), .C1(G68), .C2(new_n840), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n892), .A2(new_n483), .B1(new_n835), .B2(new_n357), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(G97), .B2(new_n828), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1255), .B(new_n1257), .C1(new_n441), .C2(new_n830), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT58), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1253), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1261), .B(new_n1092), .C1(G33), .C2(G41), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n901), .A2(new_n1207), .B1(new_n892), .B2(new_n1205), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n833), .A2(G128), .B1(new_n896), .B2(G137), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n819), .B2(new_n1208), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1264), .B(new_n1266), .C1(G150), .C2(new_n840), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT59), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n853), .A2(G159), .ZN(new_n1270));
  AOI211_X1 g1070(.A(G33), .B(G41), .C1(new_n823), .C2(G124), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1268), .A2(KEYINPUT59), .ZN(new_n1273));
  OAI221_X1 g1073(.A(new_n1263), .B1(new_n1259), .B2(new_n1258), .C1(new_n1272), .C2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n816), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n914), .A2(new_n201), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1275), .A2(new_n872), .A3(new_n1276), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n1241), .A2(new_n870), .B1(new_n1252), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1251), .A2(new_n1279), .ZN(G375));
  AOI22_X1  g1080(.A1(new_n1183), .A2(new_n1188), .B1(new_n1192), .B2(new_n1191), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1179), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1069), .B(KEYINPUT122), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1195), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1155), .A2(new_n916), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n892), .A2(new_n1207), .B1(new_n1092), .B2(new_n839), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(G159), .B2(new_n851), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n832), .A2(new_n903), .B1(new_n830), .B2(new_n902), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n411), .B(new_n1288), .C1(G128), .C2(new_n823), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1208), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n828), .A2(new_n1290), .B1(new_n853), .B2(G58), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1287), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1292));
  OAI22_X1  g1092(.A1(new_n901), .A2(new_n483), .B1(new_n486), .B2(new_n819), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1293), .B1(G294), .B2(new_n841), .ZN(new_n1294));
  OAI22_X1  g1094(.A1(new_n830), .A2(new_n562), .B1(new_n822), .B2(new_n522), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(G283), .B2(new_n833), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1294), .A2(new_n1104), .A3(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n411), .B1(new_n835), .B2(new_n298), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1298), .B(KEYINPUT123), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1292), .B1(new_n1297), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT124), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n817), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1302), .B1(new_n1301), .B2(new_n1300), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n914), .A2(new_n314), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n872), .A3(new_n1304), .ZN(new_n1305));
  OAI22_X1  g1105(.A1(new_n1281), .A2(new_n870), .B1(new_n1285), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1284), .A2(new_n1307), .ZN(G381));
  OR4_X1    g1108(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1200), .A2(new_n1219), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1310), .B1(new_n1197), .B2(new_n1196), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1251), .A2(new_n1311), .A3(new_n1279), .ZN(new_n1312));
  OR4_X1    g1112(.A1(G387), .A2(new_n1309), .A3(new_n1312), .A4(G381), .ZN(G407));
  NAND2_X1  g1113(.A1(new_n730), .A2(G213), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(new_n1314), .B(KEYINPUT125), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  OAI211_X1 g1116(.A(G407), .B(G213), .C1(new_n1312), .C2(new_n1316), .ZN(G409));
  INV_X1    g1117(.A(G390), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(G387), .A2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(G390), .B(new_n1044), .C1(new_n1071), .C2(new_n1085), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  XOR2_X1   g1121(.A(G393), .B(G396), .Z(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1322), .A2(new_n1319), .A3(new_n1320), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1326), .A2(KEYINPUT61), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1251), .A2(G378), .A3(new_n1279), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1244), .A2(new_n1249), .A3(new_n1283), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1311), .B1(new_n1329), .B2(new_n1278), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1189), .A2(new_n1193), .A3(KEYINPUT60), .A4(new_n1179), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n752), .ZN(new_n1333));
  OAI21_X1  g1133(.A(KEYINPUT60), .B1(new_n1281), .B2(new_n1179), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1333), .B1(new_n1282), .B2(new_n1334), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n918), .B1(new_n1335), .B2(new_n1306), .ZN(new_n1336));
  AND2_X1   g1136(.A1(new_n1334), .A2(new_n1282), .ZN(new_n1337));
  OAI211_X1 g1137(.A(G384), .B(new_n1307), .C1(new_n1337), .C2(new_n1333), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1336), .A2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1331), .A2(new_n1314), .A3(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT63), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1331), .A2(new_n1314), .ZN(new_n1344));
  AOI22_X1  g1144(.A1(new_n1336), .A2(new_n1338), .B1(G2897), .B2(new_n1315), .ZN(new_n1345));
  INV_X1    g1145(.A(G2897), .ZN(new_n1346));
  NOR3_X1   g1146(.A1(new_n1339), .A2(new_n1346), .A3(new_n1314), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1344), .B1(new_n1345), .B2(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1315), .B1(new_n1328), .B2(new_n1330), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1349), .A2(KEYINPUT63), .A3(new_n1340), .ZN(new_n1350));
  NAND4_X1  g1150(.A1(new_n1327), .A2(new_n1343), .A3(new_n1348), .A4(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT61), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1347), .A2(new_n1345), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1352), .B1(new_n1353), .B2(new_n1349), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1336), .A2(KEYINPUT62), .A3(new_n1338), .ZN(new_n1355));
  AOI211_X1 g1155(.A(new_n1315), .B(new_n1355), .C1(new_n1328), .C2(new_n1330), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT62), .ZN(new_n1357));
  AOI22_X1  g1157(.A1(KEYINPUT126), .A2(new_n1356), .B1(new_n1341), .B2(new_n1357), .ZN(new_n1358));
  OR2_X1    g1158(.A1(new_n1356), .A2(KEYINPUT126), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1354), .B1(new_n1358), .B2(new_n1359), .ZN(new_n1360));
  AND3_X1   g1160(.A1(new_n1322), .A2(new_n1319), .A3(new_n1320), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1322), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1351), .B1(new_n1360), .B2(new_n1363), .ZN(G405));
  NAND2_X1  g1164(.A1(new_n1339), .A2(KEYINPUT127), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1363), .A2(new_n1365), .ZN(new_n1366));
  OAI211_X1 g1166(.A(KEYINPUT127), .B(new_n1339), .C1(new_n1361), .C2(new_n1362), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1366), .A2(new_n1367), .ZN(new_n1368));
  OAI21_X1  g1168(.A(new_n1328), .B1(new_n1339), .B2(KEYINPUT127), .ZN(new_n1369));
  AOI21_X1  g1169(.A(new_n1369), .B1(new_n1311), .B2(G375), .ZN(new_n1370));
  XNOR2_X1  g1170(.A(new_n1368), .B(new_n1370), .ZN(G402));
endmodule


