//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981;
  XOR2_X1   g000(.A(KEYINPUT79), .B(KEYINPUT6), .Z(new_n202));
  INV_X1    g001(.A(G141gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT75), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT75), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G141gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n206), .A3(G148gat), .ZN(new_n207));
  INV_X1    g006(.A(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G141gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n207), .A2(new_n209), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G155gat), .B(G162gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n203), .A2(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n209), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n215), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT3), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n210), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(new_n211), .ZN(new_n221));
  XNOR2_X1  g020(.A(G141gat), .B(G148gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(KEYINPUT2), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224));
  INV_X1    g023(.A(new_n209), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT75), .B(G141gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(G148gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n220), .B1(new_n212), .B2(new_n211), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n223), .B(new_n224), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G113gat), .B(G120gat), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n230), .A2(KEYINPUT1), .A3(G134gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n232));
  INV_X1    g031(.A(G120gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G113gat), .ZN(new_n234));
  INV_X1    g033(.A(G113gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G120gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT1), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n232), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(G127gat), .B1(new_n231), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n232), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(new_n230), .B2(KEYINPUT1), .ZN(new_n242));
  INV_X1    g041(.A(G134gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n237), .A2(new_n238), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G127gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n219), .A2(new_n229), .A3(new_n240), .A4(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT5), .ZN(new_n248));
  NAND2_X1  g047(.A1(G225gat), .A2(G233gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n214), .A2(new_n218), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n245), .B1(new_n242), .B2(new_n244), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT4), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n246), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n256), .A2(new_n257), .A3(new_n251), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n250), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n255), .A2(new_n258), .A3(KEYINPUT76), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n257), .B1(new_n256), .B2(new_n251), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT76), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n249), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n260), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n223), .B1(new_n227), .B2(new_n228), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n240), .A2(new_n267), .A3(new_n246), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n254), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n249), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n248), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n259), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT78), .ZN(new_n274));
  XOR2_X1   g073(.A(G1gat), .B(G29gat), .Z(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G57gat), .B(G85gat), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n276), .B(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n202), .B1(new_n272), .B2(new_n280), .ZN(new_n281));
  AOI211_X1 g080(.A(new_n279), .B(new_n259), .C1(new_n266), .C2(new_n271), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT80), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n269), .A2(new_n270), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT5), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n264), .B1(new_n262), .B2(new_n261), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n285), .B1(new_n260), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n279), .B1(new_n287), .B2(new_n259), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n280), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT80), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .A4(new_n202), .ZN(new_n291));
  INV_X1    g090(.A(new_n202), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n279), .B(new_n292), .C1(new_n287), .C2(new_n259), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n283), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT34), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT65), .ZN(new_n296));
  AND2_X1   g095(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT23), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(G169gat), .ZN(new_n301));
  INV_X1    g100(.A(G169gat), .ZN(new_n302));
  INV_X1    g101(.A(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT23), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n299), .A2(new_n301), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n308), .A2(KEYINPUT24), .ZN(new_n309));
  INV_X1    g108(.A(G183gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G190gat), .ZN(new_n311));
  INV_X1    g110(.A(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G183gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n309), .B1(new_n314), .B2(KEYINPUT24), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT25), .B1(new_n307), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n309), .ZN(new_n317));
  XNOR2_X1  g116(.A(G183gat), .B(G190gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT24), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n302), .A2(new_n303), .A3(KEYINPUT23), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n300), .B1(G169gat), .B2(G176gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323));
  OAI211_X1 g122(.A(KEYINPUT25), .B(new_n321), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n296), .B1(new_n316), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT25), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT64), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n303), .ZN(new_n329));
  NAND2_X1  g128(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n301), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n306), .A2(new_n304), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n327), .B1(new_n320), .B2(new_n333), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n315), .A2(KEYINPUT25), .A3(new_n332), .A4(new_n321), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT65), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n326), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n310), .A2(KEYINPUT27), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT27), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G183gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n338), .A2(new_n340), .A3(new_n312), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT28), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT27), .B(G183gat), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(KEYINPUT28), .A3(new_n312), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n302), .A2(new_n303), .A3(KEYINPUT26), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT26), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n348), .B1(G169gat), .B2(G176gat), .ZN(new_n349));
  INV_X1    g148(.A(new_n305), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n347), .B(new_n308), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n346), .A2(KEYINPUT66), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT66), .B1(new_n346), .B2(new_n352), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n256), .B1(new_n337), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n351), .B1(new_n343), .B2(new_n345), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(KEYINPUT66), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n252), .A2(new_n253), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n358), .A2(new_n326), .A3(new_n336), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G227gat), .ZN(new_n362));
  INV_X1    g161(.A(G233gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n295), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  AOI211_X1 g165(.A(KEYINPUT34), .B(new_n364), .C1(new_n356), .C2(new_n360), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n356), .A2(new_n364), .A3(new_n360), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT32), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT33), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(G15gat), .B(G43gat), .Z(new_n373));
  XNOR2_X1  g172(.A(G71gat), .B(G99gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n375), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n369), .B(KEYINPUT32), .C1(new_n371), .C2(new_n377), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n368), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n366), .ZN(new_n380));
  INV_X1    g179(.A(new_n367), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n376), .A2(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G226gat), .A2(G233gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n384), .B(KEYINPUT72), .Z(new_n385));
  OAI21_X1  g184(.A(new_n385), .B1(new_n337), .B2(new_n355), .ZN(new_n386));
  INV_X1    g185(.A(new_n385), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n357), .B1(new_n334), .B2(new_n335), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n387), .B1(new_n388), .B2(KEYINPUT29), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT73), .ZN(new_n390));
  XNOR2_X1  g189(.A(G211gat), .B(G218gat), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT70), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT71), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n391), .A2(new_n392), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n391), .A2(new_n392), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(KEYINPUT71), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT69), .B(G197gat), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n400), .A2(G204gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(G204gat), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n399), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n395), .A2(new_n398), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G204gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n400), .B(new_n405), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n394), .B(new_n393), .C1(new_n406), .C2(new_n399), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT73), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n410), .B(new_n387), .C1(new_n388), .C2(KEYINPUT29), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n386), .A2(new_n390), .A3(new_n409), .A4(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n385), .A2(KEYINPUT29), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(new_n337), .B2(new_n355), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n388), .A2(new_n385), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n408), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G8gat), .B(G36gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(G64gat), .B(G92gat), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n417), .B(new_n418), .Z(new_n419));
  NAND3_X1  g218(.A1(new_n412), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT74), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n422), .B1(new_n420), .B2(new_n421), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n419), .B1(new_n412), .B2(new_n416), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(G228gat), .A2(G233gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(G22gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n429), .B(new_n430), .Z(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G78gat), .B(G106gat), .ZN(new_n433));
  INV_X1    g232(.A(G50gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT29), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n404), .A2(new_n437), .A3(new_n407), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n224), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n267), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n229), .A2(new_n437), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n408), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n436), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n251), .B1(new_n438), .B2(new_n224), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n408), .A2(new_n441), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n444), .A2(new_n445), .A3(new_n435), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n432), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n440), .A2(new_n442), .A3(new_n436), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n435), .B1(new_n444), .B2(new_n445), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n431), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n294), .A2(new_n383), .A3(new_n427), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n376), .A2(new_n378), .ZN(new_n453));
  INV_X1    g252(.A(new_n368), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT68), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n368), .A2(new_n376), .A3(new_n378), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n382), .A2(KEYINPUT68), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n293), .B1(new_n281), .B2(new_n282), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n420), .A2(new_n421), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n426), .B1(new_n462), .B2(KEYINPUT30), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT35), .B1(new_n447), .B2(new_n450), .ZN(new_n464));
  AND4_X1   g263(.A1(new_n423), .A2(new_n461), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n452), .A2(KEYINPUT35), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n451), .B1(new_n294), .B2(new_n427), .ZN(new_n467));
  INV_X1    g266(.A(new_n451), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT38), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n412), .A2(new_n416), .ZN(new_n470));
  INV_X1    g269(.A(new_n419), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(KEYINPUT37), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT37), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n475), .B1(new_n412), .B2(new_n416), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n469), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n420), .B(new_n293), .C1(new_n281), .C2(new_n282), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT82), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n358), .A2(new_n326), .A3(new_n336), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n482), .A2(new_n413), .B1(new_n385), .B2(new_n388), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n475), .B1(new_n483), .B2(new_n409), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n386), .A2(new_n390), .A3(new_n408), .A4(new_n411), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT38), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n474), .A2(new_n481), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n483), .A2(new_n409), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(KEYINPUT37), .A3(new_n485), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n469), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n471), .B1(new_n470), .B2(KEYINPUT37), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT82), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n468), .B1(new_n480), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n463), .A2(new_n423), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n272), .A2(new_n280), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT40), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n254), .A2(new_n268), .A3(new_n249), .ZN(new_n498));
  INV_X1    g297(.A(new_n247), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n499), .B1(new_n255), .B2(new_n258), .ZN(new_n500));
  OAI211_X1 g299(.A(KEYINPUT39), .B(new_n498), .C1(new_n500), .C2(new_n249), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT39), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n255), .A2(new_n258), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n502), .B(new_n270), .C1(new_n503), .C2(new_n499), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n501), .A2(new_n280), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n496), .B1(new_n497), .B2(new_n505), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n505), .A2(new_n497), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n495), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n467), .B1(new_n494), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n383), .A2(KEYINPUT36), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(new_n460), .B2(KEYINPUT36), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n466), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(G29gat), .A2(G36gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT14), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G36gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT84), .B(G29gat), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G43gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n434), .ZN(new_n520));
  NAND2_X1  g319(.A1(G43gat), .A2(G50gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT15), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT85), .B(G50gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(G43gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT86), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT86), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n530), .B(new_n526), .C1(new_n527), .C2(G43gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(KEYINPUT84), .B(G29gat), .Z(new_n533));
  NAND3_X1  g332(.A1(new_n533), .A2(KEYINPUT87), .A3(G36gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT87), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(new_n517), .B2(new_n516), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n534), .A2(new_n536), .A3(new_n515), .A4(new_n523), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n525), .B1(new_n532), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G15gat), .B(G22gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n541), .A2(G1gat), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G8gat), .ZN(new_n544));
  INV_X1    g343(.A(G1gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT16), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n543), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n544), .B1(new_n543), .B2(new_n547), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g349(.A(KEYINPUT17), .B(new_n525), .C1(new_n532), .C2(new_n537), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n540), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n548), .A2(new_n549), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n538), .ZN(new_n554));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n552), .A2(KEYINPUT18), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n550), .B(new_n525), .C1(new_n537), .C2(new_n532), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n554), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n555), .B(KEYINPUT13), .Z(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT18), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT88), .ZN(new_n565));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(G169gat), .B(G197gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT12), .Z(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n561), .B(new_n564), .C1(new_n565), .C2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n560), .A3(new_n565), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n562), .A2(new_n563), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n556), .A2(new_n560), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n574), .B(new_n571), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n512), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G120gat), .B(G148gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(G176gat), .B(G204gat), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n581), .B(new_n582), .Z(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT96), .ZN(new_n586));
  OR2_X1    g385(.A1(G57gat), .A2(G64gat), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT89), .ZN(new_n588));
  NAND2_X1  g387(.A1(G57gat), .A2(G64gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G71gat), .B(G78gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(G71gat), .ZN(new_n593));
  INV_X1    g392(.A(G78gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n595), .A2(KEYINPUT9), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n592), .A2(new_n596), .A3(new_n587), .A4(new_n589), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n587), .B(new_n589), .C1(new_n595), .C2(KEYINPUT9), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(new_n591), .A3(new_n590), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G99gat), .ZN(new_n601));
  INV_X1    g400(.A(G106gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G99gat), .A2(G106gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT92), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT92), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n603), .A2(new_n607), .A3(new_n604), .ZN(new_n608));
  INV_X1    g407(.A(G85gat), .ZN(new_n609));
  INV_X1    g408(.A(G92gat), .ZN(new_n610));
  AOI22_X1  g409(.A1(KEYINPUT8), .A2(new_n604), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G85gat), .A2(G92gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT7), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n606), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  AND4_X1   g414(.A1(new_n606), .A2(new_n614), .A3(new_n608), .A4(new_n611), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n600), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(new_n608), .A3(new_n611), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n618), .A2(KEYINPUT92), .A3(new_n605), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n612), .A2(new_n606), .A3(new_n614), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n619), .A2(new_n620), .A3(new_n597), .A4(new_n599), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(new_n621), .A3(KEYINPUT94), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n620), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT94), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(new_n624), .A3(new_n600), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT10), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT95), .B1(new_n617), .B2(new_n627), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT95), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n623), .A2(new_n630), .A3(KEYINPUT10), .A4(new_n600), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n586), .B1(new_n628), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n622), .A2(new_n586), .A3(new_n625), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n622), .A2(KEYINPUT97), .A3(new_n586), .A4(new_n625), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n584), .B1(new_n634), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n586), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT10), .B1(new_n622), .B2(new_n625), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n641), .B1(new_n642), .B2(new_n632), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n643), .A2(new_n583), .A3(new_n637), .A4(new_n638), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n640), .A2(KEYINPUT98), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT98), .B1(new_n640), .B2(new_n644), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n553), .B1(KEYINPUT21), .B2(new_n600), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n597), .A2(new_n599), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT90), .B(KEYINPUT21), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G231gat), .A2(G233gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(G127gat), .B(G155gat), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT91), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(G183gat), .B(G211gat), .Z(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n657), .A2(new_n660), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n663), .B1(new_n661), .B2(new_n664), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n652), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n667), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n669), .A2(new_n665), .A3(new_n651), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(G232gat), .A2(G233gat), .ZN(new_n672));
  AOI22_X1  g471(.A1(new_n538), .A2(new_n623), .B1(KEYINPUT41), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n540), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n551), .A2(new_n619), .A3(new_n620), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XOR2_X1   g475(.A(G190gat), .B(G218gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n672), .A2(KEYINPUT41), .ZN(new_n679));
  XNOR2_X1  g478(.A(G134gat), .B(G162gat), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n679), .B(new_n680), .Z(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT93), .Z(new_n682));
  NAND2_X1  g481(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n681), .A2(KEYINPUT93), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n683), .B1(new_n684), .B2(new_n678), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n671), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n648), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n294), .B(KEYINPUT99), .Z(new_n688));
  NAND3_X1  g487(.A1(new_n580), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT100), .B(G1gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1324gat));
  NAND3_X1  g490(.A1(new_n580), .A2(new_n495), .A3(new_n687), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n544), .A2(KEYINPUT42), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(new_n693), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n692), .A2(KEYINPUT42), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT16), .B(G8gat), .ZN(new_n699));
  NOR2_X1   g498(.A1(KEYINPUT102), .A2(KEYINPUT42), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n697), .A2(KEYINPUT103), .A3(new_n702), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1325gat));
  NAND2_X1  g506(.A1(new_n580), .A2(new_n687), .ZN(new_n708));
  OAI21_X1  g507(.A(G15gat), .B1(new_n708), .B2(new_n511), .ZN(new_n709));
  INV_X1    g508(.A(G15gat), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n460), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n708), .B2(new_n711), .ZN(G1326gat));
  NOR2_X1   g511(.A1(new_n708), .A2(new_n451), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT43), .B(G22gat), .Z(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1327gat));
  INV_X1    g514(.A(new_n671), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n647), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n685), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n580), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(new_n517), .A3(new_n688), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT45), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n512), .B2(new_n685), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n487), .A2(new_n492), .ZN(new_n725));
  OAI21_X1  g524(.A(KEYINPUT38), .B1(new_n491), .B2(new_n476), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n288), .A2(new_n289), .A3(new_n202), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n726), .A2(new_n420), .A3(new_n727), .A4(new_n293), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n508), .B(new_n451), .C1(new_n725), .C2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n467), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n511), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n452), .A2(KEYINPUT35), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n460), .A2(new_n465), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n685), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT44), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n578), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n573), .A2(new_n577), .A3(KEYINPUT104), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(new_n717), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n724), .A2(new_n736), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n688), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n533), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n722), .A2(new_n745), .ZN(G1328gat));
  NOR3_X1   g545(.A1(new_n719), .A2(G36gat), .A3(new_n427), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT46), .ZN(new_n748));
  OAI21_X1  g547(.A(G36gat), .B1(new_n743), .B2(new_n427), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1329gat));
  OAI21_X1  g549(.A(G43gat), .B1(new_n743), .B2(new_n511), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT47), .B1(new_n751), .B2(KEYINPUT105), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n720), .A2(new_n519), .A3(new_n460), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n752), .B(new_n754), .ZN(G1330gat));
  NOR2_X1   g554(.A1(new_n719), .A2(new_n451), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n468), .A2(new_n527), .ZN(new_n757));
  OAI22_X1  g556(.A1(new_n756), .A2(new_n527), .B1(new_n743), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g558(.A1(new_n512), .A2(new_n686), .A3(new_n647), .A4(new_n740), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n688), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g561(.A(new_n427), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n764), .B(new_n765), .Z(G1333gat));
  XNOR2_X1  g565(.A(new_n460), .B(KEYINPUT106), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(G71gat), .B1(new_n760), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n511), .A2(new_n593), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n760), .B2(new_n770), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g571(.A1(new_n760), .A2(new_n468), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g573(.A1(new_n716), .A2(KEYINPUT107), .A3(new_n741), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n740), .B2(new_n671), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n647), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n724), .A2(new_n736), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT108), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n724), .A2(new_n736), .A3(KEYINPUT108), .A4(new_n778), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(new_n688), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G85gat), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n731), .A2(new_n734), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n775), .A2(new_n777), .ZN(new_n786));
  INV_X1    g585(.A(new_n685), .ZN(new_n787));
  AND4_X1   g586(.A1(KEYINPUT51), .A2(new_n785), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT51), .B1(new_n735), .B2(new_n786), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n791), .A2(new_n609), .A3(new_n648), .A4(new_n688), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n784), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n784), .A2(KEYINPUT109), .A3(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1336gat));
  NOR3_X1   g596(.A1(new_n647), .A2(G92gat), .A3(new_n427), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(new_n791), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(G92gat), .B1(new_n779), .B2(new_n427), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n799), .A2(KEYINPUT111), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT111), .B1(new_n799), .B2(new_n800), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n781), .A2(new_n495), .A3(new_n782), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n798), .B(KEYINPUT110), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n803), .A2(G92gat), .B1(new_n791), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  OAI22_X1  g605(.A1(new_n801), .A2(new_n802), .B1(new_n805), .B2(new_n806), .ZN(G1337gat));
  NAND2_X1  g606(.A1(new_n781), .A2(new_n782), .ZN(new_n808));
  OAI21_X1  g607(.A(G99gat), .B1(new_n808), .B2(new_n511), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n648), .A2(new_n460), .A3(new_n601), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT112), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n790), .B2(new_n811), .ZN(G1338gat));
  NOR3_X1   g611(.A1(new_n647), .A2(G106gat), .A3(new_n451), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(KEYINPUT113), .Z(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n788), .B2(new_n789), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g616(.A(KEYINPUT114), .B(new_n814), .C1(new_n788), .C2(new_n789), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n781), .A2(new_n468), .A3(new_n782), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(G106gat), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n779), .A2(new_n451), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n602), .ZN(new_n824));
  INV_X1    g623(.A(new_n813), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n822), .B1(new_n790), .B2(new_n825), .ZN(new_n826));
  OAI22_X1  g625(.A1(new_n821), .A2(new_n822), .B1(new_n824), .B2(new_n826), .ZN(G1339gat));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n828), .B(new_n641), .C1(new_n642), .C2(new_n632), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n584), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n628), .A2(new_n633), .A3(new_n586), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(KEYINPUT54), .A3(new_n643), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(new_n832), .A3(KEYINPUT55), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(new_n644), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n830), .A2(new_n832), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n834), .A2(new_n738), .A3(new_n739), .A4(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n561), .A2(new_n572), .A3(new_n564), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n558), .A2(new_n559), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n555), .B1(new_n552), .B2(new_n554), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n570), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g643(.A(KEYINPUT115), .B(new_n570), .C1(new_n840), .C2(new_n841), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n839), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n645), .B2(new_n646), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n787), .B1(new_n838), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n837), .A2(new_n644), .A3(new_n833), .ZN(new_n849));
  INV_X1    g648(.A(new_n846), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n849), .A2(new_n850), .A3(new_n685), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n716), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n687), .A2(new_n741), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n468), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n744), .A2(new_n495), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n460), .A3(new_n855), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(KEYINPUT116), .Z(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(G113gat), .B1(new_n858), .B2(new_n579), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n744), .B1(new_n852), .B2(new_n853), .ZN(new_n860));
  AND4_X1   g659(.A1(new_n427), .A2(new_n860), .A3(new_n383), .A4(new_n451), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n740), .A2(new_n235), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT117), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n859), .A2(new_n864), .ZN(G1340gat));
  AOI21_X1  g664(.A(G120gat), .B1(new_n861), .B2(new_n648), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n647), .A2(new_n233), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n857), .B2(new_n867), .ZN(G1341gat));
  XNOR2_X1  g667(.A(KEYINPUT67), .B(G127gat), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(new_n861), .B2(new_n671), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n671), .A2(new_n869), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n857), .B2(new_n871), .ZN(G1342gat));
  OAI21_X1  g671(.A(G134gat), .B1(new_n858), .B2(new_n685), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n861), .A2(new_n243), .A3(new_n787), .ZN(new_n874));
  XOR2_X1   g673(.A(new_n874), .B(KEYINPUT56), .Z(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(G1343gat));
  AND2_X1   g675(.A1(new_n855), .A2(new_n511), .ZN(new_n877));
  XNOR2_X1  g676(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n852), .A2(new_n853), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(new_n468), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n837), .A2(new_n578), .A3(new_n644), .A4(new_n833), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n787), .B1(new_n847), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n716), .B1(new_n883), .B2(new_n851), .ZN(new_n884));
  AOI211_X1 g683(.A(new_n881), .B(new_n451), .C1(new_n884), .C2(new_n853), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n740), .B(new_n877), .C1(new_n880), .C2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887));
  INV_X1    g686(.A(new_n226), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n887), .B1(new_n886), .B2(new_n888), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n511), .A2(new_n427), .A3(new_n468), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n578), .A2(new_n203), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT120), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n860), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n889), .A2(new_n890), .A3(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT58), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n880), .A2(new_n885), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n899), .A2(new_n877), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n226), .B1(new_n900), .B2(new_n578), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT58), .B1(new_n895), .B2(KEYINPUT121), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(KEYINPUT121), .B2(new_n895), .ZN(new_n903));
  OAI22_X1  g702(.A1(new_n897), .A2(new_n898), .B1(new_n901), .B2(new_n903), .ZN(G1344gat));
  NAND2_X1  g703(.A1(new_n687), .A2(new_n579), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n884), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g705(.A(KEYINPUT122), .B(new_n881), .C1(new_n906), .C2(new_n451), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n879), .A2(new_n468), .A3(new_n878), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n451), .B1(new_n884), .B2(new_n905), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(KEYINPUT57), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n907), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n648), .A3(new_n877), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n914));
  INV_X1    g713(.A(new_n877), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n915), .A2(KEYINPUT59), .A3(new_n647), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n860), .A2(new_n891), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT59), .B1(new_n917), .B2(new_n647), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n916), .A2(new_n899), .B1(new_n208), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n914), .A2(new_n919), .ZN(G1345gat));
  INV_X1    g719(.A(G155gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n921), .B1(new_n900), .B2(new_n671), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n917), .A2(G155gat), .A3(new_n716), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n922), .A2(new_n923), .ZN(G1346gat));
  INV_X1    g723(.A(G162gat), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n685), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n860), .A2(new_n787), .A3(new_n891), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n900), .A2(new_n926), .B1(new_n927), .B2(new_n925), .ZN(G1347gat));
  AOI21_X1  g727(.A(new_n688), .B1(new_n852), .B2(new_n853), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n929), .A2(KEYINPUT123), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(KEYINPUT123), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n383), .A2(new_n495), .A3(new_n451), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT124), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n932), .A2(new_n936), .A3(new_n933), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n935), .A2(new_n302), .A3(new_n740), .A4(new_n937), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n767), .A2(new_n688), .A3(new_n427), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n854), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(G169gat), .B1(new_n940), .B2(new_n579), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT125), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n938), .A2(new_n942), .ZN(G1348gat));
  NOR3_X1   g742(.A1(new_n940), .A2(new_n299), .A3(new_n647), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n935), .A2(new_n648), .A3(new_n937), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(new_n303), .ZN(G1349gat));
  OAI21_X1  g745(.A(G183gat), .B1(new_n940), .B2(new_n716), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n671), .A2(new_n344), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n934), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g749(.A1(new_n935), .A2(new_n312), .A3(new_n787), .A4(new_n937), .ZN(new_n951));
  OAI21_X1  g750(.A(G190gat), .B1(new_n940), .B2(new_n685), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1351gat));
  NAND3_X1  g753(.A1(new_n511), .A2(new_n495), .A3(new_n468), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n955), .B1(new_n930), .B2(new_n931), .ZN(new_n956));
  AOI21_X1  g755(.A(G197gat), .B1(new_n956), .B2(new_n740), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n744), .A2(new_n511), .A3(new_n495), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n912), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n578), .A2(G197gat), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(G1352gat));
  NAND3_X1  g761(.A1(new_n956), .A2(new_n405), .A3(new_n648), .ZN(new_n963));
  OR2_X1    g762(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n964));
  OAI21_X1  g763(.A(G204gat), .B1(new_n959), .B2(new_n647), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(G1353gat));
  NAND3_X1  g766(.A1(new_n912), .A2(new_n671), .A3(new_n958), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(G211gat), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n968), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n971), .A2(KEYINPUT126), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT63), .B1(new_n968), .B2(G211gat), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n716), .A2(G211gat), .ZN(new_n976));
  AOI22_X1  g775(.A1(new_n974), .A2(new_n975), .B1(new_n956), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n973), .A2(new_n977), .ZN(G1354gat));
  OAI21_X1  g777(.A(G218gat), .B1(new_n959), .B2(new_n685), .ZN(new_n979));
  INV_X1    g778(.A(G218gat), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n956), .A2(new_n980), .A3(new_n787), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n979), .A2(new_n981), .ZN(G1355gat));
endmodule


