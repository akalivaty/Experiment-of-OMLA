//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n565, new_n566, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT65), .Z(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n464), .B1(new_n465), .B2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G101), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT69), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n466), .A2(new_n468), .A3(new_n472), .A4(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT67), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(new_n477), .A3(G2104), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n475), .A2(new_n478), .B1(KEYINPUT3), .B2(new_n465), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(G137), .A3(new_n467), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n477), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G125), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n474), .A2(new_n480), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G160));
  NAND2_X1  g064(.A1(new_n479), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n479), .A2(new_n467), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G136), .ZN(new_n495));
  OR2_X1    g070(.A1(G100), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n497), .B(KEYINPUT70), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n492), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G162));
  NAND2_X1  g075(.A1(new_n475), .A2(new_n478), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(G126), .A3(new_n482), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT71), .A2(G114), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT71), .A2(G114), .ZN(new_n504));
  NOR3_X1   g079(.A1(new_n503), .A2(new_n504), .A3(new_n465), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n467), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G138), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n508), .A2(G2105), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n501), .A2(KEYINPUT4), .A3(new_n482), .A4(new_n509), .ZN(new_n510));
  AND3_X1   g085(.A1(new_n467), .A2(G102), .A3(G2104), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n509), .A2(new_n482), .A3(new_n483), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n507), .A2(new_n515), .ZN(G164));
  XOR2_X1   g091(.A(KEYINPUT73), .B(G88), .Z(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT72), .B1(new_n518), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n518), .A2(G543), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n517), .A2(new_n523), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G50), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(G543), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n523), .A2(G62), .A3(new_n524), .ZN(new_n531));
  NAND2_X1  g106(.A1(G75), .A2(G543), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT74), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n536), .B1(new_n529), .B2(new_n533), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(G166));
  AND2_X1   g113(.A1(new_n523), .A2(new_n524), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n539), .A2(G63), .A3(G651), .ZN(new_n540));
  INV_X1    g115(.A(new_n528), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G51), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT75), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT7), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n539), .A2(G89), .A3(new_n525), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n545), .A2(KEYINPUT76), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(KEYINPUT76), .B1(new_n545), .B2(new_n546), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n540), .B(new_n542), .C1(new_n547), .C2(new_n548), .ZN(G286));
  INV_X1    g124(.A(G286), .ZN(G168));
  AOI22_X1  g125(.A1(new_n539), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n530), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n541), .A2(G52), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n539), .A2(new_n525), .ZN(new_n554));
  INV_X1    g129(.A(G90), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n552), .A2(new_n556), .ZN(G171));
  AOI22_X1  g132(.A1(new_n539), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(new_n530), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n541), .A2(G43), .ZN(new_n560));
  INV_X1    g135(.A(G81), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n554), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  AND3_X1   g139(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G36), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT77), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n565), .A2(new_n569), .ZN(G188));
  NAND3_X1  g145(.A1(new_n539), .A2(G91), .A3(new_n525), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT9), .B1(new_n528), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n525), .A2(new_n574), .A3(G53), .A4(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g151(.A1(G78), .A2(G543), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n539), .B2(G65), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n571), .B(new_n576), .C1(new_n578), .C2(new_n530), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  INV_X1    g155(.A(G166), .ZN(G303));
  INV_X1    g156(.A(new_n554), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G87), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n539), .B2(G74), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n541), .A2(G49), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  NAND3_X1  g161(.A1(new_n523), .A2(G61), .A3(new_n524), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n530), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n523), .A2(G86), .A3(new_n524), .A4(new_n525), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n525), .A2(G48), .A3(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G305));
  NAND2_X1  g169(.A1(G72), .A2(G543), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n523), .A2(new_n524), .ZN(new_n596));
  INV_X1    g171(.A(G60), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n541), .A2(G47), .ZN(new_n600));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n554), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(KEYINPUT78), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n602), .A2(KEYINPUT78), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n599), .B1(new_n604), .B2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n596), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G651), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n523), .A2(G92), .A3(new_n524), .A4(new_n525), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n541), .A2(G54), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n611), .A2(new_n612), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n610), .A2(new_n613), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G171), .B2(new_n617), .ZN(G284));
  OAI21_X1  g194(.A(new_n618), .B1(G171), .B2(new_n617), .ZN(G321));
  NAND2_X1  g195(.A1(G299), .A2(new_n617), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G168), .B2(new_n617), .ZN(G297));
  OAI21_X1  g197(.A(new_n621), .B1(G168), .B2(new_n617), .ZN(G280));
  INV_X1    g198(.A(new_n616), .ZN(new_n624));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G860), .ZN(G148));
  OAI21_X1  g201(.A(KEYINPUT80), .B1(new_n563), .B2(G868), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n616), .A2(G559), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n628), .A2(new_n617), .ZN(new_n629));
  MUX2_X1   g204(.A(new_n627), .B(KEYINPUT80), .S(new_n629), .Z(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT81), .Z(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g207(.A1(new_n469), .A2(new_n484), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT82), .B(G2100), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n491), .A2(G123), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n494), .A2(G135), .ZN(new_n639));
  NOR2_X1   g214(.A1(G99), .A2(G2105), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(new_n467), .B2(G111), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n638), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(G2096), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n637), .A2(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT85), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2427), .B(G2430), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(KEYINPUT14), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2446), .ZN(new_n653));
  XOR2_X1   g228(.A(KEYINPUT84), .B(G2443), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n651), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n658), .A2(new_n661), .A3(new_n659), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(G14), .A3(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT86), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G401));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2072), .B(G2078), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT18), .Z(new_n675));
  XOR2_X1   g250(.A(new_n672), .B(KEYINPUT87), .Z(new_n676));
  OAI21_X1  g251(.A(KEYINPUT17), .B1(new_n676), .B2(new_n671), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(new_n673), .Z(new_n678));
  AND2_X1   g253(.A1(new_n676), .A2(new_n671), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n675), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(new_n643), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(G2100), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G227));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT88), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT20), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n689), .A2(new_n690), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n693), .B1(new_n688), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n688), .A2(new_n694), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT89), .Z(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(G1986), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  OR3_X1    g275(.A1(new_n696), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n696), .B2(new_n698), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n685), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT22), .B(G1981), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n701), .A2(new_n685), .A3(new_n702), .ZN(new_n706));
  AND3_X1   g281(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n705), .B1(new_n704), .B2(new_n706), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(G229));
  NAND2_X1  g285(.A1(new_n624), .A2(G16), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G4), .B2(G16), .ZN(new_n712));
  INV_X1    g287(.A(G1348), .ZN(new_n713));
  NOR2_X1   g288(.A1(G27), .A2(G29), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G164), .B2(G29), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n712), .A2(new_n713), .B1(G2078), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(KEYINPUT98), .B1(G29), .B2(G33), .ZN(new_n717));
  OR3_X1    g292(.A1(KEYINPUT98), .A2(G29), .A3(G33), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT25), .Z(new_n720));
  INV_X1    g295(.A(G139), .ZN(new_n721));
  INV_X1    g296(.A(new_n484), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n722), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n723));
  OAI221_X1 g298(.A(new_n720), .B1(new_n493), .B2(new_n721), .C1(new_n723), .C2(new_n467), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n717), .B(new_n718), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G2072), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n716), .B(new_n727), .C1(new_n713), .C2(new_n712), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT31), .B(G11), .Z(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n730), .A2(KEYINPUT23), .A3(G20), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT23), .ZN(new_n732));
  INV_X1    g307(.A(G20), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(G16), .ZN(new_n734));
  INV_X1    g309(.A(G299), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n731), .B(new_n734), .C1(new_n735), .C2(new_n730), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1956), .ZN(new_n737));
  NOR3_X1   g312(.A1(new_n728), .A2(new_n729), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n730), .A2(G21), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G168), .B2(new_n730), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT102), .Z(new_n741));
  XOR2_X1   g316(.A(KEYINPUT103), .B(G1966), .Z(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT24), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(G34), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(G34), .ZN(new_n747));
  AOI21_X1  g322(.A(G29), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n488), .B2(G29), .ZN(new_n749));
  INV_X1    g324(.A(G2084), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n725), .A2(G35), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G162), .B2(new_n725), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT29), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n751), .B1(new_n754), .B2(G2090), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G2090), .B2(new_n754), .ZN(new_n756));
  NOR2_X1   g331(.A1(G16), .A2(G19), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n563), .B2(G16), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n758), .A2(G1341), .ZN(new_n759));
  NOR2_X1   g334(.A1(G5), .A2(G16), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G171), .B2(G16), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(G1961), .ZN(new_n762));
  NOR4_X1   g337(.A1(new_n743), .A2(new_n756), .A3(new_n759), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n715), .A2(G2078), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n741), .B2(new_n742), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT97), .B(KEYINPUT28), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n725), .A2(G26), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  AOI22_X1  g343(.A1(G128), .A2(new_n491), .B1(new_n494), .B2(G140), .ZN(new_n769));
  OR2_X1    g344(.A1(G104), .A2(G2105), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n770), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT96), .Z(new_n772));
  NAND2_X1  g347(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n768), .B1(new_n773), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2067), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n761), .A2(G1961), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT30), .B(G28), .Z(new_n777));
  MUX2_X1   g352(.A(new_n777), .B(new_n642), .S(G29), .Z(new_n778));
  NAND3_X1  g353(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  AND4_X1   g355(.A1(new_n738), .A2(new_n763), .A3(new_n765), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n749), .A2(new_n750), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n730), .A2(G23), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT93), .ZN(new_n784));
  NAND2_X1  g359(.A1(G288), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n583), .A2(KEYINPUT93), .A3(new_n584), .A4(new_n585), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n783), .B1(new_n787), .B2(new_n730), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT33), .B(G1976), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n788), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G16), .A2(G22), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G166), .B2(G16), .ZN(new_n794));
  INV_X1    g369(.A(G1971), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(G6), .A2(G16), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n593), .B2(G16), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT32), .B(G1981), .Z(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT91), .B(KEYINPUT92), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n798), .B(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n792), .A2(new_n796), .A3(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT34), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n730), .A2(G24), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n602), .A2(KEYINPUT78), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n808), .A2(new_n603), .B1(G651), .B2(new_n598), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n807), .B1(new_n809), .B2(new_n730), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(G1986), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(G1986), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n725), .A2(G25), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n491), .A2(G119), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n494), .A2(G131), .ZN(new_n816));
  OR2_X1    g391(.A1(G95), .A2(G2105), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n817), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n814), .B1(new_n820), .B2(new_n725), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT35), .B(G1991), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT90), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n821), .B(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n812), .A2(new_n813), .A3(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  AND3_X1   g401(.A1(new_n805), .A2(new_n806), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n806), .B1(new_n805), .B2(new_n826), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n781), .B(new_n782), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n758), .A2(G1341), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n494), .A2(G141), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT99), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n466), .A2(G105), .A3(new_n468), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT100), .B(KEYINPUT26), .ZN(new_n834));
  NAND3_X1  g409(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  AOI211_X1 g411(.A(new_n833), .B(new_n836), .C1(G129), .C2(new_n491), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G29), .ZN(new_n840));
  NOR2_X1   g415(.A1(G29), .A2(G32), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(KEYINPUT101), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(KEYINPUT101), .B2(new_n840), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT27), .B(G1996), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n829), .A2(new_n830), .A3(new_n845), .ZN(G311));
  OR3_X1    g421(.A1(new_n829), .A2(new_n830), .A3(new_n845), .ZN(G150));
  AOI22_X1  g422(.A1(new_n539), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n848), .A2(new_n530), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(KEYINPUT105), .B(G55), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n541), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(G93), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n554), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G860), .ZN(new_n857));
  XOR2_X1   g432(.A(KEYINPUT107), .B(KEYINPUT37), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n616), .A2(new_n625), .ZN(new_n860));
  XOR2_X1   g435(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n563), .B1(new_n849), .B2(new_n854), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n850), .B(new_n855), .C1(new_n559), .C2(new_n562), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n862), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT106), .ZN(new_n869));
  INV_X1    g444(.A(G860), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(new_n867), .B2(KEYINPUT39), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n859), .B1(new_n869), .B2(new_n871), .ZN(G145));
  XNOR2_X1  g447(.A(new_n642), .B(new_n499), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(G160), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n505), .B1(new_n479), .B2(G126), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n514), .B(new_n510), .C1(new_n875), .C2(new_n467), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n724), .B(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n874), .A2(new_n877), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(G142), .ZN(new_n881));
  NOR2_X1   g456(.A1(G106), .A2(G2105), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(new_n467), .B2(G118), .ZN(new_n883));
  OAI22_X1  g458(.A1(new_n493), .A2(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(G130), .B2(new_n491), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n820), .B(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n839), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n880), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n878), .A2(new_n887), .A3(new_n879), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n773), .B(new_n634), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n889), .A2(new_n892), .A3(new_n890), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g473(.A(KEYINPUT108), .B1(new_n624), .B2(G299), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT108), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n735), .A2(new_n616), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n624), .A2(G299), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n903), .A2(KEYINPUT110), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT110), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n624), .A2(KEYINPUT108), .A3(G299), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n900), .B1(new_n735), .B2(new_n616), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT109), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT109), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n899), .A2(new_n910), .A3(new_n901), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n911), .A3(new_n902), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n906), .B1(new_n912), .B2(new_n904), .ZN(new_n913));
  INV_X1    g488(.A(new_n903), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT41), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n905), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n865), .B(new_n628), .Z(new_n917));
  MUX2_X1   g492(.A(new_n903), .B(new_n916), .S(new_n917), .Z(new_n918));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n787), .B(KEYINPUT111), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n809), .A2(G166), .ZN(new_n923));
  NAND2_X1  g498(.A1(G290), .A2(G303), .ZN(new_n924));
  AOI21_X1  g499(.A(G305), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n924), .A3(G305), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n922), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n927), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n921), .B1(new_n929), .B2(new_n925), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n918), .A2(new_n919), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n920), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n920), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g510(.A(G868), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n856), .A2(new_n617), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(G295));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n937), .ZN(G331));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n912), .A2(new_n904), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(KEYINPUT110), .A3(new_n915), .ZN(new_n943));
  INV_X1    g518(.A(new_n905), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n863), .A2(new_n864), .A3(G301), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(G301), .B1(new_n863), .B2(new_n864), .ZN(new_n947));
  OAI21_X1  g522(.A(G286), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n865), .A2(G171), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n949), .A2(G168), .A3(new_n945), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n943), .A2(new_n944), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n948), .A2(new_n950), .A3(new_n903), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n931), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n895), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n931), .B1(new_n952), .B2(new_n953), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n941), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n953), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n916), .B2(new_n951), .ZN(new_n959));
  AOI21_X1  g534(.A(G37), .B1(new_n959), .B2(new_n931), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n953), .A2(KEYINPUT112), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n948), .A2(new_n950), .A3(new_n962), .A4(new_n903), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n912), .A2(KEYINPUT41), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n914), .A2(new_n904), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n951), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n932), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n960), .A2(KEYINPUT43), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n940), .B1(new_n957), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT43), .B1(new_n955), .B2(new_n956), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n960), .A2(new_n941), .A3(new_n968), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT44), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT113), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n956), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT43), .B1(new_n960), .B2(new_n975), .ZN(new_n976));
  AND4_X1   g551(.A1(KEYINPUT43), .A2(new_n968), .A3(new_n895), .A4(new_n954), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT44), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n941), .B1(new_n960), .B2(new_n975), .ZN(new_n979));
  AND4_X1   g554(.A1(new_n941), .A2(new_n968), .A3(new_n895), .A4(new_n954), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n940), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n978), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n974), .A2(new_n983), .ZN(G397));
  OR2_X1    g559(.A1(new_n773), .A2(G2067), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n773), .A2(G2067), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1996), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n839), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n838), .A2(G1996), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n822), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n819), .B(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT114), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  OR2_X1    g570(.A1(G290), .A2(G1986), .ZN(new_n996));
  NAND2_X1  g571(.A1(G290), .A2(G1986), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(new_n507), .B2(new_n515), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n474), .A2(new_n487), .A3(G40), .A4(new_n480), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n998), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G286), .A2(G8), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT122), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT122), .ZN(new_n1009));
  NAND3_X1  g584(.A1(G286), .A2(new_n1009), .A3(G8), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1003), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n876), .A2(KEYINPUT117), .A3(KEYINPUT45), .A4(new_n999), .ZN(new_n1013));
  OAI211_X1 g588(.A(KEYINPUT45), .B(new_n999), .C1(new_n507), .C2(new_n515), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1012), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n742), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1017), .A2(KEYINPUT118), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT118), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1000), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n876), .A2(KEYINPUT50), .A3(new_n999), .ZN(new_n1023));
  AOI211_X1 g598(.A(G2084), .B(new_n1003), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1019), .A2(new_n1020), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G8), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1006), .B(new_n1011), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT123), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT51), .B1(new_n1025), .B2(new_n1011), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1024), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1017), .A2(KEYINPUT118), .A3(new_n1018), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1030), .B1(new_n1036), .B2(G8), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1027), .B(new_n1028), .C1(new_n1029), .C2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1011), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1006), .B1(new_n1036), .B2(new_n1030), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1028), .B1(new_n1042), .B2(new_n1027), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1003), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1961), .ZN(new_n1048));
  INV_X1    g623(.A(G2078), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1012), .A2(new_n1049), .A3(new_n1014), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1047), .A2(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1051), .A2(G2078), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1052), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1057), .A2(G171), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1012), .A2(new_n1016), .A3(new_n1013), .A4(new_n1055), .ZN(new_n1059));
  AOI21_X1  g634(.A(G301), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1045), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1976), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n785), .B2(new_n786), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1064), .A2(new_n1026), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT52), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G1981), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n593), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT49), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n589), .A2(new_n592), .A3(G1981), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT49), .B1(new_n1073), .B2(KEYINPUT115), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n593), .A2(new_n1068), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1072), .B(new_n1074), .C1(new_n1068), .C2(new_n593), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1065), .A3(new_n1078), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1067), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G2090), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1081), .A2(new_n1046), .B1(new_n1053), .B2(new_n795), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n535), .A2(G8), .A3(new_n537), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n1086), .A3(G8), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n1084), .B(KEYINPUT55), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n1082), .B2(new_n1026), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT52), .B1(G288), .B2(new_n1062), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1080), .A2(new_n1087), .A3(new_n1089), .A4(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(G301), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1097), .A2(new_n1098), .A3(G301), .A4(new_n1059), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1095), .A2(new_n1096), .A3(KEYINPUT54), .A4(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(KEYINPUT54), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT124), .B1(new_n1101), .B2(new_n1094), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1093), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1044), .A2(KEYINPUT125), .A3(new_n1061), .A4(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n1105));
  OR3_X1    g680(.A1(new_n1046), .A2(new_n1105), .A3(G1956), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1105), .B1(new_n1046), .B2(G1956), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT56), .B(G2072), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1106), .A2(new_n1107), .B1(new_n1054), .B2(new_n1108), .ZN(new_n1109));
  XOR2_X1   g684(.A(G299), .B(KEYINPUT57), .Z(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1111), .A2(KEYINPUT61), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT58), .B(G1341), .Z(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1116), .B(new_n1117), .C1(G1996), .C2(new_n1053), .ZN(new_n1118));
  NAND2_X1  g693(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(new_n563), .A3(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1064), .ZN(new_n1123));
  OAI22_X1  g698(.A1(new_n1046), .A2(G1348), .B1(new_n1123), .B2(G2067), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n624), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n616), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1126), .A2(KEYINPUT60), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1121), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1118), .A2(new_n563), .A3(new_n1129), .A4(new_n1119), .ZN(new_n1130));
  OR3_X1    g705(.A1(new_n1124), .A2(KEYINPUT60), .A3(new_n616), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1122), .A2(new_n1128), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1112), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1125), .A2(new_n616), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1111), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1136), .B1(new_n1133), .B2(KEYINPUT61), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1027), .B1(new_n1029), .B2(new_n1037), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT123), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1140), .A2(new_n1103), .A3(new_n1038), .A4(new_n1061), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1104), .A2(new_n1138), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1093), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1140), .A2(KEYINPUT62), .A3(new_n1038), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .A4(new_n1060), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT63), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1147), .A2(new_n1150), .A3(G168), .A4(new_n1151), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1088), .A2(new_n1082), .A3(new_n1026), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1080), .A2(new_n1153), .A3(new_n1092), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1079), .A2(new_n1062), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1069), .B1(new_n1155), .B2(G288), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT116), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1152), .B(new_n1154), .C1(new_n1157), .C2(new_n1066), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1093), .A2(new_n1026), .A3(new_n1025), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1150), .B1(new_n1159), .B2(G168), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1149), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1005), .B1(new_n1144), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1004), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n996), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT126), .ZN(new_n1166));
  XOR2_X1   g741(.A(new_n1166), .B(KEYINPUT48), .Z(new_n1167));
  OAI21_X1  g742(.A(new_n1167), .B1(new_n1164), .B2(new_n995), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1164), .B1(new_n987), .B2(new_n839), .ZN(new_n1169));
  AOI21_X1  g744(.A(KEYINPUT46), .B1(new_n1004), .B2(new_n988), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n1004), .A2(KEYINPUT46), .A3(new_n988), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  XOR2_X1   g747(.A(new_n1172), .B(KEYINPUT47), .Z(new_n1173));
  NAND2_X1  g748(.A1(new_n820), .A2(new_n992), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n985), .B1(new_n991), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1004), .ZN(new_n1176));
  AND3_X1   g751(.A1(new_n1168), .A2(new_n1173), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1163), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g753(.A(new_n462), .B1(new_n667), .B2(new_n668), .ZN(new_n1180));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n1181));
  NAND4_X1  g755(.A1(new_n709), .A2(new_n1180), .A3(new_n1181), .A4(new_n682), .ZN(new_n1182));
  NAND2_X1  g756(.A1(new_n1182), .A2(new_n897), .ZN(new_n1183));
  NOR3_X1   g757(.A1(new_n707), .A2(new_n708), .A3(G227), .ZN(new_n1184));
  AOI21_X1  g758(.A(new_n1181), .B1(new_n1184), .B2(new_n1180), .ZN(new_n1185));
  NOR2_X1   g759(.A1(new_n979), .A2(new_n980), .ZN(new_n1186));
  NOR3_X1   g760(.A1(new_n1183), .A2(new_n1185), .A3(new_n1186), .ZN(G308));
  OR3_X1    g761(.A1(new_n1183), .A2(new_n1185), .A3(new_n1186), .ZN(G225));
endmodule


