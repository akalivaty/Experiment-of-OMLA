//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  AND2_X1   g0022(.A1(new_n222), .A2(new_n209), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT64), .Z(new_n226));
  OAI211_X1 g0026(.A(new_n217), .B(new_n226), .C1(new_n224), .C2(new_n223), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT65), .Z(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G68), .Z(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G169), .ZN(new_n246));
  AND2_X1   g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n247), .A2(new_n213), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  AOI21_X1  g0053(.A(G1698), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n254), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(new_n253), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G232), .A3(G1698), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n249), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT13), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT68), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(new_n247), .B2(new_n213), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n265), .A2(KEYINPUT68), .A3(G1), .A4(G13), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n262), .A2(new_n264), .A3(G274), .A4(new_n266), .ZN(new_n267));
  AND3_X1   g0067(.A1(new_n262), .A2(new_n263), .A3(new_n266), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G238), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n259), .A2(new_n260), .A3(new_n267), .A4(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n267), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT13), .B1(new_n271), .B2(new_n258), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n246), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT14), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n270), .A2(new_n272), .ZN(new_n275));
  INV_X1    g0075(.A(G179), .ZN(new_n276));
  OAI22_X1  g0076(.A1(new_n273), .A2(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n273), .A2(new_n274), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT80), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT80), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n273), .A2(new_n280), .A3(new_n274), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n277), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G13), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n283), .A2(new_n207), .A3(G1), .ZN(new_n284));
  INV_X1    g0084(.A(G68), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n286), .B(KEYINPUT12), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n213), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n284), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n206), .A2(G20), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(G68), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT70), .B1(new_n251), .B2(G20), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT70), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n294), .A2(new_n207), .A3(G33), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G77), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n207), .A2(new_n251), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n299), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n289), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT11), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n287), .B(new_n292), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n301), .A2(new_n302), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n282), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n275), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G190), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n275), .A2(G200), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(new_n305), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G200), .ZN(new_n313));
  INV_X1    g0113(.A(G1698), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n252), .B2(new_n253), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n315), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n316));
  AND2_X1   g0116(.A1(KEYINPUT3), .A2(G33), .ZN(new_n317));
  NOR2_X1   g0117(.A1(KEYINPUT3), .A2(G33), .ZN(new_n318));
  OAI211_X1 g0118(.A(G223), .B(new_n314), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n249), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n262), .A2(G232), .A3(new_n263), .A4(new_n266), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n267), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n313), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  OAI211_X1 g0123(.A(G226), .B(G1698), .C1(new_n317), .C2(new_n318), .ZN(new_n324));
  INV_X1    g0124(.A(G87), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n319), .B(new_n324), .C1(new_n251), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n248), .ZN(new_n327));
  INV_X1    g0127(.A(G190), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n327), .A2(new_n328), .A3(new_n267), .A4(new_n321), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT8), .B(G58), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n206), .B2(G20), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n332), .A2(new_n290), .B1(new_n331), .B2(new_n284), .ZN(new_n333));
  NAND3_X1  g0133(.A1(KEYINPUT81), .A2(G58), .A3(G68), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT81), .B1(G58), .B2(G68), .ZN(new_n336));
  NOR3_X1   g0136(.A1(new_n335), .A2(new_n336), .A3(new_n201), .ZN(new_n337));
  INV_X1    g0137(.A(G159), .ZN(new_n338));
  OAI22_X1  g0138(.A1(new_n337), .A2(new_n207), .B1(new_n338), .B2(new_n299), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n317), .A2(new_n318), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT7), .B1(new_n340), .B2(new_n207), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n253), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(G68), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT82), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n339), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n252), .A2(new_n207), .A3(new_n253), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT7), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n285), .B1(new_n349), .B2(new_n342), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT82), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT16), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n336), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n353), .B(new_n334), .C1(G58), .C2(G68), .ZN(new_n354));
  INV_X1    g0154(.A(new_n299), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n354), .A2(G20), .B1(G159), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n344), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT16), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n289), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n330), .B(new_n333), .C1(new_n352), .C2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT17), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n333), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n356), .B1(new_n350), .B2(KEYINPUT82), .ZN(new_n364));
  AOI211_X1 g0164(.A(new_n345), .B(new_n285), .C1(new_n349), .C2(new_n342), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n358), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n289), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n350), .A2(new_n339), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n367), .B1(new_n368), .B2(KEYINPUT16), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n363), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(KEYINPUT17), .A3(new_n330), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT84), .B1(new_n362), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n362), .A2(KEYINPUT84), .A3(new_n371), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n333), .B1(new_n352), .B2(new_n359), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT83), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT83), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n370), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n327), .A2(new_n267), .A3(new_n321), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G169), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n380), .B2(new_n276), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n377), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT18), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT18), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n377), .A2(new_n379), .A3(new_n385), .A4(new_n382), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n312), .A2(new_n375), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G150), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n299), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n331), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n293), .A2(new_n295), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n393), .A2(KEYINPUT71), .B1(G20), .B2(new_n203), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT71), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n296), .A2(new_n331), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n395), .B1(new_n396), .B2(new_n390), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n367), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n290), .A2(G50), .A3(new_n291), .ZN(new_n399));
  INV_X1    g0199(.A(new_n284), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n399), .B1(G50), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT9), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT9), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n398), .B2(new_n401), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n268), .A2(G226), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n267), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n254), .A2(G222), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n315), .A2(G223), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n340), .A2(G77), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n249), .B1(new_n411), .B2(KEYINPUT69), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT69), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n408), .A2(new_n409), .A3(new_n413), .A4(new_n410), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n407), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G190), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n403), .A2(new_n405), .A3(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(KEYINPUT10), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n412), .A2(new_n414), .ZN(new_n419));
  INV_X1    g0219(.A(new_n407), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT76), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(G200), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT76), .B1(new_n415), .B2(new_n313), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT77), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT77), .B1(new_n423), .B2(new_n424), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n418), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT78), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(KEYINPUT10), .C1(new_n417), .C2(new_n425), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n402), .A2(KEYINPUT9), .B1(G190), .B2(new_n415), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n433), .A2(new_n423), .A3(new_n424), .A4(new_n405), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n430), .B1(new_n434), .B2(KEYINPUT10), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n429), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n402), .B1(new_n246), .B2(new_n421), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(G179), .B2(new_n421), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n268), .A2(G244), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n267), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT72), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT72), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n439), .A2(new_n442), .A3(new_n267), .ZN(new_n443));
  XNOR2_X1  g0243(.A(KEYINPUT73), .B(G107), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n315), .A2(G238), .B1(new_n340), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n256), .A2(G232), .A3(new_n314), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n248), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n441), .A2(new_n443), .A3(new_n448), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n449), .A2(new_n328), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(G200), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n297), .B1(new_n206), .B2(G20), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n290), .A2(new_n452), .B1(new_n297), .B2(new_n284), .ZN(new_n453));
  XNOR2_X1  g0253(.A(KEYINPUT15), .B(G87), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n296), .A2(new_n454), .ZN(new_n455));
  OAI22_X1  g0255(.A1(new_n331), .A2(new_n299), .B1(new_n207), .B2(new_n297), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n289), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n457), .A2(KEYINPUT74), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(KEYINPUT74), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n453), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT75), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(KEYINPUT75), .B(new_n453), .C1(new_n458), .C2(new_n459), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n450), .A2(new_n451), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n449), .A2(new_n246), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n465), .B(new_n460), .C1(G179), .C2(new_n449), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n436), .A2(new_n438), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT79), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT79), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n436), .A2(new_n470), .A3(new_n438), .A4(new_n467), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n388), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n262), .A2(G274), .A3(new_n266), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT5), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G41), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n476), .A2(KEYINPUT86), .A3(new_n206), .A4(G45), .ZN(new_n477));
  INV_X1    g0277(.A(G41), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n206), .B(G45), .C1(new_n478), .C2(KEYINPUT5), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT86), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n479), .A2(new_n480), .B1(KEYINPUT5), .B2(new_n478), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n474), .A2(KEYINPUT87), .A3(new_n477), .A4(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT87), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n479), .A2(new_n480), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n478), .A2(KEYINPUT5), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n484), .A2(new_n477), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n262), .A2(G274), .A3(new_n266), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n483), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n262), .A2(new_n266), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n476), .A2(new_n485), .A3(new_n206), .A4(G45), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G270), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n400), .A2(G116), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n206), .A2(G33), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n290), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n495), .B1(new_n498), .B2(G116), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G283), .ZN(new_n500));
  INV_X1    g0300(.A(G97), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n500), .B(new_n207), .C1(G33), .C2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n502), .B(new_n289), .C1(new_n207), .C2(G116), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT20), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n254), .A2(G257), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n315), .A2(G264), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n340), .A2(G303), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n276), .B1(new_n510), .B2(new_n248), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n494), .A2(new_n506), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n246), .B1(new_n499), .B2(new_n505), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n248), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n489), .A2(new_n493), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT21), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n516), .B1(new_n513), .B2(new_n515), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n512), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n515), .A2(G200), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n515), .A2(new_n328), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n520), .A2(new_n521), .A3(new_n506), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n254), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n524));
  AND4_X1   g0324(.A1(KEYINPUT90), .A2(new_n256), .A3(G257), .A4(G1698), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT90), .B1(new_n315), .B2(G257), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n248), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n492), .A2(G264), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n528), .A2(new_n489), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT91), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n531), .A3(G179), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n528), .A2(new_n489), .A3(new_n529), .ZN(new_n533));
  AOI21_X1  g0333(.A(KEYINPUT91), .B1(new_n533), .B2(G169), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n533), .A2(new_n276), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT89), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT23), .ZN(new_n538));
  AND2_X1   g0338(.A1(KEYINPUT73), .A2(G107), .ZN(new_n539));
  NOR2_X1   g0339(.A1(KEYINPUT73), .A2(G107), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n538), .B1(new_n541), .B2(G20), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n251), .A2(G20), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G116), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n207), .A2(G107), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n538), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n537), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(KEYINPUT23), .B1(new_n444), .B2(new_n207), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n538), .A2(new_n545), .B1(new_n543), .B2(G116), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(KEYINPUT89), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT88), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n256), .A2(new_n207), .A3(G87), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT22), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT22), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n256), .A2(new_n556), .A3(new_n207), .A4(G87), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n552), .A2(new_n553), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n553), .B1(new_n552), .B2(new_n558), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT24), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n542), .A2(new_n547), .A3(new_n537), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT89), .B1(new_n549), .B2(new_n550), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n558), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT88), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT24), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n567), .A3(new_n559), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n367), .B1(new_n562), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n283), .A2(G1), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n545), .ZN(new_n571));
  XNOR2_X1  g0371(.A(new_n571), .B(KEYINPUT25), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(G107), .B2(new_n498), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n536), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n566), .A2(new_n567), .A3(new_n559), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n567), .B1(new_n566), .B2(new_n559), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n289), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n533), .A2(new_n313), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(G190), .B2(new_n533), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n573), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(G107), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(KEYINPUT6), .A3(G97), .ZN(new_n583));
  XOR2_X1   g0383(.A(G97), .B(G107), .Z(new_n584));
  OAI21_X1  g0384(.A(new_n583), .B1(new_n584), .B2(KEYINPUT6), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n585), .A2(G20), .B1(G77), .B2(new_n355), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n444), .B1(new_n341), .B2(new_n343), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n367), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n284), .A2(new_n501), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n497), .B2(new_n501), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(G244), .B(new_n314), .C1(new_n317), .C2(new_n318), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT4), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(KEYINPUT85), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n315), .A2(G250), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n500), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n593), .B1(new_n592), .B2(KEYINPUT85), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n248), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n492), .A2(G257), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n598), .A2(new_n489), .A3(new_n599), .A4(G190), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n598), .A2(new_n489), .A3(new_n599), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n591), .B(new_n600), .C1(new_n601), .C2(new_n313), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n598), .A2(new_n489), .A3(new_n599), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n246), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n588), .A2(new_n590), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n598), .A2(new_n489), .A3(new_n599), .A4(new_n276), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n207), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n325), .A2(new_n501), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n609), .B1(new_n444), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n256), .A2(new_n207), .A3(G68), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n501), .B1(new_n293), .B2(new_n295), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n611), .B(new_n612), .C1(KEYINPUT19), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n289), .ZN(new_n615));
  INV_X1    g0415(.A(new_n454), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n498), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n454), .A2(new_n284), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n615), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(G244), .B(G1698), .C1(new_n317), .C2(new_n318), .ZN(new_n620));
  OAI211_X1 g0420(.A(G238), .B(new_n314), .C1(new_n317), .C2(new_n318), .ZN(new_n621));
  NAND2_X1  g0421(.A1(G33), .A2(G116), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n248), .ZN(new_n624));
  INV_X1    g0424(.A(G45), .ZN(new_n625));
  OR3_X1    g0425(.A1(new_n625), .A2(G1), .A3(G274), .ZN(new_n626));
  INV_X1    g0426(.A(G250), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n625), .B2(G1), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n262), .A2(new_n626), .A3(new_n266), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n246), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n624), .A2(new_n276), .A3(new_n629), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n619), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n630), .A2(G200), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n614), .A2(new_n289), .B1(new_n284), .B2(new_n454), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n498), .A2(G87), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n624), .A2(G190), .A3(new_n629), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n634), .A2(new_n635), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n602), .A2(new_n607), .A3(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n523), .A2(new_n575), .A3(new_n581), .A4(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n473), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g0442(.A(new_n642), .B(KEYINPUT92), .Z(G372));
  NAND2_X1  g0443(.A1(new_n376), .A2(new_n382), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT18), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n376), .A2(new_n385), .A3(new_n382), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI22_X1  g0447(.A1(new_n282), .A2(new_n305), .B1(new_n311), .B2(new_n466), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n647), .B1(new_n648), .B2(new_n375), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n434), .A2(KEYINPUT10), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT78), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n425), .B(new_n426), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n651), .A2(new_n431), .B1(new_n652), .B2(new_n418), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n438), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT94), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT94), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n656), .B(new_n438), .C1(new_n649), .C2(new_n653), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n578), .A2(new_n573), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n519), .B1(new_n659), .B2(new_n536), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n581), .A2(new_n640), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n633), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n633), .A2(new_n638), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n663), .B1(new_n607), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n591), .B1(new_n246), .B2(new_n603), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n639), .A2(new_n666), .A3(KEYINPUT26), .A4(new_n606), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT93), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  OAI211_X1 g0469(.A(KEYINPUT93), .B(new_n663), .C1(new_n607), .C2(new_n664), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n662), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n658), .B1(new_n473), .B2(new_n672), .ZN(G369));
  AND2_X1   g0473(.A1(new_n575), .A2(new_n581), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n562), .A2(new_n568), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n574), .B1(new_n675), .B2(new_n289), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n570), .A2(new_n207), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n674), .B1(new_n676), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n575), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n506), .A2(new_n682), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n523), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n519), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n687), .B1(new_n688), .B2(new_n686), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n688), .A2(new_n682), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n674), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n659), .A2(new_n536), .A3(new_n683), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n692), .A2(new_n696), .ZN(G399));
  INV_X1    g0497(.A(new_n210), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G41), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G1), .ZN(new_n701));
  INV_X1    g0501(.A(G116), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n541), .A2(new_n325), .A3(new_n501), .A4(new_n702), .ZN(new_n703));
  OAI22_X1  g0503(.A1(new_n701), .A2(new_n703), .B1(new_n215), .B2(new_n700), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n683), .B1(new_n662), .B2(new_n671), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT96), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT29), .ZN(new_n709));
  OAI211_X1 g0509(.A(KEYINPUT96), .B(new_n683), .C1(new_n662), .C2(new_n671), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n633), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n575), .A2(new_n688), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n602), .A2(new_n607), .A3(new_n639), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n676), .B2(new_n580), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n712), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n665), .A2(new_n667), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n682), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT29), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n711), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n630), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n721), .A2(new_n493), .A3(new_n511), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n530), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n603), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT30), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n723), .B2(new_n603), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n721), .A2(G179), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n533), .A2(new_n603), .A3(new_n729), .A4(new_n515), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n725), .A2(new_n726), .A3(new_n728), .A4(new_n730), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n641), .A2(KEYINPUT31), .B1(new_n682), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n683), .A2(new_n726), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n728), .A2(new_n730), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n735), .A2(KEYINPUT95), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n735), .A2(KEYINPUT95), .B1(KEYINPUT30), .B2(new_n724), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(G330), .B1(new_n732), .B2(new_n738), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n720), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n705), .B1(new_n740), .B2(G1), .ZN(G364));
  AOI21_X1  g0541(.A(new_n213), .B1(G20), .B2(new_n246), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n742), .A2(KEYINPUT98), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(KEYINPUT98), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n244), .A2(new_n625), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n751), .B(KEYINPUT97), .Z(new_n752));
  NOR2_X1   g0552(.A1(new_n698), .A2(new_n256), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n752), .B(new_n753), .C1(G45), .C2(new_n215), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n698), .A2(new_n340), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n755), .A2(G355), .B1(new_n702), .B2(new_n698), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n750), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n283), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n206), .B1(new_n758), .B2(G45), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n699), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n745), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n207), .A2(new_n276), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(G190), .A3(new_n313), .ZN(new_n765));
  INV_X1    g0565(.A(G322), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G190), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G311), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n765), .A2(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n767), .A2(G20), .A3(new_n276), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n256), .B(new_n770), .C1(G329), .C2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n764), .A2(new_n328), .A3(G200), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n774), .A2(KEYINPUT99), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(KEYINPUT99), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(KEYINPUT33), .B(G317), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR4_X1   g0580(.A1(new_n207), .A2(new_n328), .A3(new_n313), .A4(G179), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n276), .A2(new_n313), .A3(G190), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n781), .A2(G303), .B1(new_n783), .B2(G294), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n764), .A2(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n328), .ZN(new_n786));
  NOR4_X1   g0586(.A1(new_n207), .A2(new_n313), .A3(G179), .A4(G190), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n786), .A2(G326), .B1(G283), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n773), .A2(new_n780), .A3(new_n784), .A4(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n786), .ZN(new_n790));
  INV_X1    g0590(.A(new_n787), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n790), .A2(new_n202), .B1(new_n582), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n781), .ZN(new_n793));
  INV_X1    g0593(.A(new_n783), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n793), .A2(new_n325), .B1(new_n501), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n778), .A2(G68), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n771), .A2(new_n338), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT32), .ZN(new_n799));
  INV_X1    g0599(.A(G58), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n256), .B1(new_n765), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n768), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(G77), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n796), .A2(new_n797), .A3(new_n799), .A4(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n763), .B1(new_n789), .B2(new_n804), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n757), .A2(new_n762), .A3(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n748), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n689), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n690), .A2(new_n762), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n689), .A2(G330), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(G396));
  NOR2_X1   g0611(.A1(new_n466), .A2(new_n682), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n460), .A2(new_n682), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n464), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n812), .B1(new_n814), .B2(new_n466), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n708), .A2(new_n710), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n671), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n682), .B1(new_n716), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n815), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n761), .B1(new_n821), .B2(new_n739), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n739), .B2(new_n821), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n763), .A2(new_n747), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n761), .B1(new_n824), .B2(G77), .ZN(new_n825));
  INV_X1    g0625(.A(G294), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n765), .A2(new_n826), .B1(new_n768), .B2(new_n702), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n256), .B(new_n827), .C1(G311), .C2(new_n772), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n778), .A2(G283), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n781), .A2(G107), .B1(new_n783), .B2(G97), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n791), .A2(new_n325), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(G303), .B2(new_n786), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n828), .A2(new_n829), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n256), .B1(new_n771), .B2(new_n834), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n793), .A2(new_n202), .B1(new_n791), .B2(new_n285), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n835), .B(new_n836), .C1(G58), .C2(new_n783), .ZN(new_n837));
  INV_X1    g0637(.A(new_n765), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n838), .A2(G143), .B1(new_n802), .B2(G159), .ZN(new_n839));
  INV_X1    g0639(.A(G137), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n839), .B1(new_n840), .B2(new_n790), .C1(new_n777), .C2(new_n389), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n837), .B1(new_n842), .B2(KEYINPUT34), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT34), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n833), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n825), .B1(new_n846), .B2(new_n745), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n815), .B2(new_n747), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n823), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G384));
  NOR2_X1   g0650(.A1(new_n758), .A2(new_n206), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT40), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n362), .A2(KEYINPUT84), .A3(new_n371), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n384), .B(new_n386), .C1(new_n853), .C2(new_n372), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n368), .A2(KEYINPUT16), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n333), .B1(new_n359), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n680), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n381), .B(new_n680), .C1(new_n380), .C2(new_n276), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n856), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n861), .B1(new_n863), .B2(new_n360), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n377), .A2(new_n379), .A3(new_n862), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT37), .B1(new_n370), .B2(new_n330), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n860), .A2(KEYINPUT38), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT105), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n867), .B1(new_n854), .B2(new_n859), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(KEYINPUT105), .A3(KEYINPUT38), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT104), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n377), .A2(new_n379), .A3(new_n857), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n360), .A2(KEYINPUT103), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT103), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n370), .A2(new_n878), .A3(new_n330), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(new_n644), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT37), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n865), .A2(new_n866), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n645), .A2(new_n362), .A3(new_n371), .A4(new_n646), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n881), .A2(new_n882), .B1(new_n876), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n875), .B1(new_n884), .B2(KEYINPUT38), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n377), .A2(new_n379), .A3(new_n857), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n887), .A2(new_n644), .A3(new_n879), .A4(new_n877), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n888), .A2(KEYINPUT37), .B1(new_n865), .B2(new_n866), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n883), .A2(new_n876), .ZN(new_n890));
  OAI211_X1 g0690(.A(KEYINPUT104), .B(new_n886), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n874), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n641), .A2(KEYINPUT31), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n731), .A2(new_n682), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n735), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n734), .B1(new_n897), .B2(new_n725), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n305), .ZN(new_n901));
  INV_X1    g0701(.A(new_n277), .ZN(new_n902));
  INV_X1    g0702(.A(new_n281), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n280), .B1(new_n273), .B2(new_n274), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n901), .B(new_n682), .C1(new_n905), .C2(new_n311), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n901), .A2(new_n682), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n310), .B(new_n907), .C1(new_n282), .C2(new_n305), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n900), .A2(new_n815), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n852), .B1(new_n893), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT38), .B1(new_n860), .B2(new_n868), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n886), .B(new_n867), .C1(new_n854), .C2(new_n859), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT102), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n872), .A2(KEYINPUT102), .A3(KEYINPUT38), .ZN(new_n917));
  NOR4_X1   g0717(.A1(new_n916), .A2(new_n910), .A3(KEYINPUT40), .A4(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(G330), .B1(new_n912), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n472), .A2(G330), .A3(new_n900), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n921), .A2(KEYINPUT106), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n885), .A2(new_n891), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n871), .B2(new_n873), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT40), .B1(new_n924), .B2(new_n910), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n915), .B1(new_n872), .B2(KEYINPUT38), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n858), .B1(new_n387), .B2(new_n375), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n886), .B1(new_n927), .B2(new_n867), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n917), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n911), .A2(new_n929), .A3(new_n852), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n925), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(new_n472), .A3(new_n900), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n921), .A2(KEYINPUT106), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n922), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n812), .B(KEYINPUT101), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n819), .B2(new_n815), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n938), .A2(new_n929), .A3(new_n930), .A4(new_n909), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n647), .A2(new_n680), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT39), .ZN(new_n941));
  AND4_X1   g0741(.A1(KEYINPUT105), .A2(new_n860), .A3(KEYINPUT38), .A4(new_n868), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT105), .B1(new_n872), .B2(KEYINPUT38), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n941), .B1(new_n944), .B2(new_n923), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT39), .B1(new_n916), .B2(new_n917), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n306), .A2(new_n683), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n939), .B(new_n940), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n711), .A2(new_n472), .A3(new_n719), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n658), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n949), .B(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n851), .B1(new_n935), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n952), .B2(new_n935), .ZN(new_n954));
  NOR4_X1   g0754(.A1(new_n335), .A2(new_n336), .A3(new_n215), .A4(new_n297), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n202), .B2(G68), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n956), .A2(new_n206), .A3(G13), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT100), .Z(new_n958));
  INV_X1    g0758(.A(KEYINPUT36), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n214), .A2(G116), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(new_n585), .B2(KEYINPUT35), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(KEYINPUT35), .B2(new_n585), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n958), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n959), .B2(new_n962), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n954), .A2(new_n964), .ZN(G367));
  OAI22_X1  g0765(.A1(new_n765), .A2(new_n389), .B1(new_n768), .B2(new_n202), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n340), .B(new_n966), .C1(G137), .C2(new_n772), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n778), .A2(G159), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n786), .A2(G143), .B1(G77), .B2(new_n787), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n794), .A2(new_n285), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G58), .B2(new_n781), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n967), .A2(new_n968), .A3(new_n969), .A4(new_n971), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n790), .A2(new_n769), .B1(new_n501), .B2(new_n791), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(new_n444), .B2(new_n783), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n781), .A2(KEYINPUT46), .A3(G116), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n256), .B1(new_n838), .B2(G303), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n802), .A2(G283), .B1(new_n772), .B2(G317), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n974), .A2(new_n975), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT46), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n793), .B2(new_n702), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n980), .A2(KEYINPUT108), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(KEYINPUT108), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n981), .B(new_n982), .C1(new_n826), .C2(new_n777), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n972), .B1(new_n978), .B2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT109), .Z(new_n985));
  OR2_X1    g0785(.A1(new_n985), .A2(KEYINPUT47), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(KEYINPUT47), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n986), .A2(new_n745), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n750), .B1(new_n698), .B2(new_n616), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n753), .A2(new_n236), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n762), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n635), .A2(new_n636), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n682), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n639), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n633), .B2(new_n993), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n988), .B(new_n991), .C1(new_n807), .C2(new_n995), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n602), .B(new_n607), .C1(new_n591), .C2(new_n683), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n666), .A2(new_n606), .A3(new_n682), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n696), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT44), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n696), .A2(new_n999), .ZN(new_n1002));
  XOR2_X1   g0802(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n1003));
  XNOR2_X1  g0803(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n692), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n694), .B1(new_n685), .B2(new_n693), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(new_n691), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n740), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n740), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n699), .B(KEYINPUT41), .Z(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n760), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n674), .A2(new_n693), .A3(new_n999), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1015), .A2(KEYINPUT42), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n607), .B1(new_n575), .B2(new_n997), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n1015), .A2(KEYINPUT42), .B1(new_n683), .B2(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n1016), .A2(new_n1018), .B1(KEYINPUT43), .B2(new_n995), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n995), .A2(KEYINPUT43), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n999), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n692), .A2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1021), .B(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n996), .B1(new_n1014), .B2(new_n1024), .ZN(G387));
  OR2_X1    g0825(.A1(new_n685), .A2(new_n807), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n753), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n233), .B2(G45), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n703), .B2(new_n755), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n391), .A2(new_n202), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT50), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n625), .B1(new_n285), .B2(new_n297), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n1031), .A2(new_n703), .A3(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n1029), .A2(new_n1033), .B1(G107), .B2(new_n210), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n762), .B1(new_n1034), .B2(new_n749), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT110), .Z(new_n1036));
  AOI22_X1  g0836(.A1(new_n838), .A2(G317), .B1(new_n802), .B2(G303), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n766), .B2(new_n790), .C1(new_n777), .C2(new_n769), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT48), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n781), .A2(G294), .B1(new_n783), .B2(G283), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT49), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n791), .A2(new_n702), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n256), .B(new_n1047), .C1(G326), .C2(new_n772), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  XOR2_X1   g0849(.A(KEYINPUT111), .B(G150), .Z(new_n1050));
  OAI22_X1  g0850(.A1(new_n765), .A2(new_n202), .B1(new_n1050), .B2(new_n771), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n340), .B(new_n1051), .C1(G68), .C2(new_n802), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n778), .A2(new_n391), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n786), .A2(G159), .B1(G97), .B2(new_n787), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n793), .A2(new_n297), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n616), .B2(new_n783), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n763), .B1(new_n1049), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1036), .A2(new_n1058), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1009), .A2(new_n760), .B1(new_n1026), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1010), .A2(new_n699), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n740), .A2(new_n1009), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(G393));
  OR2_X1    g0863(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(KEYINPUT112), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1066), .B(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1010), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n699), .B(new_n1064), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G317), .A2(new_n786), .B1(new_n838), .B2(G311), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT52), .ZN(new_n1072));
  INV_X1    g0872(.A(G283), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n793), .A2(new_n1073), .B1(new_n791), .B2(new_n582), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G116), .B2(new_n783), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n340), .B1(new_n768), .B2(new_n826), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G322), .B2(new_n772), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1072), .B(new_n1078), .C1(G303), .C2(new_n778), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n256), .B1(new_n768), .B2(new_n331), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1080), .B(new_n831), .C1(G77), .C2(new_n783), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n202), .B2(new_n777), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G150), .A2(new_n786), .B1(new_n838), .B2(G159), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT51), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n781), .A2(G68), .B1(new_n772), .B2(G143), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT113), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1082), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1079), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n763), .B1(new_n1088), .B2(KEYINPUT114), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(KEYINPUT114), .B2(new_n1088), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n749), .B1(new_n501), .B2(new_n210), .C1(new_n241), .C2(new_n1027), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1090), .A2(new_n761), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n748), .B2(new_n1022), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n1068), .B2(new_n760), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1070), .A2(new_n1094), .ZN(G390));
  AOI21_X1  g0895(.A(new_n936), .B1(new_n718), .B2(new_n815), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n909), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n948), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n924), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n948), .B1(new_n937), .B2(new_n1097), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1099), .B1(new_n947), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n815), .A2(G330), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n909), .C1(new_n732), .C2(new_n898), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1104), .A2(KEYINPUT115), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(KEYINPUT39), .B1(new_n874), .B2(new_n892), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n941), .B1(new_n929), .B2(new_n930), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1100), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n924), .A2(new_n1098), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n736), .A2(new_n737), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n733), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1102), .B1(new_n896), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n900), .A2(new_n1103), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT115), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n909), .B(new_n1113), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1109), .A2(new_n1110), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1106), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n947), .A2(new_n746), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n761), .B1(new_n824), .B2(new_n391), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n765), .A2(new_n702), .B1(new_n768), .B2(new_n501), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n256), .B(new_n1122), .C1(G294), .C2(new_n772), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n778), .A2(new_n444), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n781), .A2(G87), .B1(new_n787), .B2(G68), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n786), .A2(G283), .B1(G77), .B2(new_n783), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n793), .A2(new_n1050), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT53), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n840), .B2(new_n777), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n786), .A2(G128), .B1(G159), .B2(new_n783), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n838), .A2(G132), .B1(G125), .B2(new_n772), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT54), .B(G143), .Z(new_n1133));
  AOI21_X1  g0933(.A(new_n340), .B1(new_n802), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n787), .A2(G50), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1127), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1121), .B1(new_n1137), .B2(new_n745), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1119), .A2(new_n760), .B1(new_n1120), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n950), .A2(new_n920), .A3(new_n658), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1114), .A2(new_n1097), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1103), .B(new_n909), .C1(new_n732), .C2(new_n738), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n936), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n717), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n683), .B(new_n815), .C1(new_n662), .C2(new_n1144), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1104), .B1(new_n1113), .B2(new_n909), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1141), .A2(new_n1146), .B1(new_n1147), .B2(new_n938), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1140), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n1106), .B2(new_n1118), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1117), .B(new_n1149), .C1(new_n1101), .C2(new_n1105), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n699), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1139), .A2(new_n1153), .ZN(G378));
  INV_X1    g0954(.A(new_n1140), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT118), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1152), .A2(KEYINPUT118), .A3(new_n1155), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n436), .A2(new_n438), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n857), .B1(new_n398), .B2(new_n401), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1162), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g0969(.A(G330), .B(new_n1169), .C1(new_n912), .C2(new_n918), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1169), .B1(new_n932), .B2(G330), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n949), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n947), .A2(new_n948), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n939), .A2(new_n940), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1169), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n919), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1178), .A3(new_n1170), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1173), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1158), .A2(new_n1159), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT57), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1158), .A2(new_n1180), .A3(KEYINPUT57), .A4(new_n1159), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1183), .A2(new_n699), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1180), .A2(new_n760), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1177), .A2(new_n746), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n761), .B1(new_n824), .B2(G50), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n777), .A2(new_n501), .B1(new_n454), .B2(new_n768), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT116), .Z(new_n1190));
  OAI22_X1  g0990(.A1(new_n790), .A2(new_n702), .B1(new_n800), .B2(new_n791), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n256), .A2(G41), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n1073), .B2(new_n771), .C1(new_n582), .C2(new_n765), .ZN(new_n1193));
  NOR4_X1   g0993(.A1(new_n1191), .A2(new_n1193), .A3(new_n970), .A4(new_n1055), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT58), .B1(new_n1190), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1190), .A2(KEYINPUT58), .A3(new_n1194), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(G128), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n765), .A2(new_n1198), .B1(new_n768), .B2(new_n840), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G150), .B2(new_n783), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n786), .A2(G125), .B1(new_n781), .B2(new_n1133), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(new_n777), .C2(new_n834), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1202), .A2(KEYINPUT59), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(KEYINPUT59), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n787), .A2(G159), .ZN(new_n1205));
  AOI211_X1 g1005(.A(G33), .B(G41), .C1(new_n772), .C2(G124), .ZN(new_n1206));
  AND4_X1   g1006(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  AOI211_X1 g1007(.A(G50), .B(new_n1192), .C1(new_n251), .C2(new_n478), .ZN(new_n1208));
  OR4_X1    g1008(.A1(new_n1195), .A2(new_n1197), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1188), .B1(new_n1209), .B2(new_n745), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1187), .A2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT117), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1186), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1185), .A2(new_n1214), .ZN(G375));
  OAI21_X1  g1015(.A(new_n761), .B1(new_n824), .B2(G68), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n778), .A2(new_n1133), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n768), .A2(new_n389), .B1(new_n771), .B2(new_n1198), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n340), .B(new_n1218), .C1(G137), .C2(new_n838), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n786), .A2(G132), .B1(G58), .B2(new_n787), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n781), .A2(G159), .B1(new_n783), .B2(G50), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1217), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n777), .A2(new_n702), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n786), .A2(G294), .B1(G97), .B2(new_n781), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n838), .A2(G283), .B1(new_n802), .B2(new_n444), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n256), .B1(new_n772), .B2(G303), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n616), .A2(new_n783), .B1(new_n787), .B2(G77), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1222), .B1(new_n1223), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1216), .B1(new_n1229), .B2(new_n745), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n909), .B2(new_n747), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1148), .B2(new_n759), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1012), .B(KEYINPUT119), .Z(new_n1233));
  NOR2_X1   g1033(.A1(new_n1149), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1140), .A2(new_n1148), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1232), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(G381));
  XNOR2_X1  g1037(.A(G375), .B(KEYINPUT121), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT120), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1139), .A2(new_n1153), .A3(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1239), .B1(new_n1139), .B2(new_n1153), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(G390), .A2(G387), .ZN(new_n1243));
  NOR4_X1   g1043(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1238), .A2(new_n1245), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT122), .ZN(G407));
  INV_X1    g1047(.A(G213), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1242), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(G343), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1248), .B1(new_n1238), .B2(new_n1252), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1246), .A2(KEYINPUT122), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1246), .A2(KEYINPUT122), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1253), .B1(new_n1254), .B2(new_n1255), .ZN(G409));
  INV_X1    g1056(.A(new_n1243), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G390), .A2(G387), .ZN(new_n1258));
  XOR2_X1   g1058(.A(G393), .B(G396), .Z(new_n1259));
  OR2_X1    g1059(.A1(new_n1259), .A2(KEYINPUT126), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1257), .A2(new_n1258), .A3(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(KEYINPUT126), .A3(new_n1259), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(KEYINPUT126), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1257), .A2(new_n1263), .A3(new_n1260), .A4(new_n1258), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1250), .A2(G2897), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT123), .ZN(new_n1267));
  AOI21_X1  g1067(.A(KEYINPUT60), .B1(new_n1140), .B2(new_n1148), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1267), .B1(new_n1268), .B2(new_n1149), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1140), .A2(new_n1148), .A3(KEYINPUT60), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1270), .A2(new_n699), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1268), .A2(new_n1149), .A3(new_n1267), .ZN(new_n1273));
  OAI21_X1  g1073(.A(KEYINPUT124), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  OR3_X1    g1074(.A1(new_n1268), .A2(new_n1149), .A3(new_n1267), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT124), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1275), .A2(new_n1269), .A3(new_n1276), .A4(new_n1271), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1232), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n849), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1278), .A2(G384), .A3(new_n1279), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1266), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G384), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n849), .B(new_n1232), .C1(new_n1274), .C2(new_n1277), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1266), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1284), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1283), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n700), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1213), .B1(new_n1289), .B2(new_n1184), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1211), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1186), .B(new_n1291), .C1(new_n1181), .C2(new_n1233), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n1290), .A2(G378), .B1(new_n1242), .B2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1288), .B1(new_n1293), .B2(new_n1250), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1185), .A2(G378), .A3(new_n1214), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1242), .A2(new_n1292), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT62), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1297), .A2(new_n1298), .A3(new_n1251), .A4(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT61), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1294), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  XOR2_X1   g1102(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1303));
  AOI21_X1  g1103(.A(new_n1250), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(new_n1304), .B2(new_n1299), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1265), .B1(new_n1302), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1304), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT61), .B1(new_n1307), .B2(new_n1288), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1304), .A2(new_n1299), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1304), .A2(KEYINPUT63), .A3(new_n1299), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1308), .A2(new_n1311), .A3(new_n1312), .A4(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1306), .A2(new_n1314), .ZN(G405));
  OAI21_X1  g1115(.A(new_n1295), .B1(new_n1290), .B2(new_n1249), .ZN(new_n1316));
  OR2_X1    g1116(.A1(new_n1316), .A2(new_n1299), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1299), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1265), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1312), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(G402));
endmodule


