

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U323 ( .A(KEYINPUT94), .B(KEYINPUT26), .ZN(n455) );
  XOR2_X1 U324 ( .A(G155GAT), .B(G148GAT), .Z(n291) );
  INV_X1 U325 ( .A(KEYINPUT46), .ZN(n360) );
  XNOR2_X1 U326 ( .A(n366), .B(KEYINPUT111), .ZN(n367) );
  XNOR2_X1 U327 ( .A(KEYINPUT31), .B(KEYINPUT76), .ZN(n347) );
  XNOR2_X1 U328 ( .A(n420), .B(n291), .ZN(n421) );
  XNOR2_X1 U329 ( .A(n422), .B(n421), .ZN(n426) );
  INV_X1 U330 ( .A(KEYINPUT101), .ZN(n472) );
  XNOR2_X1 U331 ( .A(n399), .B(n357), .ZN(n358) );
  XNOR2_X1 U332 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U333 ( .A(n456), .B(n455), .ZN(n570) );
  XNOR2_X1 U334 ( .A(n475), .B(n474), .ZN(n522) );
  XNOR2_X1 U335 ( .A(n452), .B(n451), .ZN(n565) );
  INV_X1 U336 ( .A(G43GAT), .ZN(n477) );
  XNOR2_X1 U337 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n453) );
  XNOR2_X1 U338 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U339 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(n480), .B(n479), .ZN(G1330GAT) );
  INV_X1 U341 ( .A(KEYINPUT120), .ZN(n452) );
  XOR2_X1 U342 ( .A(KEYINPUT81), .B(KEYINPUT65), .Z(n293) );
  NAND2_X1 U343 ( .A1(G232GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U344 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U345 ( .A(n294), .B(KEYINPUT11), .Z(n298) );
  XNOR2_X1 U346 ( .A(G29GAT), .B(G134GAT), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n295), .B(KEYINPUT80), .ZN(n409) );
  XNOR2_X1 U348 ( .A(G36GAT), .B(G190GAT), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n296), .B(KEYINPUT82), .ZN(n380) );
  XNOR2_X1 U350 ( .A(n409), .B(n380), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n305) );
  XOR2_X1 U352 ( .A(G106GAT), .B(KEYINPUT9), .Z(n300) );
  XNOR2_X1 U353 ( .A(KEYINPUT83), .B(KEYINPUT10), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U355 ( .A(n301), .B(KEYINPUT79), .Z(n303) );
  XOR2_X1 U356 ( .A(G50GAT), .B(G162GAT), .Z(n420) );
  XNOR2_X1 U357 ( .A(n420), .B(G218GAT), .ZN(n302) );
  XNOR2_X1 U358 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U359 ( .A(n305), .B(n304), .Z(n311) );
  XOR2_X1 U360 ( .A(G43GAT), .B(KEYINPUT8), .Z(n307) );
  XNOR2_X1 U361 ( .A(KEYINPUT7), .B(KEYINPUT70), .ZN(n306) );
  XNOR2_X1 U362 ( .A(n307), .B(n306), .ZN(n344) );
  XOR2_X1 U363 ( .A(G92GAT), .B(KEYINPUT78), .Z(n309) );
  XNOR2_X1 U364 ( .A(G99GAT), .B(G85GAT), .ZN(n308) );
  XNOR2_X1 U365 ( .A(n309), .B(n308), .ZN(n348) );
  XNOR2_X1 U366 ( .A(n344), .B(n348), .ZN(n310) );
  XNOR2_X1 U367 ( .A(n311), .B(n310), .ZN(n562) );
  XOR2_X1 U368 ( .A(KEYINPUT75), .B(KEYINPUT13), .Z(n313) );
  XNOR2_X1 U369 ( .A(G71GAT), .B(G57GAT), .ZN(n312) );
  XNOR2_X1 U370 ( .A(n313), .B(n312), .ZN(n354) );
  XOR2_X1 U371 ( .A(G1GAT), .B(G127GAT), .Z(n314) );
  XOR2_X1 U372 ( .A(G155GAT), .B(n314), .Z(n402) );
  XOR2_X1 U373 ( .A(n354), .B(n402), .Z(n327) );
  XOR2_X1 U374 ( .A(KEYINPUT14), .B(KEYINPUT84), .Z(n316) );
  XNOR2_X1 U375 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n315) );
  XNOR2_X1 U376 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U377 ( .A(KEYINPUT12), .B(G78GAT), .Z(n318) );
  NAND2_X1 U378 ( .A1(G231GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U380 ( .A(n320), .B(n319), .Z(n325) );
  XOR2_X1 U381 ( .A(G15GAT), .B(G22GAT), .Z(n322) );
  XNOR2_X1 U382 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n322), .B(n321), .ZN(n343) );
  XNOR2_X1 U384 ( .A(G8GAT), .B(G183GAT), .ZN(n323) );
  XNOR2_X1 U385 ( .A(n323), .B(G211GAT), .ZN(n389) );
  XNOR2_X1 U386 ( .A(n343), .B(n389), .ZN(n324) );
  XNOR2_X1 U387 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U388 ( .A(n327), .B(n326), .Z(n580) );
  XOR2_X1 U389 ( .A(KEYINPUT109), .B(n580), .Z(n543) );
  XOR2_X1 U390 ( .A(G113GAT), .B(G50GAT), .Z(n329) );
  XNOR2_X1 U391 ( .A(G29GAT), .B(G36GAT), .ZN(n328) );
  XNOR2_X1 U392 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U393 ( .A(KEYINPUT74), .B(G8GAT), .Z(n331) );
  XNOR2_X1 U394 ( .A(G141GAT), .B(G1GAT), .ZN(n330) );
  XNOR2_X1 U395 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U396 ( .A(n333), .B(n332), .Z(n338) );
  XOR2_X1 U397 ( .A(KEYINPUT30), .B(G197GAT), .Z(n335) );
  NAND2_X1 U398 ( .A1(G229GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U399 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U400 ( .A(KEYINPUT29), .B(n336), .ZN(n337) );
  XNOR2_X1 U401 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U402 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n340) );
  XNOR2_X1 U403 ( .A(G169GAT), .B(KEYINPUT73), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U405 ( .A(n342), .B(n341), .Z(n346) );
  XNOR2_X1 U406 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U407 ( .A(n346), .B(n345), .Z(n553) );
  INV_X1 U408 ( .A(n553), .ZN(n572) );
  XNOR2_X1 U409 ( .A(n348), .B(n347), .ZN(n351) );
  XNOR2_X1 U410 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n349) );
  XOR2_X1 U411 ( .A(G176GAT), .B(G64GAT), .Z(n383) );
  XNOR2_X1 U412 ( .A(n349), .B(n383), .ZN(n350) );
  XOR2_X1 U413 ( .A(n351), .B(n350), .Z(n356) );
  XOR2_X1 U414 ( .A(G204GAT), .B(KEYINPUT77), .Z(n353) );
  XNOR2_X1 U415 ( .A(G106GAT), .B(G78GAT), .ZN(n352) );
  XNOR2_X1 U416 ( .A(n353), .B(n352), .ZN(n428) );
  XNOR2_X1 U417 ( .A(n354), .B(n428), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n359) );
  XOR2_X1 U419 ( .A(G120GAT), .B(G148GAT), .Z(n399) );
  AND2_X1 U420 ( .A1(G230GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n369) );
  XNOR2_X1 U422 ( .A(KEYINPUT41), .B(n369), .ZN(n557) );
  NAND2_X1 U423 ( .A1(n572), .A2(n557), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n361), .B(n360), .ZN(n362) );
  NOR2_X1 U425 ( .A1(n543), .A2(n362), .ZN(n364) );
  INV_X1 U426 ( .A(KEYINPUT110), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n365) );
  NOR2_X1 U428 ( .A1(n562), .A2(n365), .ZN(n368) );
  INV_X1 U429 ( .A(KEYINPUT47), .ZN(n366) );
  XNOR2_X1 U430 ( .A(n368), .B(n367), .ZN(n376) );
  XOR2_X1 U431 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n371) );
  XNOR2_X1 U432 ( .A(n562), .B(KEYINPUT36), .ZN(n582) );
  NAND2_X1 U433 ( .A1(n580), .A2(n582), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n371), .B(n370), .ZN(n372) );
  NAND2_X1 U435 ( .A1(n369), .A2(n372), .ZN(n373) );
  XOR2_X1 U436 ( .A(KEYINPUT112), .B(n373), .Z(n374) );
  NAND2_X1 U437 ( .A1(n374), .A2(n553), .ZN(n375) );
  NAND2_X1 U438 ( .A1(n376), .A2(n375), .ZN(n378) );
  XNOR2_X1 U439 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n378), .B(n377), .ZN(n532) );
  XNOR2_X1 U441 ( .A(G197GAT), .B(G218GAT), .ZN(n379) );
  XNOR2_X1 U442 ( .A(n379), .B(KEYINPUT21), .ZN(n427) );
  XOR2_X1 U443 ( .A(n380), .B(KEYINPUT93), .Z(n382) );
  NAND2_X1 U444 ( .A1(G226GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n382), .B(n381), .ZN(n386) );
  XNOR2_X1 U446 ( .A(G92GAT), .B(G204GAT), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U448 ( .A(n386), .B(n385), .Z(n391) );
  XOR2_X1 U449 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n388) );
  XNOR2_X1 U450 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n388), .B(n387), .ZN(n436) );
  XNOR2_X1 U452 ( .A(n436), .B(n389), .ZN(n390) );
  XNOR2_X1 U453 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U454 ( .A(n427), .B(n392), .ZN(n524) );
  NOR2_X1 U455 ( .A1(n532), .A2(n524), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n393), .B(KEYINPUT54), .ZN(n414) );
  XOR2_X1 U457 ( .A(KEYINPUT6), .B(KEYINPUT89), .Z(n395) );
  XNOR2_X1 U458 ( .A(KEYINPUT4), .B(KEYINPUT90), .ZN(n394) );
  XNOR2_X1 U459 ( .A(n395), .B(n394), .ZN(n413) );
  XOR2_X1 U460 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n397) );
  XNOR2_X1 U461 ( .A(KEYINPUT91), .B(G57GAT), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U463 ( .A(n398), .B(G85GAT), .Z(n401) );
  XNOR2_X1 U464 ( .A(n399), .B(G162GAT), .ZN(n400) );
  XNOR2_X1 U465 ( .A(n401), .B(n400), .ZN(n406) );
  XOR2_X1 U466 ( .A(G113GAT), .B(KEYINPUT0), .Z(n435) );
  XOR2_X1 U467 ( .A(n435), .B(n402), .Z(n404) );
  NAND2_X1 U468 ( .A1(G225GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U469 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U470 ( .A(n406), .B(n405), .Z(n411) );
  XOR2_X1 U471 ( .A(KEYINPUT2), .B(KEYINPUT88), .Z(n408) );
  XNOR2_X1 U472 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n407) );
  XNOR2_X1 U473 ( .A(n408), .B(n407), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n409), .B(n417), .ZN(n410) );
  XNOR2_X1 U475 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U476 ( .A(n413), .B(n412), .Z(n462) );
  XNOR2_X1 U477 ( .A(KEYINPUT92), .B(n462), .ZN(n533) );
  AND2_X1 U478 ( .A1(n414), .A2(n533), .ZN(n416) );
  INV_X1 U479 ( .A(KEYINPUT64), .ZN(n415) );
  XNOR2_X1 U480 ( .A(n416), .B(n415), .ZN(n571) );
  XOR2_X1 U481 ( .A(KEYINPUT23), .B(n417), .Z(n419) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U483 ( .A(n419), .B(n418), .ZN(n422) );
  XOR2_X1 U484 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n424) );
  XNOR2_X1 U485 ( .A(G22GAT), .B(G211GAT), .ZN(n423) );
  XNOR2_X1 U486 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U487 ( .A(n426), .B(n425), .Z(n430) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n464) );
  NOR2_X1 U490 ( .A1(n571), .A2(n464), .ZN(n432) );
  XNOR2_X1 U491 ( .A(KEYINPUT119), .B(KEYINPUT55), .ZN(n431) );
  XNOR2_X1 U492 ( .A(n432), .B(n431), .ZN(n450) );
  XOR2_X1 U493 ( .A(G120GAT), .B(G127GAT), .Z(n434) );
  XNOR2_X1 U494 ( .A(G43GAT), .B(G99GAT), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n449) );
  XOR2_X1 U496 ( .A(n436), .B(n435), .Z(n438) );
  XNOR2_X1 U497 ( .A(G134GAT), .B(G190GAT), .ZN(n437) );
  XNOR2_X1 U498 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U499 ( .A(KEYINPUT87), .B(KEYINPUT20), .Z(n440) );
  NAND2_X1 U500 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U502 ( .A(n442), .B(n441), .Z(n447) );
  XOR2_X1 U503 ( .A(G176GAT), .B(G183GAT), .Z(n444) );
  XNOR2_X1 U504 ( .A(G15GAT), .B(G71GAT), .ZN(n443) );
  XNOR2_X1 U505 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U506 ( .A(n445), .B(KEYINPUT86), .ZN(n446) );
  XNOR2_X1 U507 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U508 ( .A(n449), .B(n448), .ZN(n526) );
  INV_X1 U509 ( .A(n526), .ZN(n534) );
  NAND2_X1 U510 ( .A1(n450), .A2(n534), .ZN(n451) );
  NAND2_X1 U511 ( .A1(n565), .A2(n562), .ZN(n454) );
  INV_X1 U512 ( .A(n580), .ZN(n487) );
  XOR2_X1 U513 ( .A(KEYINPUT27), .B(n524), .Z(n466) );
  INV_X1 U514 ( .A(n466), .ZN(n457) );
  NAND2_X1 U515 ( .A1(n526), .A2(n464), .ZN(n456) );
  NOR2_X1 U516 ( .A1(n457), .A2(n570), .ZN(n552) );
  NOR2_X1 U517 ( .A1(n524), .A2(n526), .ZN(n458) );
  NOR2_X1 U518 ( .A1(n464), .A2(n458), .ZN(n459) );
  XOR2_X1 U519 ( .A(KEYINPUT25), .B(n459), .Z(n460) );
  NOR2_X1 U520 ( .A1(n552), .A2(n460), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n461), .B(KEYINPUT95), .ZN(n463) );
  NAND2_X1 U522 ( .A1(n463), .A2(n462), .ZN(n469) );
  XNOR2_X1 U523 ( .A(n464), .B(KEYINPUT67), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n465), .B(KEYINPUT28), .ZN(n529) );
  NAND2_X1 U525 ( .A1(n529), .A2(n466), .ZN(n536) );
  NOR2_X1 U526 ( .A1(n533), .A2(n536), .ZN(n467) );
  NAND2_X1 U527 ( .A1(n467), .A2(n526), .ZN(n468) );
  NAND2_X1 U528 ( .A1(n469), .A2(n468), .ZN(n490) );
  NAND2_X1 U529 ( .A1(n487), .A2(n490), .ZN(n470) );
  XOR2_X1 U530 ( .A(KEYINPUT100), .B(n470), .Z(n471) );
  NAND2_X1 U531 ( .A1(n471), .A2(n582), .ZN(n475) );
  XOR2_X1 U532 ( .A(KEYINPUT102), .B(KEYINPUT37), .Z(n473) );
  NAND2_X1 U533 ( .A1(n572), .A2(n369), .ZN(n492) );
  NOR2_X1 U534 ( .A1(n522), .A2(n492), .ZN(n476) );
  XOR2_X1 U535 ( .A(KEYINPUT38), .B(n476), .Z(n508) );
  NOR2_X1 U536 ( .A1(n508), .A2(n526), .ZN(n480) );
  XNOR2_X1 U537 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n478) );
  NAND2_X1 U538 ( .A1(n565), .A2(n543), .ZN(n482) );
  XNOR2_X1 U539 ( .A(G183GAT), .B(KEYINPUT122), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n482), .B(n481), .ZN(G1350GAT) );
  XNOR2_X1 U541 ( .A(KEYINPUT106), .B(n557), .ZN(n539) );
  NAND2_X1 U542 ( .A1(n539), .A2(n565), .ZN(n486) );
  XOR2_X1 U543 ( .A(G176GAT), .B(KEYINPUT121), .Z(n484) );
  XOR2_X1 U544 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(G1349GAT) );
  NOR2_X1 U547 ( .A1(n562), .A2(n487), .ZN(n488) );
  XOR2_X1 U548 ( .A(KEYINPUT16), .B(n488), .Z(n489) );
  XNOR2_X1 U549 ( .A(n489), .B(KEYINPUT85), .ZN(n491) );
  NAND2_X1 U550 ( .A1(n491), .A2(n490), .ZN(n511) );
  OR2_X1 U551 ( .A1(n492), .A2(n511), .ZN(n500) );
  NOR2_X1 U552 ( .A1(n533), .A2(n500), .ZN(n494) );
  XNOR2_X1 U553 ( .A(KEYINPUT34), .B(KEYINPUT96), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U555 ( .A(G1GAT), .B(n495), .Z(G1324GAT) );
  NOR2_X1 U556 ( .A1(n524), .A2(n500), .ZN(n496) );
  XOR2_X1 U557 ( .A(G8GAT), .B(n496), .Z(G1325GAT) );
  NOR2_X1 U558 ( .A1(n526), .A2(n500), .ZN(n498) );
  XNOR2_X1 U559 ( .A(KEYINPUT97), .B(KEYINPUT35), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U561 ( .A(G15GAT), .B(n499), .Z(G1326GAT) );
  NOR2_X1 U562 ( .A1(n529), .A2(n500), .ZN(n502) );
  XNOR2_X1 U563 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U565 ( .A(G22GAT), .B(n503), .ZN(G1327GAT) );
  NOR2_X1 U566 ( .A1(n508), .A2(n533), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  NOR2_X1 U569 ( .A1(n508), .A2(n524), .ZN(n507) );
  XNOR2_X1 U570 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(G1329GAT) );
  XNOR2_X1 U572 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n510) );
  NOR2_X1 U573 ( .A1(n529), .A2(n508), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(G1331GAT) );
  NAND2_X1 U575 ( .A1(n539), .A2(n553), .ZN(n521) );
  NOR2_X1 U576 ( .A1(n511), .A2(n521), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(KEYINPUT107), .ZN(n517) );
  NOR2_X1 U578 ( .A1(n533), .A2(n517), .ZN(n513) );
  XOR2_X1 U579 ( .A(KEYINPUT42), .B(n513), .Z(n514) );
  XNOR2_X1 U580 ( .A(G57GAT), .B(n514), .ZN(G1332GAT) );
  NOR2_X1 U581 ( .A1(n524), .A2(n517), .ZN(n515) );
  XOR2_X1 U582 ( .A(G64GAT), .B(n515), .Z(G1333GAT) );
  NOR2_X1 U583 ( .A1(n526), .A2(n517), .ZN(n516) );
  XOR2_X1 U584 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  NOR2_X1 U585 ( .A1(n529), .A2(n517), .ZN(n519) );
  XNOR2_X1 U586 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n518) );
  XNOR2_X1 U587 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(n520), .ZN(G1335GAT) );
  OR2_X1 U589 ( .A1(n522), .A2(n521), .ZN(n528) );
  NOR2_X1 U590 ( .A1(n533), .A2(n528), .ZN(n523) );
  XOR2_X1 U591 ( .A(G85GAT), .B(n523), .Z(G1336GAT) );
  NOR2_X1 U592 ( .A1(n524), .A2(n528), .ZN(n525) );
  XOR2_X1 U593 ( .A(G92GAT), .B(n525), .Z(G1337GAT) );
  NOR2_X1 U594 ( .A1(n526), .A2(n528), .ZN(n527) );
  XOR2_X1 U595 ( .A(G99GAT), .B(n527), .Z(G1338GAT) );
  NOR2_X1 U596 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U597 ( .A(KEYINPUT44), .B(n530), .Z(n531) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NOR2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n551) );
  NAND2_X1 U600 ( .A1(n534), .A2(n551), .ZN(n535) );
  NOR2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n572), .A2(n547), .ZN(n537) );
  XNOR2_X1 U603 ( .A(KEYINPUT114), .B(n537), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U606 ( .A1(n547), .A2(n539), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U608 ( .A(G120GAT), .B(n542), .Z(G1341GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n545) );
  NAND2_X1 U610 ( .A1(n547), .A2(n543), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U612 ( .A(G127GAT), .B(n546), .Z(G1342GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U614 ( .A1(n547), .A2(n562), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U616 ( .A(G134GAT), .B(n550), .Z(G1343GAT) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n556) );
  NOR2_X1 U618 ( .A1(n553), .A2(n556), .ZN(n554) );
  XOR2_X1 U619 ( .A(G141GAT), .B(n554), .Z(n555) );
  XNOR2_X1 U620 ( .A(KEYINPUT118), .B(n555), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n559) );
  INV_X1 U622 ( .A(n556), .ZN(n563) );
  NAND2_X1 U623 ( .A1(n563), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  NAND2_X1 U626 ( .A1(n563), .A2(n580), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n572), .A2(n565), .ZN(n566) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(n566), .ZN(G1348GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U635 ( .A(KEYINPUT59), .B(n569), .Z(n574) );
  NOR2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n583) );
  NAND2_X1 U637 ( .A1(n583), .A2(n572), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  INV_X1 U639 ( .A(n583), .ZN(n575) );
  NOR2_X1 U640 ( .A1(n575), .A2(n369), .ZN(n579) );
  XOR2_X1 U641 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n577) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n583), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n585) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

