

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U557 ( .A1(n785), .A2(n784), .ZN(n811) );
  AND2_X1 U558 ( .A1(n792), .A2(n818), .ZN(n525) );
  NOR2_X2 U559 ( .A1(G2105), .A2(G2104), .ZN(n539) );
  NOR2_X1 U560 ( .A1(G651), .A2(n648), .ZN(n657) );
  NOR2_X1 U561 ( .A1(n547), .A2(n546), .ZN(G164) );
  NOR2_X1 U562 ( .A1(G651), .A2(G543), .ZN(n652) );
  NAND2_X1 U563 ( .A1(n652), .A2(G89), .ZN(n526) );
  XNOR2_X1 U564 ( .A(n526), .B(KEYINPUT4), .ZN(n528) );
  XOR2_X1 U565 ( .A(G543), .B(KEYINPUT0), .Z(n648) );
  INV_X1 U566 ( .A(G651), .ZN(n530) );
  NOR2_X1 U567 ( .A1(n648), .A2(n530), .ZN(n653) );
  NAND2_X1 U568 ( .A1(G76), .A2(n653), .ZN(n527) );
  NAND2_X1 U569 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U570 ( .A(n529), .B(KEYINPUT5), .ZN(n536) );
  NAND2_X1 U571 ( .A1(G51), .A2(n657), .ZN(n533) );
  NOR2_X1 U572 ( .A1(G543), .A2(n530), .ZN(n531) );
  XOR2_X1 U573 ( .A(KEYINPUT1), .B(n531), .Z(n658) );
  NAND2_X1 U574 ( .A1(G63), .A2(n658), .ZN(n532) );
  NAND2_X1 U575 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U576 ( .A(KEYINPUT6), .B(n534), .Z(n535) );
  NAND2_X1 U577 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U578 ( .A(n537), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U579 ( .A(G168), .B(KEYINPUT8), .Z(n538) );
  XNOR2_X1 U580 ( .A(KEYINPUT74), .B(n538), .ZN(G286) );
  XOR2_X2 U581 ( .A(KEYINPUT17), .B(n539), .Z(n884) );
  NAND2_X1 U582 ( .A1(n884), .A2(G138), .ZN(n540) );
  XNOR2_X1 U583 ( .A(KEYINPUT85), .B(n540), .ZN(n547) );
  AND2_X1 U584 ( .A1(G2105), .A2(G2104), .ZN(n888) );
  NAND2_X1 U585 ( .A1(n888), .A2(G114), .ZN(n545) );
  INV_X1 U586 ( .A(G2105), .ZN(n541) );
  AND2_X1 U587 ( .A1(n541), .A2(G2104), .ZN(n885) );
  NAND2_X1 U588 ( .A1(G102), .A2(n885), .ZN(n543) );
  NOR2_X1 U589 ( .A1(G2104), .A2(n541), .ZN(n889) );
  NAND2_X1 U590 ( .A1(G126), .A2(n889), .ZN(n542) );
  AND2_X1 U591 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U592 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U593 ( .A1(G101), .A2(n885), .ZN(n548) );
  XOR2_X1 U594 ( .A(KEYINPUT23), .B(n548), .Z(n551) );
  NAND2_X1 U595 ( .A1(G137), .A2(n884), .ZN(n549) );
  XOR2_X1 U596 ( .A(n549), .B(KEYINPUT65), .Z(n550) );
  NAND2_X1 U597 ( .A1(n551), .A2(n550), .ZN(n555) );
  NAND2_X1 U598 ( .A1(G113), .A2(n888), .ZN(n553) );
  NAND2_X1 U599 ( .A1(G125), .A2(n889), .ZN(n552) );
  NAND2_X1 U600 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X2 U601 ( .A1(n555), .A2(n554), .ZN(G160) );
  XOR2_X1 U602 ( .A(G2435), .B(G2454), .Z(n557) );
  XNOR2_X1 U603 ( .A(KEYINPUT105), .B(G2438), .ZN(n556) );
  XNOR2_X1 U604 ( .A(n557), .B(n556), .ZN(n564) );
  XOR2_X1 U605 ( .A(G2446), .B(G2430), .Z(n559) );
  XNOR2_X1 U606 ( .A(G2451), .B(G2443), .ZN(n558) );
  XNOR2_X1 U607 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U608 ( .A(n560), .B(G2427), .Z(n562) );
  XNOR2_X1 U609 ( .A(G1341), .B(G1348), .ZN(n561) );
  XNOR2_X1 U610 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U611 ( .A(n564), .B(n563), .ZN(n565) );
  AND2_X1 U612 ( .A1(n565), .A2(G14), .ZN(G401) );
  AND2_X1 U613 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U614 ( .A(G57), .ZN(G237) );
  NAND2_X1 U615 ( .A1(G52), .A2(n657), .ZN(n567) );
  NAND2_X1 U616 ( .A1(G64), .A2(n658), .ZN(n566) );
  NAND2_X1 U617 ( .A1(n567), .A2(n566), .ZN(n572) );
  NAND2_X1 U618 ( .A1(G90), .A2(n652), .ZN(n569) );
  NAND2_X1 U619 ( .A1(G77), .A2(n653), .ZN(n568) );
  NAND2_X1 U620 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U621 ( .A(KEYINPUT9), .B(n570), .Z(n571) );
  NOR2_X1 U622 ( .A1(n572), .A2(n571), .ZN(G171) );
  NAND2_X1 U623 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U624 ( .A(n573), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U625 ( .A(G223), .ZN(n833) );
  NAND2_X1 U626 ( .A1(n833), .A2(G567), .ZN(n574) );
  XOR2_X1 U627 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  XOR2_X1 U628 ( .A(KEYINPUT14), .B(KEYINPUT71), .Z(n576) );
  NAND2_X1 U629 ( .A1(G56), .A2(n658), .ZN(n575) );
  XNOR2_X1 U630 ( .A(n576), .B(n575), .ZN(n586) );
  NAND2_X1 U631 ( .A1(G43), .A2(n657), .ZN(n577) );
  XNOR2_X1 U632 ( .A(n577), .B(KEYINPUT73), .ZN(n584) );
  NAND2_X1 U633 ( .A1(G81), .A2(n652), .ZN(n578) );
  XNOR2_X1 U634 ( .A(n578), .B(KEYINPUT72), .ZN(n579) );
  XNOR2_X1 U635 ( .A(n579), .B(KEYINPUT12), .ZN(n581) );
  NAND2_X1 U636 ( .A1(G68), .A2(n653), .ZN(n580) );
  NAND2_X1 U637 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U638 ( .A(KEYINPUT13), .B(n582), .Z(n583) );
  NOR2_X1 U639 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U640 ( .A1(n586), .A2(n585), .ZN(n971) );
  INV_X1 U641 ( .A(G860), .ZN(n840) );
  OR2_X1 U642 ( .A1(n971), .A2(n840), .ZN(G153) );
  INV_X1 U643 ( .A(G171), .ZN(G301) );
  NAND2_X1 U644 ( .A1(G868), .A2(G301), .ZN(n595) );
  NAND2_X1 U645 ( .A1(G54), .A2(n657), .ZN(n588) );
  NAND2_X1 U646 ( .A1(G66), .A2(n658), .ZN(n587) );
  NAND2_X1 U647 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U648 ( .A1(G92), .A2(n652), .ZN(n590) );
  NAND2_X1 U649 ( .A1(G79), .A2(n653), .ZN(n589) );
  NAND2_X1 U650 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U651 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U652 ( .A(KEYINPUT15), .B(n593), .Z(n911) );
  INV_X1 U653 ( .A(n911), .ZN(n972) );
  INV_X1 U654 ( .A(G868), .ZN(n671) );
  NAND2_X1 U655 ( .A1(n972), .A2(n671), .ZN(n594) );
  NAND2_X1 U656 ( .A1(n595), .A2(n594), .ZN(G284) );
  NAND2_X1 U657 ( .A1(G53), .A2(n657), .ZN(n597) );
  NAND2_X1 U658 ( .A1(G65), .A2(n658), .ZN(n596) );
  NAND2_X1 U659 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U660 ( .A1(G91), .A2(n652), .ZN(n599) );
  NAND2_X1 U661 ( .A1(G78), .A2(n653), .ZN(n598) );
  NAND2_X1 U662 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U663 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U664 ( .A(KEYINPUT70), .B(n602), .Z(G299) );
  NAND2_X1 U665 ( .A1(G868), .A2(G286), .ZN(n604) );
  NAND2_X1 U666 ( .A1(G299), .A2(n671), .ZN(n603) );
  NAND2_X1 U667 ( .A1(n604), .A2(n603), .ZN(G297) );
  NAND2_X1 U668 ( .A1(G559), .A2(n840), .ZN(n605) );
  XOR2_X1 U669 ( .A(KEYINPUT75), .B(n605), .Z(n606) );
  NAND2_X1 U670 ( .A1(n606), .A2(n911), .ZN(n607) );
  XNOR2_X1 U671 ( .A(n607), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U672 ( .A1(G868), .A2(n971), .ZN(n610) );
  NAND2_X1 U673 ( .A1(G868), .A2(n911), .ZN(n608) );
  NOR2_X1 U674 ( .A1(G559), .A2(n608), .ZN(n609) );
  NOR2_X1 U675 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U676 ( .A1(G123), .A2(n889), .ZN(n611) );
  XNOR2_X1 U677 ( .A(n611), .B(KEYINPUT18), .ZN(n613) );
  NAND2_X1 U678 ( .A1(n888), .A2(G111), .ZN(n612) );
  NAND2_X1 U679 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U680 ( .A1(G135), .A2(n884), .ZN(n615) );
  NAND2_X1 U681 ( .A1(G99), .A2(n885), .ZN(n614) );
  NAND2_X1 U682 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U683 ( .A1(n617), .A2(n616), .ZN(n928) );
  XNOR2_X1 U684 ( .A(n928), .B(G2096), .ZN(n619) );
  INV_X1 U685 ( .A(G2100), .ZN(n618) );
  NAND2_X1 U686 ( .A1(n619), .A2(n618), .ZN(G156) );
  NAND2_X1 U687 ( .A1(n652), .A2(G85), .ZN(n620) );
  XNOR2_X1 U688 ( .A(n620), .B(KEYINPUT66), .ZN(n622) );
  NAND2_X1 U689 ( .A1(G72), .A2(n653), .ZN(n621) );
  NAND2_X1 U690 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U691 ( .A(n623), .B(KEYINPUT67), .ZN(n625) );
  NAND2_X1 U692 ( .A1(G60), .A2(n658), .ZN(n624) );
  NAND2_X1 U693 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U694 ( .A1(G47), .A2(n657), .ZN(n626) );
  XOR2_X1 U695 ( .A(KEYINPUT68), .B(n626), .Z(n627) );
  NOR2_X1 U696 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U697 ( .A(KEYINPUT69), .B(n629), .ZN(G290) );
  NAND2_X1 U698 ( .A1(G86), .A2(n652), .ZN(n631) );
  NAND2_X1 U699 ( .A1(G61), .A2(n658), .ZN(n630) );
  NAND2_X1 U700 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U701 ( .A(KEYINPUT78), .B(n632), .ZN(n636) );
  NAND2_X1 U702 ( .A1(G73), .A2(n653), .ZN(n633) );
  XNOR2_X1 U703 ( .A(n633), .B(KEYINPUT2), .ZN(n634) );
  XNOR2_X1 U704 ( .A(n634), .B(KEYINPUT79), .ZN(n635) );
  NOR2_X1 U705 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U706 ( .A1(n657), .A2(G48), .ZN(n637) );
  NAND2_X1 U707 ( .A1(n638), .A2(n637), .ZN(G305) );
  NAND2_X1 U708 ( .A1(G88), .A2(n652), .ZN(n640) );
  NAND2_X1 U709 ( .A1(G75), .A2(n653), .ZN(n639) );
  NAND2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U711 ( .A1(G50), .A2(n657), .ZN(n642) );
  NAND2_X1 U712 ( .A1(G62), .A2(n658), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U714 ( .A1(n644), .A2(n643), .ZN(G166) );
  NAND2_X1 U715 ( .A1(G49), .A2(n657), .ZN(n646) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n645) );
  NAND2_X1 U717 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U718 ( .A1(n658), .A2(n647), .ZN(n650) );
  NAND2_X1 U719 ( .A1(n648), .A2(G87), .ZN(n649) );
  NAND2_X1 U720 ( .A1(n650), .A2(n649), .ZN(G288) );
  NAND2_X1 U721 ( .A1(G559), .A2(n911), .ZN(n651) );
  XOR2_X1 U722 ( .A(n971), .B(n651), .Z(n839) );
  NAND2_X1 U723 ( .A1(G93), .A2(n652), .ZN(n655) );
  NAND2_X1 U724 ( .A1(G80), .A2(n653), .ZN(n654) );
  NAND2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U726 ( .A(KEYINPUT76), .B(n656), .ZN(n662) );
  NAND2_X1 U727 ( .A1(G55), .A2(n657), .ZN(n660) );
  NAND2_X1 U728 ( .A1(G67), .A2(n658), .ZN(n659) );
  NAND2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U730 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U731 ( .A(KEYINPUT77), .B(n663), .ZN(n841) );
  XOR2_X1 U732 ( .A(n841), .B(G290), .Z(n669) );
  XNOR2_X1 U733 ( .A(KEYINPUT19), .B(KEYINPUT80), .ZN(n665) );
  XNOR2_X1 U734 ( .A(G305), .B(G166), .ZN(n664) );
  XNOR2_X1 U735 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U736 ( .A(G299), .B(n666), .ZN(n667) );
  XNOR2_X1 U737 ( .A(n667), .B(G288), .ZN(n668) );
  XNOR2_X1 U738 ( .A(n669), .B(n668), .ZN(n910) );
  XNOR2_X1 U739 ( .A(n839), .B(n910), .ZN(n670) );
  NAND2_X1 U740 ( .A1(n670), .A2(G868), .ZN(n673) );
  NAND2_X1 U741 ( .A1(n671), .A2(n841), .ZN(n672) );
  NAND2_X1 U742 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U743 ( .A1(G2078), .A2(G2084), .ZN(n674) );
  XOR2_X1 U744 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U745 ( .A1(G2090), .A2(n675), .ZN(n676) );
  XNOR2_X1 U746 ( .A(KEYINPUT21), .B(n676), .ZN(n677) );
  NAND2_X1 U747 ( .A1(n677), .A2(G2072), .ZN(n678) );
  XOR2_X1 U748 ( .A(KEYINPUT81), .B(n678), .Z(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U750 ( .A1(G132), .A2(G82), .ZN(n679) );
  XNOR2_X1 U751 ( .A(n679), .B(KEYINPUT22), .ZN(n680) );
  XNOR2_X1 U752 ( .A(n680), .B(KEYINPUT82), .ZN(n681) );
  NOR2_X1 U753 ( .A1(G218), .A2(n681), .ZN(n682) );
  XOR2_X1 U754 ( .A(KEYINPUT83), .B(n682), .Z(n683) );
  NAND2_X1 U755 ( .A1(G96), .A2(n683), .ZN(n837) );
  NAND2_X1 U756 ( .A1(G2106), .A2(n837), .ZN(n684) );
  XNOR2_X1 U757 ( .A(KEYINPUT84), .B(n684), .ZN(n688) );
  NAND2_X1 U758 ( .A1(G69), .A2(G120), .ZN(n685) );
  NOR2_X1 U759 ( .A1(G237), .A2(n685), .ZN(n686) );
  NAND2_X1 U760 ( .A1(G108), .A2(n686), .ZN(n838) );
  NAND2_X1 U761 ( .A1(G567), .A2(n838), .ZN(n687) );
  NAND2_X1 U762 ( .A1(n688), .A2(n687), .ZN(n843) );
  NAND2_X1 U763 ( .A1(G483), .A2(G661), .ZN(n689) );
  NOR2_X1 U764 ( .A1(n843), .A2(n689), .ZN(n836) );
  NAND2_X1 U765 ( .A1(n836), .A2(G36), .ZN(G176) );
  XOR2_X1 U766 ( .A(KEYINPUT86), .B(G166), .Z(G303) );
  NOR2_X1 U767 ( .A1(G164), .A2(G1384), .ZN(n721) );
  NAND2_X1 U768 ( .A1(G160), .A2(G40), .ZN(n690) );
  NOR2_X1 U769 ( .A1(n721), .A2(n690), .ZN(n805) );
  XNOR2_X1 U770 ( .A(G2067), .B(KEYINPUT37), .ZN(n803) );
  NAND2_X1 U771 ( .A1(G140), .A2(n884), .ZN(n692) );
  NAND2_X1 U772 ( .A1(G104), .A2(n885), .ZN(n691) );
  NAND2_X1 U773 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U774 ( .A(KEYINPUT34), .B(n693), .ZN(n699) );
  NAND2_X1 U775 ( .A1(n889), .A2(G128), .ZN(n694) );
  XOR2_X1 U776 ( .A(KEYINPUT87), .B(n694), .Z(n696) );
  NAND2_X1 U777 ( .A1(n888), .A2(G116), .ZN(n695) );
  NAND2_X1 U778 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U779 ( .A(KEYINPUT35), .B(n697), .Z(n698) );
  NOR2_X1 U780 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U781 ( .A(KEYINPUT36), .B(n700), .ZN(n907) );
  NOR2_X1 U782 ( .A1(n803), .A2(n907), .ZN(n926) );
  NAND2_X1 U783 ( .A1(n805), .A2(n926), .ZN(n801) );
  NAND2_X1 U784 ( .A1(G105), .A2(n885), .ZN(n701) );
  XNOR2_X1 U785 ( .A(n701), .B(KEYINPUT38), .ZN(n708) );
  NAND2_X1 U786 ( .A1(G141), .A2(n884), .ZN(n703) );
  NAND2_X1 U787 ( .A1(G129), .A2(n889), .ZN(n702) );
  NAND2_X1 U788 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U789 ( .A1(n888), .A2(G117), .ZN(n704) );
  XOR2_X1 U790 ( .A(KEYINPUT90), .B(n704), .Z(n705) );
  NOR2_X1 U791 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U792 ( .A1(n708), .A2(n707), .ZN(n901) );
  NAND2_X1 U793 ( .A1(G1996), .A2(n901), .ZN(n709) );
  XNOR2_X1 U794 ( .A(n709), .B(KEYINPUT91), .ZN(n718) );
  XNOR2_X1 U795 ( .A(KEYINPUT89), .B(G1991), .ZN(n946) );
  NAND2_X1 U796 ( .A1(G131), .A2(n884), .ZN(n711) );
  NAND2_X1 U797 ( .A1(G95), .A2(n885), .ZN(n710) );
  NAND2_X1 U798 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U799 ( .A(KEYINPUT88), .B(n712), .ZN(n716) );
  NAND2_X1 U800 ( .A1(G107), .A2(n888), .ZN(n714) );
  NAND2_X1 U801 ( .A1(G119), .A2(n889), .ZN(n713) );
  NAND2_X1 U802 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U803 ( .A1(n716), .A2(n715), .ZN(n900) );
  NOR2_X1 U804 ( .A1(n946), .A2(n900), .ZN(n717) );
  NOR2_X1 U805 ( .A1(n718), .A2(n717), .ZN(n930) );
  INV_X1 U806 ( .A(n805), .ZN(n719) );
  NOR2_X1 U807 ( .A1(n930), .A2(n719), .ZN(n798) );
  INV_X1 U808 ( .A(n798), .ZN(n720) );
  NAND2_X1 U809 ( .A1(n801), .A2(n720), .ZN(n824) );
  AND2_X1 U810 ( .A1(G160), .A2(G40), .ZN(n722) );
  NAND2_X2 U811 ( .A1(n722), .A2(n721), .ZN(n767) );
  NAND2_X1 U812 ( .A1(n767), .A2(G8), .ZN(n723) );
  XNOR2_X2 U813 ( .A(n723), .B(KEYINPUT92), .ZN(n789) );
  NOR2_X1 U814 ( .A1(n789), .A2(G1966), .ZN(n779) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n767), .ZN(n780) );
  NOR2_X1 U816 ( .A1(n779), .A2(n780), .ZN(n724) );
  NAND2_X1 U817 ( .A1(n724), .A2(G8), .ZN(n726) );
  XNOR2_X1 U818 ( .A(KEYINPUT96), .B(KEYINPUT30), .ZN(n725) );
  XNOR2_X1 U819 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U820 ( .A1(G168), .A2(n727), .ZN(n728) );
  XNOR2_X1 U821 ( .A(n728), .B(KEYINPUT97), .ZN(n732) );
  XOR2_X1 U822 ( .A(G2078), .B(KEYINPUT25), .Z(n947) );
  NOR2_X1 U823 ( .A1(n947), .A2(n767), .ZN(n730) );
  INV_X1 U824 ( .A(n767), .ZN(n746) );
  NOR2_X1 U825 ( .A1(n746), .A2(G1961), .ZN(n729) );
  NOR2_X1 U826 ( .A1(n730), .A2(n729), .ZN(n762) );
  NAND2_X1 U827 ( .A1(n762), .A2(G301), .ZN(n731) );
  NAND2_X1 U828 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U829 ( .A(n733), .B(KEYINPUT31), .ZN(n777) );
  INV_X1 U830 ( .A(n767), .ZN(n734) );
  NAND2_X1 U831 ( .A1(G2072), .A2(n734), .ZN(n735) );
  XOR2_X1 U832 ( .A(n735), .B(KEYINPUT27), .Z(n736) );
  XNOR2_X1 U833 ( .A(KEYINPUT93), .B(n736), .ZN(n738) );
  INV_X1 U834 ( .A(G1956), .ZN(n1001) );
  NOR2_X1 U835 ( .A1(n746), .A2(n1001), .ZN(n737) );
  NOR2_X1 U836 ( .A1(n738), .A2(n737), .ZN(n742) );
  INV_X1 U837 ( .A(G299), .ZN(n741) );
  NOR2_X1 U838 ( .A1(n742), .A2(n741), .ZN(n740) );
  XOR2_X1 U839 ( .A(KEYINPUT28), .B(KEYINPUT94), .Z(n739) );
  XNOR2_X1 U840 ( .A(n740), .B(n739), .ZN(n760) );
  NAND2_X1 U841 ( .A1(n742), .A2(n741), .ZN(n758) );
  NAND2_X1 U842 ( .A1(G1348), .A2(n767), .ZN(n744) );
  NAND2_X1 U843 ( .A1(G2067), .A2(n746), .ZN(n743) );
  NAND2_X1 U844 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U845 ( .A(KEYINPUT95), .B(n745), .ZN(n754) );
  OR2_X1 U846 ( .A1(n911), .A2(n754), .ZN(n753) );
  AND2_X1 U847 ( .A1(n746), .A2(G1996), .ZN(n748) );
  XOR2_X1 U848 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n747) );
  XNOR2_X1 U849 ( .A(n748), .B(n747), .ZN(n750) );
  NAND2_X1 U850 ( .A1(n767), .A2(G1341), .ZN(n749) );
  NAND2_X1 U851 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U852 ( .A1(n971), .A2(n751), .ZN(n752) );
  NAND2_X1 U853 ( .A1(n753), .A2(n752), .ZN(n756) );
  NAND2_X1 U854 ( .A1(n754), .A2(n911), .ZN(n755) );
  AND2_X1 U855 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U856 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U857 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U858 ( .A(n761), .B(KEYINPUT29), .Z(n764) );
  OR2_X1 U859 ( .A1(G301), .A2(n762), .ZN(n763) );
  NAND2_X1 U860 ( .A1(n764), .A2(n763), .ZN(n776) );
  NAND2_X1 U861 ( .A1(n777), .A2(n776), .ZN(n765) );
  NAND2_X1 U862 ( .A1(n765), .A2(G286), .ZN(n766) );
  XNOR2_X1 U863 ( .A(n766), .B(KEYINPUT99), .ZN(n773) );
  NOR2_X1 U864 ( .A1(n789), .A2(G1971), .ZN(n769) );
  NOR2_X1 U865 ( .A1(G2090), .A2(n767), .ZN(n768) );
  NOR2_X1 U866 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U867 ( .A1(G303), .A2(n770), .ZN(n771) );
  XOR2_X1 U868 ( .A(KEYINPUT100), .B(n771), .Z(n772) );
  OR2_X1 U869 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U870 ( .A1(n774), .A2(G8), .ZN(n775) );
  XNOR2_X1 U871 ( .A(KEYINPUT32), .B(n775), .ZN(n785) );
  AND2_X1 U872 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U873 ( .A1(n779), .A2(n778), .ZN(n782) );
  NAND2_X1 U874 ( .A1(G8), .A2(n780), .ZN(n781) );
  NAND2_X1 U875 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U876 ( .A(KEYINPUT98), .B(n783), .ZN(n784) );
  NOR2_X1 U877 ( .A1(G303), .A2(G2090), .ZN(n786) );
  NAND2_X1 U878 ( .A1(G8), .A2(n786), .ZN(n787) );
  XOR2_X1 U879 ( .A(KEYINPUT104), .B(n787), .Z(n788) );
  NOR2_X1 U880 ( .A1(n811), .A2(n788), .ZN(n790) );
  INV_X1 U881 ( .A(n789), .ZN(n818) );
  NOR2_X1 U882 ( .A1(n790), .A2(n818), .ZN(n793) );
  NOR2_X1 U883 ( .A1(G1981), .A2(G305), .ZN(n791) );
  XNOR2_X1 U884 ( .A(KEYINPUT24), .B(n791), .ZN(n792) );
  OR2_X1 U885 ( .A1(n793), .A2(n525), .ZN(n794) );
  XNOR2_X1 U886 ( .A(G1986), .B(G290), .ZN(n985) );
  NAND2_X1 U887 ( .A1(n985), .A2(n805), .ZN(n826) );
  NAND2_X1 U888 ( .A1(n794), .A2(n826), .ZN(n795) );
  NOR2_X1 U889 ( .A1(n824), .A2(n795), .ZN(n808) );
  NOR2_X1 U890 ( .A1(G1996), .A2(n901), .ZN(n922) );
  AND2_X1 U891 ( .A1(n946), .A2(n900), .ZN(n932) );
  NOR2_X1 U892 ( .A1(G1986), .A2(G290), .ZN(n796) );
  NOR2_X1 U893 ( .A1(n932), .A2(n796), .ZN(n797) );
  NOR2_X1 U894 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U895 ( .A1(n922), .A2(n799), .ZN(n800) );
  XNOR2_X1 U896 ( .A(KEYINPUT39), .B(n800), .ZN(n802) );
  NAND2_X1 U897 ( .A1(n802), .A2(n801), .ZN(n804) );
  NAND2_X1 U898 ( .A1(n803), .A2(n907), .ZN(n939) );
  NAND2_X1 U899 ( .A1(n804), .A2(n939), .ZN(n806) );
  AND2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U901 ( .A1(n808), .A2(n807), .ZN(n831) );
  NOR2_X1 U902 ( .A1(G303), .A2(G1971), .ZN(n809) );
  XNOR2_X1 U903 ( .A(n809), .B(KEYINPUT101), .ZN(n810) );
  NOR2_X1 U904 ( .A1(G1976), .A2(G288), .ZN(n819) );
  INV_X1 U905 ( .A(n819), .ZN(n982) );
  NAND2_X1 U906 ( .A1(n810), .A2(n982), .ZN(n812) );
  OR2_X2 U907 ( .A1(n812), .A2(n811), .ZN(n817) );
  INV_X1 U908 ( .A(KEYINPUT33), .ZN(n814) );
  NAND2_X1 U909 ( .A1(G288), .A2(G1976), .ZN(n813) );
  XNOR2_X1 U910 ( .A(n813), .B(KEYINPUT102), .ZN(n983) );
  AND2_X1 U911 ( .A1(n814), .A2(n983), .ZN(n815) );
  AND2_X1 U912 ( .A1(n815), .A2(n818), .ZN(n816) );
  NAND2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n822) );
  NAND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n820), .A2(KEYINPUT33), .ZN(n821) );
  NAND2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U917 ( .A(KEYINPUT103), .B(n823), .Z(n829) );
  XOR2_X1 U918 ( .A(G1981), .B(G305), .Z(n978) );
  INV_X1 U919 ( .A(n824), .ZN(n825) );
  AND2_X1 U920 ( .A1(n978), .A2(n825), .ZN(n827) );
  AND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U923 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U924 ( .A(n832), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U927 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U929 ( .A1(n836), .A2(n835), .ZN(G188) );
  INV_X1 U931 ( .A(G132), .ZN(G219) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(G82), .ZN(G220) );
  INV_X1 U935 ( .A(G69), .ZN(G235) );
  NOR2_X1 U936 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  NAND2_X1 U938 ( .A1(n840), .A2(n839), .ZN(n842) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(G145) );
  INV_X1 U940 ( .A(n843), .ZN(G319) );
  XOR2_X1 U941 ( .A(KEYINPUT109), .B(G1961), .Z(n845) );
  XNOR2_X1 U942 ( .A(G1981), .B(G1966), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U944 ( .A(n846), .B(KEYINPUT41), .Z(n848) );
  XNOR2_X1 U945 ( .A(G1996), .B(G1991), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U947 ( .A(G1976), .B(G1971), .Z(n850) );
  XNOR2_X1 U948 ( .A(G1986), .B(G1956), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U950 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U951 ( .A(KEYINPUT108), .B(G2474), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(G229) );
  XOR2_X1 U953 ( .A(KEYINPUT43), .B(KEYINPUT42), .Z(n856) );
  XNOR2_X1 U954 ( .A(G2678), .B(KEYINPUT107), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U956 ( .A(KEYINPUT106), .B(G2090), .Z(n858) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2072), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U959 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U960 ( .A(G2096), .B(G2100), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n864) );
  XOR2_X1 U962 ( .A(G2078), .B(G2084), .Z(n863) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(G227) );
  NAND2_X1 U964 ( .A1(G124), .A2(n889), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n865), .B(KEYINPUT110), .ZN(n866) );
  XNOR2_X1 U966 ( .A(KEYINPUT44), .B(n866), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G112), .A2(n888), .ZN(n867) );
  XOR2_X1 U968 ( .A(KEYINPUT111), .B(n867), .Z(n868) );
  NAND2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n873) );
  NAND2_X1 U970 ( .A1(G136), .A2(n884), .ZN(n871) );
  NAND2_X1 U971 ( .A1(G100), .A2(n885), .ZN(n870) );
  NAND2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U973 ( .A1(n873), .A2(n872), .ZN(G162) );
  NAND2_X1 U974 ( .A1(n885), .A2(G106), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n874), .B(KEYINPUT114), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G142), .A2(n884), .ZN(n875) );
  NAND2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n877), .B(KEYINPUT45), .ZN(n883) );
  NAND2_X1 U979 ( .A1(G118), .A2(n888), .ZN(n878) );
  XNOR2_X1 U980 ( .A(n878), .B(KEYINPUT113), .ZN(n881) );
  NAND2_X1 U981 ( .A1(G130), .A2(n889), .ZN(n879) );
  XOR2_X1 U982 ( .A(KEYINPUT112), .B(n879), .Z(n880) );
  NOR2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n882) );
  NAND2_X1 U984 ( .A1(n883), .A2(n882), .ZN(n895) );
  NAND2_X1 U985 ( .A1(G139), .A2(n884), .ZN(n887) );
  NAND2_X1 U986 ( .A1(G103), .A2(n885), .ZN(n886) );
  NAND2_X1 U987 ( .A1(n887), .A2(n886), .ZN(n894) );
  NAND2_X1 U988 ( .A1(G115), .A2(n888), .ZN(n891) );
  NAND2_X1 U989 ( .A1(G127), .A2(n889), .ZN(n890) );
  NAND2_X1 U990 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U991 ( .A(KEYINPUT47), .B(n892), .Z(n893) );
  NOR2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n935) );
  XNOR2_X1 U993 ( .A(n895), .B(n935), .ZN(n896) );
  XNOR2_X1 U994 ( .A(G164), .B(n896), .ZN(n905) );
  XOR2_X1 U995 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n898) );
  XNOR2_X1 U996 ( .A(G160), .B(G162), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n928), .B(n899), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1002 ( .A(n907), .B(n906), .Z(n908) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n908), .ZN(n909) );
  XOR2_X1 U1004 ( .A(KEYINPUT115), .B(n909), .Z(G395) );
  XNOR2_X1 U1005 ( .A(G286), .B(n910), .ZN(n913) );
  XNOR2_X1 U1006 ( .A(G171), .B(n911), .ZN(n912) );
  XNOR2_X1 U1007 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1008 ( .A(n914), .B(n971), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n915), .ZN(G397) );
  NOR2_X1 U1010 ( .A1(G229), .A2(G227), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(G401), .A2(n917), .ZN(n918) );
  AND2_X1 U1013 ( .A1(G319), .A2(n918), .ZN(n920) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1015 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1018 ( .A(G2090), .B(G162), .Z(n921) );
  NOR2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1020 ( .A(KEYINPUT116), .B(n923), .Z(n924) );
  XOR2_X1 U1021 ( .A(KEYINPUT51), .B(n924), .Z(n925) );
  NOR2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n934) );
  XOR2_X1 U1023 ( .A(G2084), .B(G160), .Z(n927) );
  NOR2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1026 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1027 ( .A1(n934), .A2(n933), .ZN(n942) );
  XOR2_X1 U1028 ( .A(G2072), .B(n935), .Z(n937) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n936) );
  NOR2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1031 ( .A(n938), .B(KEYINPUT50), .ZN(n940) );
  NAND2_X1 U1032 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1033 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1034 ( .A(KEYINPUT52), .B(n943), .ZN(n944) );
  INV_X1 U1035 ( .A(KEYINPUT55), .ZN(n967) );
  NAND2_X1 U1036 ( .A1(n944), .A2(n967), .ZN(n945) );
  NAND2_X1 U1037 ( .A1(n945), .A2(G29), .ZN(n1029) );
  XOR2_X1 U1038 ( .A(n946), .B(G25), .Z(n949) );
  XNOR2_X1 U1039 ( .A(G27), .B(n947), .ZN(n948) );
  NOR2_X1 U1040 ( .A1(n949), .A2(n948), .ZN(n957) );
  XNOR2_X1 U1041 ( .A(G2067), .B(G26), .ZN(n951) );
  XNOR2_X1 U1042 ( .A(G33), .B(G2072), .ZN(n950) );
  NOR2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1044 ( .A1(G28), .A2(n952), .ZN(n955) );
  XOR2_X1 U1045 ( .A(G32), .B(G1996), .Z(n953) );
  XNOR2_X1 U1046 ( .A(KEYINPUT117), .B(n953), .ZN(n954) );
  NOR2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1048 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(n958), .B(KEYINPUT53), .ZN(n959) );
  XNOR2_X1 U1050 ( .A(KEYINPUT118), .B(n959), .ZN(n965) );
  XOR2_X1 U1051 ( .A(KEYINPUT119), .B(G34), .Z(n961) );
  XNOR2_X1 U1052 ( .A(G2084), .B(KEYINPUT54), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(n961), .B(n960), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(G35), .B(G2090), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1057 ( .A(n967), .B(n966), .ZN(n969) );
  INV_X1 U1058 ( .A(G29), .ZN(n968) );
  NAND2_X1 U1059 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1060 ( .A1(G11), .A2(n970), .ZN(n1027) );
  XNOR2_X1 U1061 ( .A(G16), .B(KEYINPUT56), .ZN(n997) );
  XNOR2_X1 U1062 ( .A(n971), .B(G1341), .ZN(n977) );
  XNOR2_X1 U1063 ( .A(G301), .B(G1961), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(n972), .B(G1348), .ZN(n973) );
  NOR2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(KEYINPUT121), .B(n975), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n995) );
  XNOR2_X1 U1068 ( .A(G1966), .B(G168), .ZN(n979) );
  NAND2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(n980), .B(KEYINPUT120), .ZN(n981) );
  XOR2_X1 U1071 ( .A(KEYINPUT57), .B(n981), .Z(n993) );
  XNOR2_X1 U1072 ( .A(G299), .B(n1001), .ZN(n987) );
  NAND2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1075 ( .A1(n987), .A2(n986), .ZN(n990) );
  XNOR2_X1 U1076 ( .A(G1971), .B(G303), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(KEYINPUT122), .B(n988), .ZN(n989) );
  NOR2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(KEYINPUT123), .B(n991), .ZN(n992) );
  NOR2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1082 ( .A1(n997), .A2(n996), .ZN(n1025) );
  INV_X1 U1083 ( .A(G16), .ZN(n1023) );
  XNOR2_X1 U1084 ( .A(G1981), .B(G6), .ZN(n999) );
  XNOR2_X1 U1085 ( .A(G1341), .B(G19), .ZN(n998) );
  NOR2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(KEYINPUT124), .B(n1000), .ZN(n1003) );
  XNOR2_X1 U1088 ( .A(n1001), .B(G20), .ZN(n1002) );
  NAND2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(n1007) );
  XNOR2_X1 U1090 ( .A(KEYINPUT59), .B(KEYINPUT125), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(n1004), .B(G4), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(n1005), .B(G1348), .ZN(n1006) );
  NOR2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1094 ( .A(KEYINPUT60), .B(n1008), .ZN(n1012) );
  XNOR2_X1 U1095 ( .A(G1966), .B(G21), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(G5), .B(G1961), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1020) );
  XNOR2_X1 U1099 ( .A(G1986), .B(G24), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(G23), .B(G1976), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XOR2_X1 U1102 ( .A(G1971), .B(KEYINPUT126), .Z(n1015) );
  XNOR2_X1 U1103 ( .A(G22), .B(n1015), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(KEYINPUT58), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(KEYINPUT61), .B(n1021), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1110 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1111 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1112 ( .A(n1030), .B(KEYINPUT127), .ZN(n1031) );
  XNOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1031), .ZN(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

