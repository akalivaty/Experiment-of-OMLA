//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n211), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n202), .A2(new_n203), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(new_n215), .A2(new_n216), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n213), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n222), .B1(new_n216), .B2(new_n215), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(G20), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT64), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT64), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n257), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(new_n217), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n254), .A2(new_n259), .B1(new_n201), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n259), .B1(new_n210), .B2(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G50), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT9), .ZN(new_n266));
  INV_X1    g0066(.A(G200), .ZN(new_n267));
  OR2_X1    g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  AOI21_X1  g0069(.A(G1698), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n270), .A2(G222), .B1(new_n273), .B2(G77), .ZN(new_n274));
  INV_X1    g0074(.A(G223), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G1698), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(G1), .A2(G13), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n284));
  INV_X1    g0084(.A(G274), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n281), .A2(new_n284), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n286), .B1(new_n288), .B2(G226), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n267), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n283), .A2(G190), .A3(new_n289), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n266), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT10), .B1(new_n290), .B2(KEYINPUT68), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n266), .A2(new_n294), .A3(new_n291), .A4(new_n292), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n283), .A2(new_n289), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G169), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(new_n298), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n296), .A2(new_n297), .B1(new_n265), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT66), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n260), .A2(G77), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  AND3_X1   g0105(.A1(new_n256), .A2(new_n217), .A3(new_n258), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(G1), .B2(new_n211), .ZN(new_n307));
  INV_X1    g0107(.A(G77), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n253), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n310), .A2(new_n248), .B1(G20), .B2(G77), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT15), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n312), .A2(G87), .ZN(new_n313));
  INV_X1    g0113(.A(G87), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(KEYINPUT15), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT65), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(KEYINPUT15), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n312), .A2(G87), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT65), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n316), .A2(new_n251), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n306), .B1(new_n311), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n303), .B1(new_n309), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n304), .B1(new_n263), .B2(G77), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n311), .A2(new_n321), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n324), .B(KEYINPUT66), .C1(new_n325), .C2(new_n306), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n270), .A2(G232), .B1(new_n273), .B2(G107), .ZN(new_n327));
  INV_X1    g0127(.A(G1698), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(new_n268), .B2(new_n269), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G238), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n282), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n286), .B1(new_n288), .B2(G244), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n323), .B(new_n326), .C1(new_n334), .C2(new_n267), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n335), .A2(KEYINPUT67), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(G190), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n335), .B2(KEYINPUT67), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n334), .A2(G179), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n332), .A2(new_n333), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G169), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n340), .A2(new_n342), .B1(new_n323), .B2(new_n326), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n302), .A2(new_n339), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT69), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n310), .A2(new_n261), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(new_n307), .B2(new_n310), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT75), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G58), .A2(G68), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT74), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT74), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(G58), .A3(G68), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n354), .A3(new_n219), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(G20), .B1(G159), .B2(new_n248), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n271), .A2(new_n272), .A3(G20), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT7), .ZN(new_n358));
  OAI21_X1  g0158(.A(G68), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n273), .A2(new_n360), .A3(new_n211), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n356), .B(KEYINPUT16), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n259), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n268), .A2(new_n358), .A3(new_n211), .A4(new_n269), .ZN(new_n364));
  OAI211_X1 g0164(.A(G68), .B(new_n364), .C1(new_n357), .C2(new_n360), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT16), .B1(new_n365), .B2(new_n356), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n350), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n366), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n368), .A2(KEYINPUT75), .A3(new_n259), .A4(new_n362), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n349), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT76), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n281), .A2(new_n371), .A3(G232), .A4(new_n284), .ZN(new_n372));
  INV_X1    g0172(.A(new_n286), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT76), .B1(new_n287), .B2(new_n235), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT77), .ZN(new_n377));
  INV_X1    g0177(.A(G190), .ZN(new_n378));
  OAI211_X1 g0178(.A(G226), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n379));
  OAI211_X1 g0179(.A(G223), .B(new_n328), .C1(new_n271), .C2(new_n272), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n379), .B(new_n380), .C1(new_n250), .C2(new_n314), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n282), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n376), .A2(new_n377), .A3(new_n378), .A4(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n382), .A2(new_n375), .A3(new_n374), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT77), .B1(new_n384), .B2(new_n267), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(G190), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n370), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT17), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n367), .A2(new_n369), .ZN(new_n391));
  INV_X1    g0191(.A(new_n349), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT18), .ZN(new_n394));
  INV_X1    g0194(.A(G169), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n384), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(G179), .B2(new_n384), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n393), .A2(new_n394), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT18), .B1(new_n370), .B2(new_n397), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n370), .A2(KEYINPUT17), .A3(new_n387), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n390), .A2(new_n399), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n347), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n276), .A2(G226), .A3(new_n328), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G97), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n405), .B(new_n406), .C1(new_n277), .C2(new_n235), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n282), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT13), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n286), .B1(new_n288), .B2(G238), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n409), .B1(new_n408), .B2(new_n410), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n267), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n408), .A2(new_n410), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT13), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n416), .A2(new_n378), .A3(new_n411), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n248), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n252), .B2(new_n308), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n259), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT11), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n263), .A2(G68), .ZN(new_n423));
  INV_X1    g0223(.A(G13), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(G1), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(G20), .A3(new_n203), .ZN(new_n426));
  OR3_X1    g0226(.A1(new_n426), .A2(KEYINPUT70), .A3(KEYINPUT12), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT70), .B1(new_n426), .B2(KEYINPUT12), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(KEYINPUT12), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n422), .A2(new_n423), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT71), .B1(new_n418), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT71), .ZN(new_n434));
  AOI211_X1 g0234(.A(new_n434), .B(new_n431), .C1(new_n414), .C2(new_n417), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT14), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n416), .A2(new_n411), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n437), .B1(new_n438), .B2(new_n300), .ZN(new_n439));
  AND2_X1   g0239(.A1(KEYINPUT72), .A2(G169), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n438), .A2(new_n437), .A3(new_n440), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n432), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n436), .B(new_n445), .C1(new_n345), .C2(new_n346), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n404), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(G20), .B1(new_n250), .B2(G97), .ZN(new_n448));
  AND3_X1   g0248(.A1(KEYINPUT79), .A2(G33), .A3(G283), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT79), .B1(G33), .B2(G283), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G116), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G20), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n259), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT20), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n259), .A2(new_n451), .A3(KEYINPUT20), .A4(new_n453), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n210), .A2(G33), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n260), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  AND3_X1   g0261(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n279), .B1(new_n462), .B2(new_n257), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n461), .A2(new_n463), .A3(G116), .A4(new_n256), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n261), .A2(new_n452), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n458), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT21), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT5), .B(G41), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n468), .A2(new_n470), .B1(new_n279), .B2(new_n280), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n210), .A2(G45), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n471), .A2(G270), .B1(G274), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(G264), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n478));
  OAI211_X1 g0278(.A(G257), .B(new_n328), .C1(new_n271), .C2(new_n272), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n268), .A2(G303), .A3(new_n269), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n282), .ZN(new_n482));
  AOI211_X1 g0282(.A(new_n467), .B(new_n395), .C1(new_n477), .C2(new_n482), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n477), .A2(G179), .A3(new_n482), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n466), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n464), .A2(new_n465), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n486), .B1(new_n456), .B2(new_n457), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n477), .A2(new_n482), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(G190), .ZN(new_n489));
  AOI21_X1  g0289(.A(G200), .B1(new_n477), .B2(new_n482), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n488), .A2(G169), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n467), .B1(new_n492), .B2(new_n487), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n485), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(G250), .B(new_n328), .C1(new_n271), .C2(new_n272), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT84), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT84), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n276), .A2(new_n497), .A3(G250), .A4(new_n328), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G294), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n276), .A2(G257), .A3(G1698), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n496), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n282), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n476), .A2(G274), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n471), .A2(G264), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G169), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n501), .A2(new_n282), .B1(G264), .B2(new_n471), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n507), .A2(G179), .A3(new_n503), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n211), .B(G87), .C1(new_n271), .C2(new_n272), .ZN(new_n509));
  NAND2_X1  g0309(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n510), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n276), .A2(new_n211), .A3(G87), .A4(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT23), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(new_n207), .A3(G20), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n211), .A2(G33), .A3(G116), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n511), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT24), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n511), .A2(new_n513), .A3(KEYINPUT24), .A4(new_n518), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n259), .A3(new_n522), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n259), .A2(new_n207), .A3(new_n460), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n425), .A2(G20), .A3(new_n207), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n525), .A2(KEYINPUT25), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n525), .A2(KEYINPUT25), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n506), .A2(new_n508), .B1(new_n523), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n523), .A2(new_n528), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n505), .A2(new_n267), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n507), .A2(new_n378), .A3(new_n503), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n494), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(G244), .B(new_n328), .C1(new_n271), .C2(new_n272), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT4), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT4), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n276), .A2(new_n537), .A3(G244), .A4(new_n328), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n449), .A2(new_n450), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n329), .B2(G250), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n281), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n475), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n470), .B1(new_n543), .B2(new_n473), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n544), .A2(G257), .A3(new_n281), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n503), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n395), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n546), .ZN(new_n548));
  OR2_X1    g0348(.A1(new_n449), .A2(new_n450), .ZN(new_n549));
  OAI211_X1 g0349(.A(G250), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n536), .B2(new_n538), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n548), .B(new_n300), .C1(new_n552), .C2(new_n281), .ZN(new_n553));
  OAI211_X1 g0353(.A(G107), .B(new_n364), .C1(new_n357), .C2(new_n360), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G97), .A2(G107), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(G97), .A2(G107), .ZN(new_n557));
  OAI22_X1  g0357(.A1(new_n556), .A2(new_n557), .B1(KEYINPUT78), .B2(KEYINPUT6), .ZN(new_n558));
  NOR2_X1   g0358(.A1(KEYINPUT78), .A2(KEYINPUT6), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n208), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n558), .A2(new_n560), .A3(G20), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n248), .A2(G77), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n554), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n260), .A2(new_n206), .ZN(new_n565));
  OAI21_X1  g0365(.A(G97), .B1(new_n259), .B2(new_n460), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n564), .A2(new_n259), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n547), .B(new_n553), .C1(new_n567), .C2(KEYINPUT81), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(KEYINPUT81), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(KEYINPUT80), .B1(new_n542), .B2(new_n546), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT80), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n548), .B(new_n572), .C1(new_n552), .C2(new_n281), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n267), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n548), .B1(new_n552), .B2(new_n281), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n567), .B1(new_n575), .B2(new_n378), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n568), .A2(new_n570), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT82), .ZN(new_n578));
  OAI211_X1 g0378(.A(G238), .B(new_n328), .C1(new_n271), .C2(new_n272), .ZN(new_n579));
  OAI211_X1 g0379(.A(G244), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G33), .A2(G116), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n282), .ZN(new_n583));
  OAI21_X1  g0383(.A(G250), .B1(new_n469), .B2(G1), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n210), .A2(G45), .A3(G274), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n281), .ZN(new_n587));
  AOI21_X1  g0387(.A(G169), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n584), .A2(new_n585), .B1(new_n279), .B2(new_n280), .ZN(new_n589));
  AOI211_X1 g0389(.A(G179), .B(new_n589), .C1(new_n582), .C2(new_n282), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n578), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n583), .A2(new_n300), .A3(new_n587), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n589), .B1(new_n582), .B2(new_n282), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n592), .B(KEYINPUT82), .C1(G169), .C2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n211), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n314), .A2(new_n206), .A3(new_n207), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n211), .B(G68), .C1(new_n271), .C2(new_n272), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n211), .A2(G33), .A3(G97), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT19), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n598), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n259), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n306), .A2(new_n320), .A3(new_n316), .A4(new_n461), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n316), .A2(new_n320), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n261), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n591), .A2(new_n594), .A3(new_n608), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n596), .A2(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n610), .A2(new_n599), .B1(new_n256), .B2(new_n463), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n259), .A2(new_n314), .A3(new_n460), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n260), .B1(new_n316), .B2(new_n320), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n593), .A2(G190), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n614), .B(new_n615), .C1(new_n267), .C2(new_n593), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n609), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n577), .A2(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n447), .A2(new_n534), .A3(new_n618), .ZN(G372));
  NAND2_X1  g0419(.A1(new_n296), .A2(new_n297), .ZN(new_n620));
  INV_X1    g0420(.A(new_n401), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT17), .B1(new_n370), .B2(new_n387), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n436), .A2(new_n343), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n624), .B1(new_n625), .B2(new_n445), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n399), .A2(new_n400), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n620), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n301), .A2(new_n265), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT85), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n587), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n589), .A2(KEYINPUT85), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n633), .A2(new_n634), .B1(new_n582), .B2(new_n282), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n608), .B(new_n592), .C1(new_n635), .C2(G169), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT86), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n633), .A2(new_n634), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n583), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n395), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n641), .A2(KEYINPUT86), .A3(new_n592), .A4(new_n608), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n614), .B(new_n615), .C1(new_n635), .C2(new_n267), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n636), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n564), .A2(new_n259), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n566), .A2(new_n565), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(new_n547), .A3(new_n553), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n643), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT81), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n654), .A2(new_n569), .A3(new_n553), .A4(new_n547), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT26), .B1(new_n617), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT87), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n652), .A2(new_n656), .A3(KEYINPUT87), .ZN(new_n660));
  INV_X1    g0460(.A(new_n577), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n506), .A2(new_n508), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n530), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n663), .A2(new_n493), .A3(new_n485), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n533), .A2(new_n645), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n661), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n659), .A2(new_n660), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n447), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n631), .A2(new_n668), .ZN(G369));
  INV_X1    g0469(.A(KEYINPUT88), .ZN(new_n670));
  INV_X1    g0470(.A(new_n425), .ZN(new_n671));
  OR3_X1    g0471(.A1(new_n671), .A2(KEYINPUT27), .A3(G20), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT27), .B1(new_n671), .B2(G20), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(G343), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(new_n487), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n494), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n485), .A2(new_n493), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n678), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n670), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n679), .A2(new_n670), .A3(new_n681), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n529), .A2(new_n677), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n533), .B1(new_n530), .B2(new_n676), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n687), .B1(new_n688), .B2(new_n529), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n680), .A2(new_n677), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n693), .B1(new_n529), .B2(new_n677), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n694), .ZN(G399));
  INV_X1    g0495(.A(new_n214), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT89), .B1(new_n698), .B2(new_n220), .ZN(new_n699));
  NOR4_X1   g0499(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n697), .A2(new_n210), .A3(new_n701), .ZN(new_n702));
  MUX2_X1   g0502(.A(new_n699), .B(KEYINPUT89), .S(new_n702), .Z(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n618), .A2(new_n534), .A3(new_n677), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT31), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n542), .A2(new_n546), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n507), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n484), .A2(new_n593), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n707), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(G179), .B1(new_n477), .B2(new_n482), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n505), .A2(new_n575), .A3(new_n640), .A4(new_n712), .ZN(new_n713));
  AND4_X1   g0513(.A1(G179), .A2(new_n593), .A3(new_n482), .A4(new_n477), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(KEYINPUT30), .A3(new_n507), .A4(new_n708), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n711), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n706), .B1(new_n716), .B2(new_n676), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n705), .A2(new_n717), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n716), .A2(new_n706), .A3(new_n676), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G330), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n661), .A2(KEYINPUT90), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n661), .A2(KEYINPUT90), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n724), .A2(new_n664), .A3(new_n665), .A4(new_n725), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n617), .A2(new_n655), .A3(KEYINPUT26), .ZN(new_n727));
  INV_X1    g0527(.A(new_n643), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(new_n650), .B2(new_n651), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n676), .B1(new_n726), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT29), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n667), .A2(new_n677), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n723), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n704), .B1(new_n736), .B2(G1), .ZN(G364));
  NOR2_X1   g0537(.A1(new_n696), .A2(new_n273), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n738), .A2(G355), .B1(new_n452), .B2(new_n696), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n221), .A2(G45), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n740), .B1(new_n243), .B2(G45), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n214), .A2(new_n273), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n279), .B1(new_n211), .B2(G169), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT92), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G13), .A2(G33), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n743), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n424), .A2(G20), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n210), .B1(new_n752), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n697), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g0555(.A(new_n755), .B(KEYINPUT91), .Z(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n211), .A2(new_n378), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n300), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT93), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT32), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n211), .A2(G190), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G159), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n763), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n766), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(KEYINPUT32), .A3(G159), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n762), .A2(G58), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n300), .A2(new_n267), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n758), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n267), .A2(G179), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n758), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI22_X1  g0577(.A1(G50), .A2(new_n774), .B1(new_n777), .B2(G87), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n775), .A2(new_n764), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n207), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n211), .B1(new_n765), .B2(G190), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n206), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n780), .A2(new_n782), .A3(new_n273), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n772), .A2(new_n764), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n764), .A2(new_n759), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(G68), .A2(new_n785), .B1(new_n787), .B2(G77), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n771), .A2(new_n778), .A3(new_n783), .A4(new_n788), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n789), .A2(KEYINPUT94), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(KEYINPUT94), .ZN(new_n791));
  INV_X1    g0591(.A(G322), .ZN(new_n792));
  INV_X1    g0592(.A(G311), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n760), .A2(new_n792), .B1(new_n786), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(KEYINPUT33), .B(G317), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n276), .B(new_n794), .C1(new_n785), .C2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n779), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G283), .A2(new_n797), .B1(new_n769), .B2(G329), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G326), .A2(new_n774), .B1(new_n777), .B2(G303), .ZN(new_n799));
  INV_X1    g0599(.A(new_n781), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G294), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n796), .A2(new_n798), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n790), .A2(new_n791), .A3(new_n802), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n751), .B(new_n757), .C1(new_n803), .C2(new_n746), .ZN(new_n804));
  INV_X1    g0604(.A(new_n749), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n685), .B2(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT95), .Z(new_n807));
  INV_X1    g0607(.A(new_n686), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n755), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(G330), .B2(new_n685), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n807), .A2(new_n810), .ZN(G396));
  NAND2_X1  g0611(.A1(new_n745), .A2(new_n748), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT96), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n757), .B1(new_n814), .B2(new_n308), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G87), .A2(new_n797), .B1(new_n769), .B2(G311), .ZN(new_n816));
  INV_X1    g0616(.A(G294), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n273), .C1(new_n817), .C2(new_n760), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n776), .A2(new_n207), .B1(new_n786), .B2(new_n452), .ZN(new_n819));
  INV_X1    g0619(.A(G303), .ZN(new_n820));
  INV_X1    g0620(.A(G283), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n773), .A2(new_n820), .B1(new_n784), .B2(new_n821), .ZN(new_n822));
  NOR4_X1   g0622(.A1(new_n818), .A2(new_n782), .A3(new_n819), .A4(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G137), .A2(new_n774), .B1(new_n787), .B2(G159), .ZN(new_n824));
  INV_X1    g0624(.A(G150), .ZN(new_n825));
  INV_X1    g0625(.A(G143), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n824), .B1(new_n825), .B2(new_n784), .C1(new_n761), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT34), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n273), .B1(new_n777), .B2(G50), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n769), .A2(G132), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n797), .A2(G68), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n800), .A2(G58), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n830), .A2(new_n831), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n827), .B2(new_n828), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n823), .B1(new_n829), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n343), .A2(new_n677), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n326), .A2(new_n323), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n676), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n336), .B2(new_n338), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n838), .B1(new_n841), .B2(new_n344), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n815), .B1(new_n745), .B2(new_n836), .C1(new_n842), .C2(new_n748), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n660), .A2(new_n666), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT87), .B1(new_n652), .B2(new_n656), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n677), .B(new_n842), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(KEYINPUT97), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT97), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n667), .A2(new_n848), .A3(new_n677), .A4(new_n842), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n842), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n733), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n755), .B1(new_n854), .B2(new_n723), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n854), .A2(new_n723), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n843), .B1(new_n856), .B2(new_n857), .ZN(G384));
  OR2_X1    g0658(.A1(new_n359), .A2(new_n361), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT16), .B1(new_n859), .B2(new_n356), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n392), .B1(new_n860), .B2(new_n363), .ZN(new_n861));
  INV_X1    g0661(.A(new_n674), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n402), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n861), .B1(new_n398), .B2(new_n862), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n388), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT37), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n393), .B1(new_n398), .B2(new_n862), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n869), .A2(new_n870), .A3(new_n388), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n865), .A2(KEYINPUT38), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT38), .B1(new_n865), .B2(new_n872), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT99), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n865), .A2(new_n872), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT99), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n865), .A2(KEYINPUT38), .A3(new_n872), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n432), .A2(new_n677), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n436), .A2(new_n445), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n433), .A2(new_n435), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n883), .B1(new_n886), .B2(new_n444), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT102), .B1(new_n718), .B2(new_n720), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT102), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n890), .B(new_n719), .C1(new_n705), .C2(new_n717), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n842), .B(new_n888), .C1(new_n889), .C2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n882), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT40), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n721), .A2(new_n890), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n718), .A2(KEYINPUT102), .A3(new_n720), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n851), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n402), .A2(new_n393), .A3(new_n862), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT100), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n869), .A2(new_n901), .A3(KEYINPUT37), .A4(new_n388), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n370), .B1(new_n397), .B2(new_n674), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT37), .B1(new_n903), .B2(new_n901), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n869), .A2(new_n388), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n900), .A2(new_n902), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n877), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n880), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n899), .A2(new_n909), .A3(KEYINPUT40), .A4(new_n888), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n896), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n897), .A2(new_n898), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n447), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n911), .B(new_n913), .Z(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(G330), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT103), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT98), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n850), .B2(new_n837), .ZN(new_n918));
  AOI211_X1 g0718(.A(KEYINPUT98), .B(new_n838), .C1(new_n847), .C2(new_n849), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n888), .B(new_n882), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT101), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT39), .B1(new_n873), .B2(new_n874), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n909), .B2(KEYINPUT39), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n445), .A2(new_n676), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n923), .A2(new_n924), .B1(new_n628), .B2(new_n674), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n920), .A2(new_n921), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n921), .B1(new_n920), .B2(new_n925), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n447), .A2(new_n735), .A3(new_n732), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n631), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n928), .B(new_n930), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n916), .A2(new_n931), .B1(new_n210), .B2(new_n752), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n916), .B2(new_n931), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n221), .A2(G77), .A3(new_n354), .A4(new_n352), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n201), .A2(G68), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n210), .B(G13), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT35), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n939), .A2(G116), .A3(new_n218), .A4(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT36), .Z(new_n942));
  NOR3_X1   g0742(.A1(new_n933), .A2(new_n936), .A3(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT104), .Z(G367));
  OAI21_X1  g0744(.A(new_n750), .B1(new_n239), .B2(new_n742), .ZN(new_n945));
  INV_X1    g0745(.A(new_n606), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n945), .B1(new_n696), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(G137), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n779), .A2(new_n308), .B1(new_n766), .B2(new_n948), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n273), .B(new_n949), .C1(G58), .C2(new_n777), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n784), .A2(new_n767), .B1(new_n786), .B2(new_n201), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n773), .A2(new_n826), .B1(new_n760), .B2(new_n825), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n781), .A2(new_n203), .ZN(new_n954));
  NOR4_X1   g0754(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n276), .B1(new_n769), .B2(G317), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n777), .A2(G116), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT46), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n956), .B1(new_n207), .B2(new_n781), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  AOI22_X1  g0759(.A1(G294), .A2(new_n785), .B1(new_n787), .B2(G283), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n960), .B1(new_n206), .B2(new_n779), .C1(new_n793), .C2(new_n773), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n959), .B(new_n961), .C1(G303), .C2(new_n762), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n957), .A2(new_n958), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT107), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n955), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n965), .A2(KEYINPUT47), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n745), .B1(new_n965), .B2(KEYINPUT47), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n757), .B(new_n947), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n677), .A2(new_n614), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n970), .A2(new_n636), .A3(new_n644), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT105), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n643), .A2(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n972), .B2(new_n971), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n968), .B1(new_n805), .B2(new_n974), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n724), .B(new_n725), .C1(new_n567), .C2(new_n677), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n649), .A2(new_n677), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n693), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT42), .Z(new_n980));
  INV_X1    g0780(.A(new_n978), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n655), .B1(new_n981), .B2(new_n663), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n677), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n980), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n980), .A2(new_n983), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n974), .B(KEYINPUT43), .Z(new_n987));
  AND3_X1   g0787(.A1(new_n986), .A2(KEYINPUT106), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(KEYINPUT106), .B1(new_n986), .B2(new_n987), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n691), .A2(new_n981), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n991), .B(new_n985), .C1(new_n988), .C2(new_n989), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n978), .A2(new_n694), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT44), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n978), .A2(new_n694), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT45), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n690), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1000), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1002), .A2(new_n691), .A3(new_n997), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n689), .B(new_n692), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n686), .B(new_n1004), .Z(new_n1005));
  NAND4_X1  g0805(.A1(new_n1001), .A2(new_n1003), .A3(new_n736), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n736), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n697), .B(KEYINPUT41), .Z(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n754), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n975), .B1(new_n995), .B2(new_n1010), .ZN(G387));
  INV_X1    g0811(.A(KEYINPUT108), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1005), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n736), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1005), .A2(new_n736), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n697), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n1005), .A2(KEYINPUT108), .A3(new_n736), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n750), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n214), .A2(G107), .ZN(new_n1022));
  AOI211_X1 g0822(.A(G45), .B(new_n701), .C1(G68), .C2(G77), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n253), .A2(G50), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT50), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n742), .B(new_n1026), .C1(new_n236), .C2(G45), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1022), .B(new_n1027), .C1(new_n701), .C2(new_n738), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n760), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G50), .A2(new_n1029), .B1(new_n769), .B2(G150), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n203), .B2(new_n786), .C1(new_n253), .C2(new_n784), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n606), .A2(new_n781), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n276), .B1(new_n779), .B2(new_n206), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n777), .A2(G77), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n767), .B2(new_n773), .ZN(new_n1035));
  NOR4_X1   g0835(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n273), .B1(new_n779), .B2(new_n452), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G322), .A2(new_n774), .B1(new_n787), .B2(G303), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n793), .B2(new_n784), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G317), .B2(new_n762), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1040), .A2(KEYINPUT48), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(KEYINPUT48), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n777), .A2(G294), .B1(new_n800), .B2(G283), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT49), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1037), .B(new_n1046), .C1(G326), .C2(new_n769), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1036), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n756), .B1(new_n1021), .B2(new_n1028), .C1(new_n1049), .C2(new_n745), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n689), .B2(new_n749), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n1005), .B2(new_n754), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1020), .A2(new_n1052), .ZN(G393));
  NAND2_X1  g0853(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n1016), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(new_n1006), .A3(new_n697), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1001), .A2(new_n754), .A3(new_n1003), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G317), .A2(new_n774), .B1(new_n1029), .B2(G311), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT52), .Z(new_n1059));
  AOI22_X1  g0859(.A1(G303), .A2(new_n785), .B1(new_n769), .B2(G322), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G283), .A2(new_n777), .B1(new_n787), .B2(G294), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n276), .B(new_n780), .C1(G116), .C2(new_n800), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n773), .A2(new_n825), .B1(new_n760), .B2(new_n767), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT51), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G68), .A2(new_n777), .B1(new_n769), .B2(G143), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n785), .A2(G50), .B1(new_n787), .B2(new_n310), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n781), .A2(new_n308), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n273), .B(new_n1068), .C1(G87), .C2(new_n797), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n745), .B1(new_n1063), .B2(new_n1070), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n750), .B1(new_n206), .B2(new_n214), .C1(new_n246), .C2(new_n742), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1072), .A2(KEYINPUT109), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1072), .A2(KEYINPUT109), .ZN(new_n1074));
  NOR4_X1   g0874(.A1(new_n1071), .A2(new_n1073), .A3(new_n757), .A4(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n978), .B2(new_n805), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1056), .A2(new_n1057), .A3(new_n1076), .ZN(G390));
  NAND3_X1  g0877(.A1(new_n723), .A2(new_n842), .A3(new_n888), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT110), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1078), .B(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n841), .A2(new_n344), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n838), .B1(new_n731), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n888), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n924), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n909), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n838), .B1(new_n847), .B2(new_n849), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(new_n917), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n924), .B1(new_n1090), .B2(new_n888), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1080), .B(new_n1088), .C1(new_n1091), .C2(new_n923), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n899), .A2(G330), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1093), .A2(new_n1083), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n888), .B1(new_n918), .B2(new_n919), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n923), .B1(new_n1095), .B2(new_n1085), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1094), .B1(new_n1096), .B2(new_n1087), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1092), .A2(new_n1097), .A3(new_n754), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n757), .B1(new_n814), .B2(new_n253), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G283), .A2(new_n774), .B1(new_n787), .B2(G97), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n207), .B2(new_n784), .C1(new_n452), .C2(new_n760), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n273), .B1(new_n776), .B2(new_n314), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n832), .B1(new_n817), .B2(new_n766), .ZN(new_n1103));
  NOR4_X1   g0903(.A1(new_n1101), .A2(new_n1068), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1104), .A2(KEYINPUT112), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT54), .B(G143), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n774), .A2(G128), .B1(new_n787), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n948), .B2(new_n784), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(G132), .ZN(new_n1111));
  INV_X1    g0911(.A(G125), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n760), .A2(new_n1111), .B1(new_n766), .B2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n273), .B(new_n1113), .C1(G50), .C2(new_n797), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n800), .A2(G159), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n776), .A2(new_n825), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT53), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1110), .A2(new_n1114), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1105), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(KEYINPUT112), .B2(new_n1104), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1099), .B1(new_n745), .B2(new_n1120), .C1(new_n923), .C2(new_n748), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1098), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1092), .A2(new_n1097), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT111), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n913), .B2(new_n722), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n447), .A2(new_n912), .A3(KEYINPUT111), .A4(G330), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n930), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n888), .B1(new_n723), .B2(new_n842), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n1094), .A2(new_n1128), .B1(new_n919), .B2(new_n918), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1093), .A2(new_n1083), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1080), .A2(new_n1082), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1127), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n698), .B1(new_n1123), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1092), .A2(new_n1097), .A3(new_n1132), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1122), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(G378));
  NAND2_X1  g0937(.A1(new_n920), .A2(new_n925), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(KEYINPUT101), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n920), .A2(new_n921), .A3(new_n925), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n892), .B1(new_n875), .B2(new_n881), .ZN(new_n1141));
  OAI211_X1 g0941(.A(G330), .B(new_n910), .C1(new_n1141), .C2(KEYINPUT40), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n265), .A2(new_n862), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n302), .B(new_n1143), .Z(new_n1144));
  XOR2_X1   g0944(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1145));
  XNOR2_X1  g0945(.A(new_n1144), .B(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1142), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1146), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n896), .A2(G330), .A3(new_n910), .A4(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1139), .A2(new_n1140), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n926), .B2(new_n927), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1150), .A2(new_n1152), .A3(new_n754), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n755), .B1(new_n813), .B2(G50), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n779), .A2(new_n202), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT113), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1034), .B1(new_n207), .B2(new_n760), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n276), .A2(G41), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1158), .B1(new_n821), .B2(new_n766), .C1(new_n452), .C2(new_n773), .ZN(new_n1159));
  NOR4_X1   g0959(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .A4(new_n954), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n946), .A2(new_n787), .B1(G97), .B2(new_n785), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1161), .A2(KEYINPUT114), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1161), .A2(KEYINPUT114), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1160), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT58), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1158), .ZN(new_n1166));
  INV_X1    g0966(.A(G41), .ZN(new_n1167));
  AOI21_X1  g0967(.A(G50), .B1(new_n250), .B2(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1164), .A2(new_n1165), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT115), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n773), .A2(new_n1112), .B1(new_n784), .B2(new_n1111), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1107), .A2(new_n777), .B1(new_n1029), .B2(G128), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n948), .B2(new_n786), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(G150), .C2(new_n800), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n250), .B(new_n1167), .C1(new_n779), .C2(new_n767), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G124), .B2(new_n769), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT59), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1178), .B1(new_n1174), .B2(new_n1179), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1170), .B1(new_n1165), .B2(new_n1164), .C1(new_n1176), .C2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1154), .B1(new_n1181), .B2(new_n746), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n1148), .B2(new_n748), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1153), .A2(new_n1183), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n930), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1135), .A2(new_n1185), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT57), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT57), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1186), .A2(new_n1187), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1184), .B1(new_n1192), .B2(new_n697), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(G375));
  NAND2_X1  g0994(.A1(new_n1131), .A2(new_n1129), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1195), .A2(new_n1185), .ZN(new_n1196));
  OR3_X1    g0996(.A1(new_n1196), .A2(new_n1132), .A3(new_n1008), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT116), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1083), .A2(new_n747), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n276), .B1(new_n797), .B2(G77), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n452), .B2(new_n784), .C1(new_n817), .C2(new_n773), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n206), .A2(new_n776), .B1(new_n760), .B2(new_n821), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n786), .A2(new_n207), .B1(new_n766), .B2(new_n820), .ZN(new_n1205));
  NOR4_X1   g1005(.A1(new_n1203), .A2(new_n1032), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G132), .A2(new_n774), .B1(new_n785), .B2(new_n1107), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n273), .B1(new_n777), .B2(G159), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n769), .A2(G128), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1156), .B(new_n1210), .C1(G137), .C2(new_n762), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n786), .A2(new_n825), .B1(new_n781), .B2(new_n201), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT117), .Z(new_n1213));
  AOI21_X1  g1013(.A(new_n1206), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n756), .B1(G68), .B2(new_n813), .C1(new_n1214), .C2(new_n745), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT118), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1195), .A2(new_n754), .B1(new_n1201), .B2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1199), .A2(new_n1200), .A3(new_n1217), .ZN(G381));
  OR2_X1    g1018(.A1(G393), .A2(G396), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1219), .A2(G384), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1220), .A2(KEYINPUT119), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1221), .A2(G387), .A3(G390), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(KEYINPUT119), .B2(new_n1220), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1193), .A2(new_n1136), .ZN(new_n1224));
  OR3_X1    g1024(.A1(new_n1223), .A2(new_n1224), .A3(G381), .ZN(G407));
  OAI211_X1 g1025(.A(G407), .B(G213), .C1(G343), .C2(new_n1224), .ZN(G409));
  NAND2_X1  g1026(.A1(new_n1184), .A2(KEYINPUT120), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT120), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1153), .A2(new_n1228), .A3(new_n1183), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1186), .A2(new_n1187), .A3(new_n1009), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1227), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1136), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(KEYINPUT121), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1186), .A2(new_n1187), .A3(new_n1190), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1190), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n697), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1184), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(G378), .A3(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT121), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1231), .A2(new_n1239), .A3(new_n1136), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1233), .A2(new_n1238), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n675), .A2(G213), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1195), .A2(new_n1185), .A3(KEYINPUT60), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT60), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1196), .A2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n697), .B(new_n1133), .C1(new_n1243), .C2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(G384), .A3(new_n1217), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(G384), .B1(new_n1246), .B2(new_n1217), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1241), .A2(new_n1242), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1242), .ZN(new_n1252));
  OAI211_X1 g1052(.A(G2897), .B(new_n1252), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1249), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(G2897), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n1247), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT63), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1251), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(G390), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G387), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT123), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1008), .B1(new_n1006), .B2(new_n736), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n993), .B(new_n994), .C1(new_n1264), .C2(new_n754), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(new_n975), .A3(G390), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1262), .A2(new_n1263), .A3(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(G387), .A2(KEYINPUT123), .A3(new_n1261), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(G393), .B(G396), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT61), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1269), .B1(G387), .B2(new_n1261), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT122), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1266), .A2(new_n1273), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1265), .A2(KEYINPUT122), .A3(new_n975), .A4(G390), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1272), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1270), .A2(new_n1271), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1241), .A2(KEYINPUT63), .A3(new_n1250), .A4(new_n1242), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1279), .A2(KEYINPUT124), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(KEYINPUT124), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1260), .B(new_n1278), .C1(new_n1280), .C2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT126), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT125), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1266), .A2(new_n1263), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G390), .B1(new_n1265), .B2(new_n975), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1276), .B(new_n1284), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1284), .B1(new_n1270), .B2(new_n1276), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1283), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1276), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(KEYINPUT125), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1294), .A2(KEYINPUT126), .A3(new_n1289), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT62), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1241), .A2(new_n1297), .A3(new_n1250), .A4(new_n1242), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1239), .B1(new_n1231), .B2(new_n1136), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1299), .B1(new_n1193), .B2(G378), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1252), .B1(new_n1300), .B2(new_n1240), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1271), .B(new_n1298), .C1(new_n1301), .C2(new_n1257), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1251), .A2(KEYINPUT62), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1296), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1282), .A2(new_n1304), .ZN(G405));
  NAND2_X1  g1105(.A1(new_n1294), .A2(new_n1289), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1193), .A2(new_n1136), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1193), .A2(new_n1136), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1250), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(G375), .A2(G378), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1250), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1310), .A2(new_n1224), .A3(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1306), .A2(new_n1309), .A3(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(KEYINPUT127), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1309), .A2(new_n1312), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1315), .A2(new_n1294), .A3(new_n1289), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT127), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1306), .A2(new_n1309), .A3(new_n1312), .A4(new_n1317), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1314), .A2(new_n1316), .A3(new_n1318), .ZN(G402));
endmodule


