//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT77), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT65), .A2(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT65), .A2(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(G143), .A3(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT64), .A2(G143), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(G146), .A3(new_n195), .ZN(new_n196));
  AND2_X1   g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n191), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT0), .B(G128), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  AND2_X1   g014(.A1(KEYINPUT64), .A2(G143), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT64), .A2(G143), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n200), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  AND2_X1   g017(.A1(KEYINPUT65), .A2(G146), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT65), .A2(G146), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n193), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n199), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n188), .B1(new_n198), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n199), .ZN(new_n209));
  AOI21_X1  g023(.A(G143), .B1(new_n189), .B2(new_n190), .ZN(new_n210));
  AOI21_X1  g024(.A(G146), .B1(new_n194), .B2(new_n195), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n191), .A2(new_n196), .A3(new_n197), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(KEYINPUT77), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216));
  INV_X1    g030(.A(G134), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(G137), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT66), .ZN(new_n219));
  INV_X1    g033(.A(G137), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G134), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(new_n216), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g038(.A(KEYINPUT67), .B(G131), .Z(new_n225));
  OAI21_X1  g039(.A(KEYINPUT68), .B1(new_n220), .B2(G134), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(new_n217), .A3(G137), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n217), .A2(G137), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n226), .A2(new_n228), .B1(new_n229), .B2(KEYINPUT11), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n224), .A2(new_n225), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n224), .A2(new_n230), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n224), .A2(KEYINPUT69), .A3(new_n230), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(G131), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n215), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G128), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(KEYINPUT1), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n191), .A2(new_n196), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT71), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n191), .A2(new_n196), .A3(KEYINPUT71), .A4(new_n239), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G128), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n203), .A2(new_n206), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n242), .A2(new_n243), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT70), .B1(new_n220), .B2(G134), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n221), .ZN(new_n249));
  NOR3_X1   g063(.A1(new_n220), .A2(KEYINPUT70), .A3(G134), .ZN(new_n250));
  OAI21_X1  g064(.A(G131), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n231), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n187), .B1(new_n237), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT76), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT2), .ZN(new_n256));
  INV_X1    g070(.A(G113), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AND3_X1   g072(.A1(KEYINPUT73), .A2(KEYINPUT2), .A3(G113), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT73), .B1(KEYINPUT2), .B2(G113), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT74), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT74), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n263), .B(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n264));
  INV_X1    g078(.A(G119), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G116), .ZN(new_n266));
  INV_X1    g080(.A(G116), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G119), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n262), .A2(KEYINPUT75), .A3(new_n264), .A4(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n261), .A2(new_n269), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n266), .A2(new_n268), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n274), .B1(new_n261), .B2(KEYINPUT74), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT75), .B1(new_n275), .B2(new_n264), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n255), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT75), .ZN(new_n278));
  NAND2_X1  g092(.A1(KEYINPUT2), .A2(G113), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(KEYINPUT73), .A2(KEYINPUT2), .A3(G113), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n281), .A2(new_n282), .B1(new_n256), .B2(new_n257), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n269), .B1(new_n283), .B2(new_n263), .ZN(new_n284));
  INV_X1    g098(.A(new_n264), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n278), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n286), .A2(KEYINPUT76), .A3(new_n272), .A4(new_n270), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n277), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT79), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT79), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n277), .A2(new_n290), .A3(new_n287), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n242), .A2(new_n243), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n245), .A2(new_n246), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n252), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n231), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n235), .A2(G131), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n297), .B1(new_n298), .B2(new_n234), .ZN(new_n299));
  OAI211_X1 g113(.A(KEYINPUT81), .B(new_n296), .C1(new_n299), .C2(new_n215), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n254), .A2(new_n289), .A3(new_n291), .A4(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT28), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT82), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n291), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n296), .B1(new_n299), .B2(new_n215), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n290), .B1(new_n277), .B2(new_n287), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n235), .A2(G131), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT69), .B1(new_n224), .B2(new_n230), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n231), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n212), .A2(new_n213), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n312), .A2(new_n314), .B1(new_n294), .B2(new_n295), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(new_n277), .B2(new_n287), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT28), .B1(new_n309), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n301), .A2(KEYINPUT82), .A3(new_n302), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n305), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT80), .B(KEYINPUT27), .ZN(new_n320));
  INV_X1    g134(.A(G210), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n321), .A2(G237), .A3(G953), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n320), .B(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT26), .B(G101), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT72), .B1(new_n315), .B2(KEYINPUT30), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT72), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT30), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n313), .B1(new_n236), .B2(new_n231), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n328), .B(new_n329), .C1(new_n330), .C2(new_n253), .ZN(new_n331));
  OAI211_X1 g145(.A(KEYINPUT30), .B(new_n296), .C1(new_n299), .C2(new_n215), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n327), .A2(new_n288), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT78), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n309), .ZN(new_n336));
  INV_X1    g150(.A(new_n325), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT29), .B1(new_n326), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G902), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n307), .B1(new_n306), .B2(new_n308), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT28), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(new_n305), .A3(new_n318), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n325), .A2(KEYINPUT29), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n340), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(G472), .B1(new_n339), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n309), .A2(new_n337), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n333), .A2(new_n334), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n333), .A2(new_n334), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT31), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n319), .A2(new_n337), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT31), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n335), .A2(new_n354), .A3(new_n348), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT32), .ZN(new_n357));
  NOR2_X1   g171(.A1(G472), .A2(G902), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n357), .B1(new_n356), .B2(new_n358), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n347), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G214), .B1(G237), .B2(G902), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT6), .ZN(new_n365));
  INV_X1    g179(.A(G101), .ZN(new_n366));
  INV_X1    g180(.A(G104), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n367), .A2(KEYINPUT3), .A3(G107), .ZN(new_n368));
  INV_X1    g182(.A(G107), .ZN(new_n369));
  NAND2_X1  g183(.A1(KEYINPUT88), .A2(G104), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(KEYINPUT88), .A2(G104), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n368), .B1(new_n373), .B2(KEYINPUT3), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT88), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n367), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(G107), .A3(new_n370), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n366), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT4), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT89), .ZN(new_n381));
  INV_X1    g195(.A(new_n368), .ZN(new_n382));
  AOI21_X1  g196(.A(G107), .B1(new_n376), .B2(new_n370), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n377), .A2(new_n366), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n381), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n377), .A2(new_n366), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n374), .A2(new_n388), .A3(KEYINPUT89), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n380), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n379), .B1(new_n390), .B2(new_n378), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n288), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n387), .A2(new_n389), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT92), .B(KEYINPUT5), .ZN(new_n394));
  OAI21_X1  g208(.A(G113), .B1(new_n394), .B2(new_n266), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(new_n274), .B2(new_n394), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(new_n271), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n367), .A2(G107), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n366), .B1(new_n373), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n393), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n392), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G110), .B(G122), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n365), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n401), .B1(new_n288), .B2(new_n391), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n407), .A2(KEYINPUT93), .A3(new_n404), .ZN(new_n408));
  AOI21_X1  g222(.A(KEYINPUT93), .B1(new_n407), .B2(new_n404), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n403), .A2(new_n365), .A3(new_n405), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n313), .A2(G125), .ZN(new_n412));
  OR2_X1    g226(.A1(new_n412), .A2(KEYINPUT94), .ZN(new_n413));
  INV_X1    g227(.A(G125), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n247), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(KEYINPUT94), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G224), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(G953), .ZN(new_n419));
  XOR2_X1   g233(.A(new_n419), .B(KEYINPUT95), .Z(new_n420));
  XNOR2_X1  g234(.A(new_n417), .B(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n410), .A2(new_n411), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n392), .A2(new_n402), .A3(new_n404), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT93), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n407), .A2(KEYINPUT93), .A3(new_n404), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT7), .B1(new_n418), .B2(G953), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n417), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n417), .A2(new_n429), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n399), .B1(new_n387), .B2(new_n389), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n395), .B1(KEYINPUT5), .B2(new_n274), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n432), .B1(new_n271), .B2(new_n433), .ZN(new_n434));
  XOR2_X1   g248(.A(new_n404), .B(KEYINPUT8), .Z(new_n435));
  NOR3_X1   g249(.A1(new_n385), .A2(new_n381), .A3(new_n386), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT89), .B1(new_n374), .B2(new_n388), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n400), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n435), .B1(new_n438), .B2(new_n397), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n430), .A2(new_n431), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(G902), .B1(new_n427), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G210), .B1(G237), .B2(G902), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n422), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n442), .B1(new_n422), .B2(new_n441), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n364), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G217), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(G234), .B2(new_n340), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT87), .ZN(new_n450));
  INV_X1    g264(.A(G110), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n238), .A2(KEYINPUT23), .A3(G119), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n265), .A2(G128), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n265), .A2(G128), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n452), .B(new_n453), .C1(new_n454), .C2(KEYINPUT23), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n451), .B1(new_n455), .B2(KEYINPUT83), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(KEYINPUT83), .B2(new_n455), .ZN(new_n457));
  INV_X1    g271(.A(new_n454), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n458), .A2(new_n453), .ZN(new_n459));
  XOR2_X1   g273(.A(KEYINPUT24), .B(G110), .Z(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G140), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT16), .B1(new_n462), .B2(G125), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(G125), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT84), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n414), .A2(G140), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n462), .A2(KEYINPUT84), .A3(G125), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n463), .B1(new_n469), .B2(KEYINPUT16), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n470), .A2(new_n200), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n470), .A2(new_n200), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n457), .B(new_n461), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  OAI22_X1  g287(.A1(new_n459), .A2(new_n460), .B1(G110), .B2(new_n455), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n204), .A2(new_n205), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n464), .A3(new_n467), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n474), .B(new_n476), .C1(new_n200), .C2(new_n470), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT22), .B(G137), .ZN(new_n478));
  INV_X1    g292(.A(G953), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(G221), .A3(G234), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n478), .B(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n473), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT86), .ZN(new_n483));
  OR2_X1    g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n483), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n481), .B(KEYINPUT85), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(new_n473), .B2(new_n477), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n484), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n450), .B1(new_n488), .B2(new_n340), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n449), .B1(new_n489), .B2(KEYINPUT25), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT25), .ZN(new_n492));
  AOI211_X1 g306(.A(new_n450), .B(new_n492), .C1(new_n488), .C2(new_n340), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n449), .A2(G902), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n491), .A2(new_n494), .B1(new_n488), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n391), .A2(new_n208), .A3(new_n214), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n191), .A2(new_n196), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n498), .B1(new_n499), .B2(new_n238), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n292), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n432), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT10), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(new_n292), .B2(new_n293), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n502), .A2(new_n503), .B1(new_n432), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(KEYINPUT90), .B(new_n231), .C1(new_n310), .C2(new_n311), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT90), .B1(new_n236), .B2(new_n231), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n497), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n438), .A2(new_n247), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n502), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT12), .B1(new_n512), .B2(new_n312), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT12), .ZN(new_n514));
  AOI211_X1 g328(.A(new_n514), .B(new_n299), .C1(new_n511), .C2(new_n502), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n510), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT91), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT91), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n510), .B(new_n518), .C1(new_n513), .C2(new_n515), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(G110), .B(G140), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n479), .A2(G227), .ZN(new_n522));
  XOR2_X1   g336(.A(new_n521), .B(new_n522), .Z(new_n523));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n523), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n510), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n299), .B1(new_n497), .B2(new_n505), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n524), .A2(G469), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G469), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(new_n340), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n497), .A2(new_n505), .A3(new_n509), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n523), .B1(new_n533), .B2(new_n527), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n510), .B(new_n525), .C1(new_n513), .C2(new_n515), .ZN(new_n535));
  AOI21_X1  g349(.A(G902), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n532), .B1(new_n536), .B2(new_n531), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n530), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT9), .B(G234), .ZN(new_n539));
  OAI21_X1  g353(.A(G221), .B1(new_n539), .B2(G902), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n496), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT100), .ZN(new_n542));
  OR3_X1    g356(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT99), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT96), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n201), .A2(new_n202), .ZN(new_n545));
  INV_X1    g359(.A(G237), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n479), .A3(G214), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n544), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n547), .A2(new_n193), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n545), .A2(new_n544), .A3(new_n547), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n225), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n550), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(new_n548), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n225), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n554), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n552), .A2(KEYINPUT17), .A3(new_n553), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT99), .B1(new_n471), .B2(new_n472), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n543), .A2(new_n559), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n552), .A2(KEYINPUT18), .A3(G131), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n469), .A2(G146), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n476), .ZN(new_n565));
  NAND2_X1  g379(.A1(KEYINPUT18), .A2(G131), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n556), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n563), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(G113), .B(G122), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT98), .B(G104), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n570), .B(new_n571), .Z(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n542), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n562), .A2(KEYINPUT100), .A3(new_n568), .A4(new_n572), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT19), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n464), .A2(new_n467), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n469), .B2(KEYINPUT19), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n475), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n580), .B1(new_n200), .B2(new_n470), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT97), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n554), .A2(new_n557), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n581), .A2(KEYINPUT97), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n568), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n573), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n576), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT20), .ZN(new_n589));
  NOR2_X1   g403(.A1(G475), .A2(G902), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n574), .A2(new_n575), .B1(new_n573), .B2(new_n586), .ZN(new_n592));
  INV_X1    g406(.A(new_n590), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT20), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n539), .A2(new_n448), .A3(G953), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n194), .A2(new_n195), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n598), .A2(KEYINPUT101), .A3(new_n238), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT101), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n545), .B2(G128), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n193), .A2(G128), .ZN(new_n603));
  OAI21_X1  g417(.A(G134), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT101), .B1(new_n598), .B2(new_n238), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n545), .A2(new_n600), .A3(G128), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n607), .B(new_n217), .C1(G128), .C2(new_n193), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  OR2_X1    g423(.A1(new_n267), .A2(G122), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n369), .B1(new_n610), .B2(KEYINPUT14), .ZN(new_n611));
  XOR2_X1   g425(.A(G116), .B(G122), .Z(new_n612));
  XOR2_X1   g426(.A(new_n611), .B(new_n612), .Z(new_n613));
  AND2_X1   g427(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT13), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n603), .B1(new_n607), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n602), .A2(KEYINPUT13), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n217), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n612), .B(G107), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n608), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n597), .B1(new_n614), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n609), .A2(new_n613), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n623), .B(new_n596), .C1(new_n618), .C2(new_n620), .ZN(new_n624));
  AOI21_X1  g438(.A(G902), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(G478), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(KEYINPUT15), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n625), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(G234), .A2(G237), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(G952), .A3(new_n479), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n629), .A2(G902), .A3(G953), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT21), .B(G898), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n574), .A2(new_n575), .B1(new_n569), .B2(new_n573), .ZN(new_n637));
  OAI21_X1  g451(.A(G475), .B1(new_n637), .B2(G902), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n595), .A2(new_n628), .A3(new_n636), .A4(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n541), .A2(new_n639), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n362), .A2(new_n447), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(new_n366), .ZN(G3));
  NAND2_X1  g456(.A1(new_n595), .A2(new_n638), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT33), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n622), .B2(new_n624), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n622), .A2(new_n645), .A3(new_n624), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n647), .A2(G478), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n625), .A2(new_n626), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n626), .A2(new_n340), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n644), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n647), .A2(G478), .A3(new_n648), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n655), .A2(KEYINPUT102), .A3(new_n650), .A4(new_n652), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n643), .A2(new_n657), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n363), .B(new_n636), .C1(new_n443), .C2(new_n445), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n496), .A2(new_n538), .A3(new_n540), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n356), .A2(new_n358), .ZN(new_n662));
  INV_X1    g476(.A(G472), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n356), .B2(new_n340), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n660), .A2(new_n661), .A3(new_n662), .A4(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT34), .B(G104), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  NOR3_X1   g482(.A1(new_n659), .A2(new_n628), .A3(new_n643), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n669), .A2(new_n662), .A3(new_n661), .A4(new_n665), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT35), .B(G107), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  INV_X1    g486(.A(new_n486), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(KEYINPUT36), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n473), .A2(new_n477), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n495), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n677), .B1(new_n490), .B2(new_n493), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n525), .B1(new_n517), .B2(new_n519), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n679), .A2(new_n531), .A3(new_n528), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n534), .A2(new_n535), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n531), .A3(new_n340), .ZN(new_n682));
  INV_X1    g496(.A(new_n532), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n678), .B(new_n540), .C1(new_n680), .C2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n639), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n686), .A2(new_n662), .A3(new_n665), .A4(new_n447), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT37), .B(G110), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT103), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n687), .B(new_n689), .ZN(G12));
  INV_X1    g504(.A(new_n447), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n662), .A2(KEYINPUT32), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n359), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n691), .B1(new_n693), .B2(new_n347), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n630), .B(KEYINPUT104), .Z(new_n695));
  OAI21_X1  g509(.A(new_n695), .B1(G900), .B2(new_n632), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NOR4_X1   g511(.A1(new_n685), .A2(new_n643), .A3(new_n628), .A4(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G128), .ZN(G30));
  XNOR2_X1  g514(.A(new_n696), .B(KEYINPUT39), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n538), .A2(new_n540), .A3(new_n701), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n702), .A2(KEYINPUT40), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(KEYINPUT40), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n595), .A2(new_n638), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n628), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n363), .A2(new_n703), .A3(new_n704), .A4(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n678), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n337), .B1(new_n335), .B2(new_n336), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n340), .B1(new_n342), .B2(new_n325), .ZN(new_n710));
  OAI21_X1  g524(.A(G472), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n693), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n444), .A2(new_n446), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT38), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n707), .A2(new_n708), .A3(new_n712), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n598), .ZN(G45));
  NAND3_X1  g530(.A1(new_n643), .A2(new_n657), .A3(new_n696), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n685), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n694), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  INV_X1    g534(.A(new_n496), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n536), .B(G469), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n540), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n362), .A2(new_n660), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT105), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n362), .A2(new_n727), .A3(new_n660), .A4(new_n724), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT41), .B(G113), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  NAND3_X1  g545(.A1(new_n362), .A2(new_n669), .A3(new_n724), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n362), .A2(KEYINPUT106), .A3(new_n669), .A4(new_n724), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G116), .ZN(G18));
  NOR4_X1   g551(.A1(new_n691), .A2(new_n723), .A3(new_n708), .A4(new_n639), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n362), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G119), .ZN(G21));
  NAND2_X1  g554(.A1(new_n706), .A2(new_n447), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n741), .A2(new_n723), .A3(new_n635), .ZN(new_n742));
  INV_X1    g556(.A(new_n358), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n352), .A2(new_n355), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n344), .A2(new_n337), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n664), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n721), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n742), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G122), .ZN(G24));
  NOR4_X1   g565(.A1(new_n717), .A2(new_n746), .A3(new_n664), .A4(new_n708), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n691), .A2(new_n723), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  NOR3_X1   g569(.A1(new_n443), .A2(new_n445), .A3(new_n364), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT107), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n757), .B1(new_n680), .B2(new_n684), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n530), .A2(new_n537), .A3(KEYINPUT107), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n756), .A2(new_n758), .A3(new_n759), .A4(new_n540), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT108), .ZN(new_n761));
  INV_X1    g575(.A(new_n540), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n538), .B2(new_n757), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n763), .A2(new_n764), .A3(new_n756), .A4(new_n759), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n721), .B1(new_n693), .B2(new_n347), .ZN(new_n767));
  INV_X1    g581(.A(new_n717), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT42), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n766), .A2(new_n767), .A3(KEYINPUT42), .A4(new_n768), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G131), .ZN(G33));
  NOR3_X1   g588(.A1(new_n643), .A2(new_n628), .A3(new_n697), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n766), .A2(new_n767), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G134), .ZN(G36));
  INV_X1    g591(.A(KEYINPUT43), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n657), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n705), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n657), .A2(new_n779), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n778), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n705), .A2(KEYINPUT110), .A3(KEYINPUT43), .A4(new_n657), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n657), .A2(KEYINPUT43), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n785), .B1(new_n786), .B2(new_n643), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n708), .B1(new_n783), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n665), .A2(new_n662), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(KEYINPUT44), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT111), .B1(new_n791), .B2(KEYINPUT44), .ZN(new_n795));
  INV_X1    g609(.A(new_n756), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n791), .B2(KEYINPUT44), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT112), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n524), .A2(KEYINPUT45), .A3(new_n529), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT45), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n801), .B1(new_n679), .B2(new_n528), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(G469), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT46), .B1(new_n803), .B2(new_n683), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(new_n531), .B2(new_n536), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n803), .A2(KEYINPUT46), .A3(new_n683), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n762), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n807), .A2(new_n701), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n794), .A2(new_n809), .A3(new_n795), .A4(new_n797), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n799), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  XOR2_X1   g625(.A(KEYINPUT113), .B(G137), .Z(new_n812));
  XNOR2_X1  g626(.A(new_n811), .B(new_n812), .ZN(G39));
  XNOR2_X1  g627(.A(new_n807), .B(KEYINPUT47), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n768), .A2(new_n721), .A3(new_n756), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n815), .A2(new_n362), .A3(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(new_n462), .ZN(G42));
  NOR2_X1   g632(.A1(new_n796), .A2(new_n723), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n631), .A3(new_n496), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(new_n712), .ZN(new_n821));
  INV_X1    g635(.A(new_n658), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(G952), .A3(new_n479), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n783), .A2(new_n788), .ZN(new_n825));
  INV_X1    g639(.A(new_n695), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT116), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n825), .A2(new_n829), .A3(new_n826), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n831), .A2(new_n749), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n824), .B1(new_n832), .B2(new_n753), .ZN(new_n833));
  NOR2_X1   g647(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n819), .ZN(new_n835));
  INV_X1    g649(.A(new_n767), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XOR2_X1   g651(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n838));
  NAND4_X1  g652(.A1(new_n831), .A2(new_n767), .A3(new_n819), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n833), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT119), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n722), .A2(new_n762), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n815), .A2(new_n842), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n843), .A2(KEYINPUT117), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(KEYINPUT117), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n844), .A2(new_n756), .A3(new_n832), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n657), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n821), .A2(new_n705), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n748), .A2(new_n708), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n835), .B2(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n714), .A2(new_n363), .A3(new_n723), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n832), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT50), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n832), .A2(KEYINPUT50), .A3(new_n852), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n851), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n846), .A2(KEYINPUT51), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n843), .A2(new_n832), .A3(new_n756), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n841), .B(new_n858), .C1(new_n860), .C2(KEYINPUT51), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n694), .B1(new_n698), .B2(new_n718), .ZN(new_n862));
  INV_X1    g676(.A(new_n741), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n763), .A2(new_n696), .A3(new_n759), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(new_n712), .A3(new_n864), .A4(new_n708), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n862), .A2(new_n865), .A3(new_n754), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT52), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n766), .A2(new_n752), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n705), .A2(new_n628), .A3(new_n696), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n869), .A2(new_n796), .A3(new_n685), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n362), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n776), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n670), .A2(new_n666), .A3(new_n687), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n641), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n773), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n742), .A2(new_n749), .B1(new_n362), .B2(new_n738), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n729), .A2(new_n876), .A3(new_n736), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT114), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n877), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n766), .A2(new_n752), .B1(new_n362), .B2(new_n870), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n874), .A2(new_n776), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT114), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n879), .A2(new_n881), .A3(new_n882), .A4(new_n773), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n867), .B1(new_n878), .B2(new_n883), .ZN(new_n884));
  XNOR2_X1  g698(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n886), .B(KEYINPUT54), .C1(new_n887), .C2(new_n884), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n875), .A2(new_n887), .A3(new_n877), .ZN(new_n889));
  INV_X1    g703(.A(new_n867), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n885), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n891), .B1(new_n884), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n888), .B1(KEYINPUT54), .B2(new_n893), .ZN(new_n894));
  OAI22_X1  g708(.A1(new_n861), .A2(new_n894), .B1(G952), .B2(G953), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n847), .A2(new_n364), .A3(new_n762), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n705), .A3(new_n496), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n722), .B(KEYINPUT49), .Z(new_n898));
  OR3_X1    g712(.A1(new_n714), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n895), .B1(new_n712), .B2(new_n899), .ZN(G75));
  NOR2_X1   g714(.A1(new_n321), .A2(new_n340), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n893), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT56), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n410), .A2(new_n411), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(new_n421), .Z(new_n905));
  XNOR2_X1  g719(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n905), .B(new_n906), .Z(new_n907));
  NAND3_X1  g721(.A1(new_n902), .A2(new_n903), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n479), .A2(G952), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n893), .A2(new_n912), .A3(new_n901), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n912), .B1(new_n893), .B2(new_n901), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT56), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT122), .B1(new_n915), .B2(new_n907), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n917));
  INV_X1    g731(.A(new_n907), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n902), .A2(KEYINPUT121), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n903), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n917), .B(new_n918), .C1(new_n920), .C2(new_n913), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n911), .B1(new_n916), .B2(new_n921), .ZN(G51));
  XOR2_X1   g736(.A(new_n893), .B(KEYINPUT54), .Z(new_n923));
  XOR2_X1   g737(.A(new_n532), .B(KEYINPUT57), .Z(new_n924));
  OAI21_X1  g738(.A(new_n681), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n893), .ZN(new_n926));
  OR3_X1    g740(.A1(new_n926), .A2(new_n340), .A3(new_n803), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n909), .B1(new_n925), .B2(new_n927), .ZN(G54));
  NAND4_X1  g742(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n929), .A2(new_n592), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n592), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n930), .A2(new_n931), .A3(new_n909), .ZN(G60));
  NAND2_X1  g746(.A1(new_n647), .A2(new_n648), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT123), .ZN(new_n934));
  XNOR2_X1  g748(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n652), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n910), .B1(new_n923), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n934), .B1(new_n894), .B2(new_n936), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(G63));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT60), .Z(new_n942));
  NAND2_X1  g756(.A1(new_n893), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n488), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n909), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT61), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n676), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n945), .B1(new_n948), .B2(new_n943), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  OAI221_X1 g764(.A(new_n945), .B1(new_n946), .B2(KEYINPUT61), .C1(new_n948), .C2(new_n943), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(G66));
  NAND2_X1  g766(.A1(new_n879), .A2(new_n874), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n479), .ZN(new_n954));
  OAI21_X1  g768(.A(G953), .B1(new_n634), .B2(new_n418), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT126), .Z(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(G898), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n904), .B1(new_n958), .B2(G953), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n957), .B(new_n959), .Z(G69));
  NAND3_X1  g774(.A1(new_n327), .A2(new_n332), .A3(new_n331), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(new_n579), .Z(new_n962));
  NAND2_X1  g776(.A1(G900), .A2(G953), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n862), .A2(new_n754), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT127), .Z(new_n965));
  NAND3_X1  g779(.A1(new_n808), .A2(new_n863), .A3(new_n767), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n776), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n817), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n811), .A2(new_n773), .A3(new_n965), .A4(new_n968), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n962), .B(new_n963), .C1(new_n969), .C2(G953), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n965), .A2(new_n715), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n973));
  INV_X1    g787(.A(new_n628), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n822), .B1(new_n974), .B2(new_n705), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n975), .A2(new_n702), .A3(new_n796), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n817), .B1(new_n767), .B2(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n972), .A2(new_n811), .A3(new_n973), .A4(new_n977), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n978), .A2(new_n479), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n970), .B1(new_n979), .B2(new_n962), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n479), .B1(G227), .B2(G900), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(G72));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n978), .B2(new_n953), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n709), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n984), .B1(new_n969), .B2(new_n953), .ZN(new_n987));
  INV_X1    g801(.A(new_n338), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n986), .A2(new_n989), .A3(new_n910), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n884), .A2(new_n887), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n991), .B1(new_n884), .B2(new_n885), .ZN(new_n992));
  INV_X1    g806(.A(new_n984), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n988), .A2(new_n709), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n990), .B1(new_n992), .B2(new_n994), .ZN(G57));
endmodule


