//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT25), .ZN(new_n203));
  NAND2_X1  g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(KEYINPUT23), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(KEYINPUT23), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n205), .A2(new_n209), .A3(KEYINPUT23), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n206), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n203), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n206), .ZN(new_n214));
  INV_X1    g013(.A(new_n210), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n209), .B1(new_n205), .B2(KEYINPUT23), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n214), .B(new_n212), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  AND2_X1   g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(KEYINPUT24), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(KEYINPUT24), .B2(new_n221), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT28), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT27), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G183gat), .ZN(new_n226));
  INV_X1    g025(.A(G183gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT27), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT68), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT68), .B1(new_n227), .B2(KEYINPUT27), .ZN(new_n230));
  INV_X1    g029(.A(G190gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n224), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT69), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n226), .A2(new_n228), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n235), .A2(KEYINPUT28), .A3(new_n231), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n237), .B(new_n224), .C1(new_n229), .C2(new_n232), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n234), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G169gat), .ZN(new_n240));
  INV_X1    g039(.A(G176gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT26), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n204), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT26), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n246), .B1(new_n247), .B2(new_n205), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n221), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n219), .A2(new_n223), .B1(new_n239), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G183gat), .A2(G190gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT24), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n251), .B2(new_n253), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n222), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT67), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n222), .B(new_n258), .C1(new_n254), .C2(new_n255), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n257), .A2(new_n214), .A3(new_n207), .A4(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT25), .ZN(new_n261));
  NAND2_X1  g060(.A1(G226gat), .A2(G233gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT74), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n250), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n239), .A2(new_n249), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT25), .B1(new_n267), .B2(KEYINPUT65), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(new_n223), .A3(new_n217), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n266), .A2(new_n261), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT29), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n264), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G211gat), .ZN(new_n275));
  INV_X1    g074(.A(G218gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G197gat), .ZN(new_n278));
  INV_X1    g077(.A(G204gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(G197gat), .A2(G204gat), .ZN(new_n281));
  OAI22_X1  g080(.A1(KEYINPUT22), .A2(new_n277), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G211gat), .B(G218gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n274), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n283), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n282), .B(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n265), .A2(new_n273), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(G8gat), .B(G36gat), .Z(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(G64gat), .ZN(new_n291));
  XOR2_X1   g090(.A(new_n291), .B(G92gat), .Z(new_n292));
  NAND2_X1  g091(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n292), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n285), .A2(new_n288), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(KEYINPUT30), .A3(new_n295), .ZN(new_n296));
  OR3_X1    g095(.A1(new_n289), .A2(KEYINPUT30), .A3(new_n292), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT79), .ZN(new_n299));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302));
  INV_X1    g101(.A(G155gat), .ZN(new_n303));
  INV_X1    g102(.A(G162gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G148gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G141gat), .ZN(new_n309));
  INV_X1    g108(.A(G141gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G148gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n307), .A2(KEYINPUT76), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT76), .B1(new_n307), .B2(new_n312), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G134gat), .ZN(new_n316));
  INV_X1    g115(.A(G127gat), .ZN(new_n317));
  INV_X1    g116(.A(G120gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G113gat), .ZN(new_n319));
  INV_X1    g118(.A(G113gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G120gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT1), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n317), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AOI211_X1 g123(.A(KEYINPUT1), .B(G127gat), .C1(new_n319), .C2(new_n321), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n316), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n310), .A2(G148gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n308), .A2(G141gat), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT75), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT75), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n309), .A2(new_n311), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(new_n302), .A3(new_n331), .ZN(new_n332));
  AND2_X1   g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G113gat), .B(G120gat), .ZN(new_n337));
  OAI21_X1  g136(.A(G127gat), .B1(new_n337), .B2(KEYINPUT1), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n320), .A2(G120gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n318), .A2(G113gat), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n323), .B(new_n317), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n338), .A2(G134gat), .A3(new_n341), .ZN(new_n342));
  AND4_X1   g141(.A1(new_n315), .A2(new_n326), .A3(new_n336), .A4(new_n342), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n315), .A2(new_n336), .B1(new_n326), .B2(new_n342), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n301), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(KEYINPUT77), .A3(KEYINPUT5), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n347));
  INV_X1    g146(.A(new_n335), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n309), .A2(new_n311), .A3(new_n330), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n330), .B1(new_n309), .B2(new_n311), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n348), .B1(new_n351), .B2(new_n302), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n353));
  INV_X1    g152(.A(new_n312), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n333), .B1(new_n302), .B2(new_n334), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n307), .A2(KEYINPUT76), .A3(new_n312), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n338), .A2(G134gat), .A3(new_n341), .ZN(new_n359));
  AOI21_X1  g158(.A(G134gat), .B1(new_n338), .B2(new_n341), .ZN(new_n360));
  OAI22_X1  g159(.A1(new_n352), .A2(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n315), .A2(new_n326), .A3(new_n336), .A4(new_n342), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n300), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT5), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n347), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n346), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n343), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n362), .A2(KEYINPUT4), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT3), .B1(new_n352), .B2(new_n358), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n326), .A2(new_n342), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT3), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n315), .A2(new_n373), .A3(new_n336), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(new_n300), .A3(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT78), .B1(new_n362), .B2(KEYINPUT4), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n369), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n362), .A2(KEYINPUT78), .A3(KEYINPUT4), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n375), .A2(new_n364), .A3(new_n300), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n366), .A2(new_n376), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G1gat), .B(G29gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(KEYINPUT0), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(G57gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(G85gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n299), .B1(new_n383), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n375), .A2(new_n300), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n346), .A2(new_n365), .B1(new_n390), .B2(new_n370), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n381), .B1(new_n378), .B2(new_n379), .ZN(new_n392));
  NOR4_X1   g191(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT79), .A4(new_n387), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n389), .A2(new_n393), .A3(KEYINPUT6), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT80), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT77), .B1(new_n345), .B2(KEYINPUT5), .ZN(new_n396));
  NOR3_X1   g195(.A1(new_n363), .A2(new_n347), .A3(new_n364), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n376), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n382), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n395), .B1(new_n400), .B2(new_n387), .ZN(new_n401));
  AOI211_X1 g200(.A(KEYINPUT80), .B(new_n388), .C1(new_n398), .C2(new_n399), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n394), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n400), .A2(KEYINPUT6), .A3(new_n387), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n298), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n315), .A2(new_n336), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n284), .A2(KEYINPUT29), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT81), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n373), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n287), .A2(new_n271), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(KEYINPUT81), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n407), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n287), .B1(new_n374), .B2(new_n271), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n414), .B1(G228gat), .B2(G233gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n411), .A2(new_n373), .B1(new_n315), .B2(new_n336), .ZN(new_n417));
  OAI211_X1 g216(.A(G228gat), .B(G233gat), .C1(new_n417), .C2(new_n414), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT31), .B(G50gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n420), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n416), .A2(new_n422), .A3(new_n418), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G78gat), .B(G106gat), .ZN(new_n425));
  XOR2_X1   g224(.A(new_n425), .B(G22gat), .Z(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n421), .A2(new_n426), .A3(new_n423), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G227gat), .A2(G233gat), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n372), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n433), .B1(new_n250), .B2(new_n261), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n266), .A2(new_n261), .A3(new_n269), .A4(new_n433), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n432), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G15gat), .B(G43gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(G71gat), .ZN(new_n439));
  INV_X1    g238(.A(G99gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT33), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n437), .A2(KEYINPUT32), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n270), .A2(new_n372), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n431), .B1(new_n444), .B2(new_n435), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n441), .B1(new_n445), .B2(KEYINPUT33), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT32), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g247(.A(KEYINPUT71), .B(new_n443), .C1(new_n446), .C2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n444), .A2(new_n431), .A3(new_n435), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT34), .B1(new_n450), .B2(KEYINPUT72), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT72), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n444), .A2(new_n452), .A3(new_n431), .A4(new_n435), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n453), .A2(KEYINPUT73), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(KEYINPUT73), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n451), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n450), .A2(KEYINPUT72), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT34), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n434), .A2(new_n436), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT73), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n460), .A2(new_n452), .A3(new_n461), .A4(new_n431), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n453), .A2(KEYINPUT73), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n437), .A2(KEYINPUT32), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT33), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n437), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT71), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n465), .A2(new_n467), .A3(new_n468), .A4(new_n441), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n449), .A2(new_n456), .A3(new_n464), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n449), .A2(new_n469), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n464), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n430), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n202), .B1(new_n406), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n296), .A2(new_n297), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n473), .A2(new_n470), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n398), .A2(new_n388), .A3(new_n399), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT79), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n387), .B1(new_n391), .B2(new_n392), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n398), .A2(new_n299), .A3(new_n388), .A4(new_n399), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT35), .B1(new_n483), .B2(new_n405), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n428), .A2(new_n429), .ZN(new_n485));
  AND4_X1   g284(.A1(new_n476), .A2(new_n477), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n475), .A2(new_n486), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n473), .A2(KEYINPUT36), .A3(new_n470), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT36), .B1(new_n473), .B2(new_n470), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n481), .A2(KEYINPUT80), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n400), .A2(new_n395), .A3(new_n387), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n405), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n476), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n430), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT82), .B1(new_n490), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n499));
  INV_X1    g298(.A(new_n470), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n449), .A2(new_n469), .B1(new_n456), .B2(new_n464), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n473), .A2(KEYINPUT36), .A3(new_n470), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT82), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n485), .B1(new_n495), .B2(new_n476), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n498), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n294), .B1(new_n289), .B2(KEYINPUT37), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n509), .A2(KEYINPUT85), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n289), .A2(KEYINPUT37), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n511), .A2(KEYINPUT85), .A3(new_n292), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT37), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n285), .A2(new_n288), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT38), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT38), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n509), .A2(new_n517), .A3(new_n514), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n483), .A2(new_n405), .A3(new_n518), .A4(new_n295), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT84), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n519), .A2(new_n520), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n516), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n300), .B1(new_n380), .B2(new_n375), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT39), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n343), .A2(new_n344), .A3(new_n301), .ZN(new_n526));
  OR3_X1    g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n525), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n527), .A2(KEYINPUT40), .A3(new_n388), .A4(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT83), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n527), .A2(new_n388), .A3(new_n528), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT40), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n531), .A2(new_n481), .A3(new_n298), .A4(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n523), .A2(new_n485), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n487), .B1(new_n508), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G230gat), .A2(G233gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(G106gat), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT8), .B1(new_n440), .B2(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(KEYINPUT93), .B(G92gat), .Z(new_n542));
  OAI21_X1  g341(.A(new_n541), .B1(new_n542), .B2(G85gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT94), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G85gat), .A2(G92gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT7), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(G99gat), .B(G106gat), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(G57gat), .B(G64gat), .Z(new_n551));
  INV_X1    g350(.A(G71gat), .ZN(new_n552));
  INV_X1    g351(.A(G78gat), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n551), .B1(KEYINPUT9), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G71gat), .B(G78gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n549), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n545), .A2(new_n558), .A3(new_n547), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n550), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n557), .B1(new_n550), .B2(new_n559), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n539), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n563), .A2(KEYINPUT100), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(KEYINPUT100), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT99), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT10), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n562), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n560), .A2(new_n566), .A3(KEYINPUT10), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n569), .A2(new_n538), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n564), .A2(new_n565), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G120gat), .B(G148gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(new_n241), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(new_n279), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n576), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n564), .A2(new_n578), .A3(new_n572), .A4(new_n565), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n581), .B(KEYINPUT89), .Z(new_n582));
  XNOR2_X1  g381(.A(G15gat), .B(G22gat), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT16), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n583), .B1(new_n584), .B2(G1gat), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n585), .B1(G1gat), .B2(new_n583), .ZN(new_n586));
  INV_X1    g385(.A(G8gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G43gat), .B(G50gat), .Z(new_n589));
  INV_X1    g388(.A(KEYINPUT15), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(G29gat), .ZN(new_n592));
  INV_X1    g391(.A(G36gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(KEYINPUT14), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT14), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(G29gat), .B2(G36gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n591), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(KEYINPUT88), .ZN(new_n600));
  INV_X1    g399(.A(new_n594), .ZN(new_n601));
  INV_X1    g400(.A(new_n591), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n589), .A2(new_n590), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n588), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n599), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT17), .ZN(new_n607));
  AOI211_X1 g406(.A(new_n582), .B(new_n605), .C1(new_n607), .C2(new_n588), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT18), .B1(new_n608), .B2(KEYINPUT90), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT90), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT18), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n588), .ZN(new_n612));
  INV_X1    g411(.A(new_n605), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n610), .B(new_n611), .C1(new_n614), .C2(new_n582), .ZN(new_n615));
  INV_X1    g414(.A(new_n588), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(new_n606), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n582), .B(KEYINPUT13), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n609), .A2(new_n615), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(KEYINPUT86), .B(KEYINPUT11), .Z(new_n622));
  XNOR2_X1  g421(.A(G113gat), .B(G141gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G169gat), .B(G197gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(KEYINPUT87), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n621), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT91), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n621), .A2(KEYINPUT91), .A3(new_n628), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n609), .A2(new_n615), .A3(new_n627), .A4(new_n620), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n633), .A2(KEYINPUT92), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(KEYINPUT92), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n631), .B(new_n632), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n537), .A2(new_n580), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n550), .A2(new_n559), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n607), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT95), .ZN(new_n641));
  AND2_X1   g440(.A1(G232gat), .A2(G233gat), .ZN(new_n642));
  AOI22_X1  g441(.A1(new_n640), .A2(new_n641), .B1(KEYINPUT41), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n607), .A2(KEYINPUT95), .A3(new_n639), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n550), .A2(new_n559), .A3(new_n606), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(G190gat), .B(G218gat), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT97), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n642), .A2(KEYINPUT41), .ZN(new_n651));
  XNOR2_X1  g450(.A(G134gat), .B(G162gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n646), .A2(new_n654), .A3(new_n648), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n643), .A2(new_n644), .A3(new_n647), .A4(new_n645), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n650), .A2(new_n653), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(KEYINPUT98), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n660), .A2(KEYINPUT96), .A3(new_n647), .A4(new_n645), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT96), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n650), .A2(new_n661), .A3(new_n655), .A4(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n653), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n659), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n658), .B1(new_n666), .B2(new_n657), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n557), .A2(KEYINPUT21), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G127gat), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n616), .B1(KEYINPUT21), .B2(new_n557), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n672));
  XNOR2_X1  g471(.A(G155gat), .B(G183gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n671), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(G231gat), .A2(G233gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(new_n275), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n675), .B(new_n677), .Z(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n667), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n638), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n495), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g484(.A(new_n587), .B1(new_n682), .B2(new_n298), .ZN(new_n686));
  NOR2_X1   g485(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n584), .A2(new_n587), .ZN(new_n688));
  NOR4_X1   g487(.A1(new_n681), .A2(new_n476), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT42), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(KEYINPUT42), .B2(new_n689), .ZN(G1325gat));
  AND3_X1   g490(.A1(new_n682), .A2(G15gat), .A3(new_n504), .ZN(new_n692));
  AOI21_X1  g491(.A(G15gat), .B1(new_n682), .B2(new_n477), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(G1326gat));
  NOR2_X1   g493(.A1(new_n681), .A2(new_n485), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT43), .B(G22gat), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  INV_X1    g496(.A(new_n667), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n637), .A2(new_n678), .A3(new_n580), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n537), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n592), .A3(new_n683), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n699), .A2(KEYINPUT101), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT44), .B1(new_n537), .B2(new_n698), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n490), .A2(new_n497), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n483), .A2(new_n405), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n711), .A2(KEYINPUT84), .A3(new_n295), .A4(new_n518), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n519), .A2(new_n520), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n430), .B1(new_n714), .B2(new_n516), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n710), .B1(new_n715), .B2(new_n535), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT102), .B1(new_n475), .B2(new_n486), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n477), .A2(new_n485), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT35), .B1(new_n718), .B2(new_n496), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT102), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n474), .A2(new_n476), .A3(new_n484), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n709), .B(new_n667), .C1(new_n716), .C2(new_n723), .ZN(new_n724));
  AOI211_X1 g523(.A(KEYINPUT103), .B(new_n707), .C1(new_n708), .C2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n505), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n504), .A2(new_n506), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT82), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n536), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n487), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n698), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n724), .B1(new_n733), .B2(new_n709), .ZN(new_n734));
  INV_X1    g533(.A(new_n707), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n727), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n495), .B1(new_n726), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n703), .B1(new_n738), .B2(new_n592), .ZN(G1328gat));
  NAND3_X1  g538(.A1(new_n701), .A2(new_n593), .A3(new_n298), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT46), .Z(new_n741));
  AOI21_X1  g540(.A(new_n476), .B1(new_n726), .B2(new_n737), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n742), .B2(new_n593), .ZN(G1329gat));
  NAND2_X1  g542(.A1(new_n733), .A2(new_n699), .ZN(new_n744));
  INV_X1    g543(.A(new_n477), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n744), .A2(G43gat), .A3(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n734), .A2(new_n504), .A3(new_n735), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n747), .B2(G43gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT47), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n504), .B1(new_n725), .B2(new_n736), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n746), .B1(new_n750), .B2(G43gat), .ZN(new_n751));
  XNOR2_X1  g550(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n749), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n749), .B(KEYINPUT105), .C1(new_n751), .C2(new_n752), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(G1330gat));
  INV_X1    g556(.A(G50gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n701), .A2(new_n758), .A3(new_n430), .ZN(new_n759));
  AOI211_X1 g558(.A(new_n485), .B(new_n707), .C1(new_n708), .C2(new_n724), .ZN(new_n760));
  OAI211_X1 g559(.A(KEYINPUT48), .B(new_n759), .C1(new_n760), .C2(new_n758), .ZN(new_n761));
  INV_X1    g560(.A(new_n759), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n430), .B1(new_n725), .B2(new_n736), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(new_n763), .B2(G50gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n761), .B1(new_n764), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g564(.A1(new_n536), .A2(new_n729), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n766), .A2(new_n717), .A3(new_n722), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n667), .A2(new_n679), .A3(new_n636), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n767), .A2(new_n580), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n495), .ZN(new_n770));
  XOR2_X1   g569(.A(KEYINPUT106), .B(G57gat), .Z(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1332gat));
  NOR2_X1   g571(.A1(new_n769), .A2(new_n476), .ZN(new_n773));
  NOR2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  AND2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n773), .B2(new_n774), .ZN(G1333gat));
  OAI21_X1  g576(.A(new_n552), .B1(new_n769), .B2(new_n745), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n504), .A2(G71gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n769), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g580(.A1(new_n769), .A2(new_n485), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(new_n553), .ZN(G1335gat));
  NOR2_X1   g582(.A1(new_n636), .A2(new_n678), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n667), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n767), .A2(KEYINPUT51), .A3(new_n667), .A4(new_n784), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n785), .A2(KEYINPUT107), .A3(new_n786), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n580), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n793), .A2(new_n495), .A3(G85gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n734), .A2(new_n580), .A3(new_n784), .ZN(new_n796));
  OAI21_X1  g595(.A(G85gat), .B1(new_n796), .B2(new_n495), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(G1336gat));
  NAND3_X1  g597(.A1(new_n787), .A2(KEYINPUT108), .A3(new_n789), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n793), .A2(G92gat), .A3(new_n476), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT108), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n801), .A3(new_n786), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n799), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n734), .A2(new_n580), .A3(new_n298), .A4(new_n784), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n804), .A2(new_n542), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT52), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT52), .B1(new_n792), .B2(new_n800), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n804), .A2(new_n808), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(new_n542), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT110), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n807), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(new_n807), .B2(new_n811), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n806), .B1(new_n813), .B2(new_n814), .ZN(G1337gat));
  OAI21_X1  g614(.A(G99gat), .B1(new_n796), .B2(new_n490), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n792), .A2(new_n440), .A3(new_n477), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(new_n793), .ZN(G1338gat));
  OAI21_X1  g617(.A(G106gat), .B1(new_n796), .B2(new_n485), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n793), .A2(G106gat), .A3(new_n485), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n799), .A2(new_n802), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT53), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n790), .A2(new_n791), .A3(new_n820), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n819), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT111), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n823), .A2(new_n829), .A3(new_n826), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(G1339gat));
  NAND2_X1  g630(.A1(new_n666), .A2(new_n657), .ZN(new_n832));
  INV_X1    g631(.A(new_n658), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n614), .A2(new_n582), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n617), .A2(new_n619), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n834), .B1(new_n837), .B2(new_n626), .ZN(new_n838));
  INV_X1    g637(.A(new_n626), .ZN(new_n839));
  AOI211_X1 g638(.A(KEYINPUT112), .B(new_n839), .C1(new_n835), .C2(new_n836), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n633), .A2(KEYINPUT92), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n633), .A2(KEYINPUT92), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n572), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n578), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n539), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(KEYINPUT54), .A3(new_n572), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n848), .A2(KEYINPUT55), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT55), .B1(new_n848), .B2(new_n851), .ZN(new_n853));
  INV_X1    g652(.A(new_n579), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n832), .A2(new_n833), .A3(new_n845), .A4(new_n855), .ZN(new_n856));
  AOI22_X1  g655(.A1(new_n845), .A2(new_n580), .B1(new_n855), .B2(new_n636), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(new_n667), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n679), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n768), .A2(new_n793), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n861), .A2(new_n683), .A3(new_n476), .A4(new_n474), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n862), .B(new_n863), .ZN(new_n864));
  OR3_X1    g663(.A1(new_n864), .A2(G113gat), .A3(new_n637), .ZN(new_n865));
  OAI21_X1  g664(.A(G113gat), .B1(new_n862), .B2(new_n637), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT114), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n865), .A2(new_n869), .A3(new_n866), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1340gat));
  OAI21_X1  g670(.A(G120gat), .B1(new_n862), .B2(new_n793), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n580), .A2(new_n318), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n864), .B2(new_n873), .ZN(G1341gat));
  NOR2_X1   g673(.A1(new_n862), .A2(new_n679), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(G127gat), .ZN(new_n876));
  XOR2_X1   g675(.A(new_n876), .B(KEYINPUT115), .Z(new_n877));
  INV_X1    g676(.A(new_n875), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n317), .B2(new_n878), .ZN(G1342gat));
  OR2_X1    g678(.A1(new_n862), .A2(new_n698), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(G134gat), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT116), .Z(new_n882));
  NOR2_X1   g681(.A1(new_n880), .A2(G134gat), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT56), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(G1343gat));
  AOI22_X1  g684(.A1(new_n858), .A2(new_n679), .B1(new_n768), .B2(new_n793), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(new_n485), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n504), .A2(new_n495), .A3(new_n298), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n889), .A2(G141gat), .A3(new_n637), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(KEYINPUT58), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n855), .A2(new_n636), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n580), .B(new_n841), .C1(new_n634), .C2(new_n635), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n843), .A2(new_n844), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n896), .A2(KEYINPUT118), .A3(new_n580), .A4(new_n841), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n892), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n698), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(KEYINPUT119), .A3(new_n856), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n898), .A2(new_n698), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n900), .A2(new_n679), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n485), .B1(new_n903), .B2(new_n860), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n861), .A2(new_n430), .ZN(new_n905));
  XOR2_X1   g704(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n904), .A2(KEYINPUT57), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n888), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n908), .A2(new_n637), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n891), .B1(new_n910), .B2(new_n310), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n890), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n903), .A2(new_n860), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(KEYINPUT57), .A3(new_n430), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n905), .A2(new_n907), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT120), .B1(new_n917), .B2(new_n888), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n919));
  AOI211_X1 g718(.A(new_n919), .B(new_n909), .C1(new_n915), .C2(new_n916), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n636), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n913), .B1(new_n921), .B2(G141gat), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT58), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n911), .B1(new_n922), .B2(new_n923), .ZN(G1344gat));
  INV_X1    g723(.A(new_n889), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n308), .A3(new_n580), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT122), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n919), .B1(new_n908), .B2(new_n909), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n917), .A2(KEYINPUT120), .A3(new_n888), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n793), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n930), .A2(KEYINPUT59), .A3(new_n308), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n667), .A2(new_n855), .ZN(new_n932));
  AOI22_X1  g731(.A1(new_n932), .A2(new_n845), .B1(new_n698), .B2(new_n898), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n860), .B1(new_n933), .B2(new_n678), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT57), .B1(new_n934), .B2(new_n430), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n886), .A2(new_n485), .A3(new_n907), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n580), .B(new_n888), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G148gat), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT59), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT123), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n941), .A3(KEYINPUT59), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n927), .B1(new_n931), .B2(new_n943), .ZN(G1345gat));
  NOR2_X1   g743(.A1(new_n918), .A2(new_n920), .ZN(new_n945));
  OAI21_X1  g744(.A(G155gat), .B1(new_n945), .B2(new_n679), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n925), .A2(new_n303), .A3(new_n678), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1346gat));
  OAI21_X1  g747(.A(G162gat), .B1(new_n945), .B2(new_n698), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n889), .A2(G162gat), .A3(new_n698), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT124), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1347gat));
  NOR2_X1   g751(.A1(new_n683), .A2(new_n476), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n861), .A2(new_n474), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n954), .A2(new_n637), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(new_n240), .ZN(G1348gat));
  NOR2_X1   g755(.A1(new_n954), .A2(new_n793), .ZN(new_n957));
  XOR2_X1   g756(.A(KEYINPUT125), .B(G176gat), .Z(new_n958));
  XNOR2_X1  g757(.A(new_n957), .B(new_n958), .ZN(G1349gat));
  NOR2_X1   g758(.A1(new_n954), .A2(new_n679), .ZN(new_n960));
  MUX2_X1   g759(.A(G183gat), .B(new_n235), .S(new_n960), .Z(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT60), .ZN(G1350gat));
  XNOR2_X1  g761(.A(KEYINPUT61), .B(G190gat), .ZN(new_n963));
  NAND2_X1  g762(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n954), .A2(new_n698), .ZN(new_n965));
  MUX2_X1   g764(.A(new_n963), .B(new_n964), .S(new_n965), .Z(G1351gat));
  NAND2_X1  g765(.A1(new_n490), .A2(new_n953), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n887), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT126), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n970), .A2(new_n278), .A3(new_n636), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n935), .A2(new_n936), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n972), .A2(new_n967), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(new_n636), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n971), .B1(new_n975), .B2(new_n278), .ZN(G1352gat));
  NOR3_X1   g775(.A1(new_n969), .A2(G204gat), .A3(new_n793), .ZN(new_n977));
  INV_X1    g776(.A(new_n977), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n978), .A2(KEYINPUT127), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n978), .A2(KEYINPUT127), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT62), .ZN(new_n981));
  OR3_X1    g780(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n580), .B1(new_n935), .B2(new_n936), .ZN(new_n983));
  OAI21_X1  g782(.A(G204gat), .B1(new_n983), .B2(new_n967), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n981), .B1(new_n979), .B2(new_n980), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n982), .A2(new_n984), .A3(new_n985), .ZN(G1353gat));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n275), .A3(new_n678), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n973), .A2(new_n678), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n988), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n989));
  AOI21_X1  g788(.A(KEYINPUT63), .B1(new_n988), .B2(G211gat), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n987), .B1(new_n989), .B2(new_n990), .ZN(G1354gat));
  AOI21_X1  g790(.A(G218gat), .B1(new_n970), .B2(new_n667), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n698), .A2(new_n276), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n992), .B1(new_n973), .B2(new_n993), .ZN(G1355gat));
endmodule


