//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n567, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n616,
    new_n617, new_n620, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  NOR3_X1   g043(.A1(new_n468), .A2(new_n462), .A3(G2105), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT67), .B1(new_n470), .B2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G101), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT66), .B1(new_n460), .B2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(new_n461), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n460), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n474), .A2(new_n475), .A3(G137), .A4(new_n470), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n467), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT68), .Z(G160));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT70), .Z(new_n481));
  NAND2_X1  g056(.A1(new_n474), .A2(new_n475), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n474), .A2(KEYINPUT69), .A3(new_n475), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n486), .A2(new_n470), .ZN(new_n489));
  AOI211_X1 g064(.A(new_n481), .B(new_n488), .C1(G124), .C2(new_n489), .ZN(G162));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n470), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n495), .A2(new_n497), .A3(KEYINPUT71), .A4(G2104), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n470), .A2(KEYINPUT4), .A3(G138), .ZN(new_n500));
  NAND2_X1  g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n474), .A2(new_n475), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n461), .A2(new_n463), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n470), .A2(G138), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n499), .A2(new_n503), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G62), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT73), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G543), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n518), .A2(new_n519), .A3(G62), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n516), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G651), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT74), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT72), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT6), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n526), .B2(G651), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(KEYINPUT72), .A3(KEYINPUT6), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n526), .A2(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n530), .A2(new_n531), .A3(new_n518), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n530), .A2(G543), .A3(new_n531), .ZN(new_n534));
  AOI22_X1  g109(.A1(G88), .A2(new_n533), .B1(new_n534), .B2(G50), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n521), .A2(KEYINPUT74), .A3(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n524), .A2(new_n535), .A3(new_n536), .ZN(G303));
  INV_X1    g112(.A(G303), .ZN(G166));
  NAND2_X1  g113(.A1(new_n514), .A2(KEYINPUT75), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT75), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n518), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n542), .A2(G63), .A3(G651), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT76), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n533), .A2(G89), .ZN(new_n546));
  NAND3_X1  g121(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n547));
  XOR2_X1   g122(.A(new_n547), .B(KEYINPUT7), .Z(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n534), .A2(G51), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n545), .A2(new_n546), .A3(new_n549), .A4(new_n550), .ZN(G286));
  INV_X1    g126(.A(G286), .ZN(G168));
  NAND2_X1  g127(.A1(new_n542), .A2(G64), .ZN(new_n553));
  NAND2_X1  g128(.A1(G77), .A2(G543), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n528), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(G52), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n530), .A2(G543), .A3(new_n531), .ZN(new_n557));
  INV_X1    g132(.A(G90), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n556), .A2(new_n557), .B1(new_n532), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n555), .A2(new_n559), .ZN(G171));
  AOI22_X1  g135(.A1(new_n542), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(new_n528), .ZN(new_n562));
  AOI22_X1  g137(.A1(G81), .A2(new_n533), .B1(new_n534), .B2(G43), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(G188));
  NAND2_X1  g146(.A1(new_n534), .A2(G53), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n533), .A2(G91), .ZN(new_n574));
  AND2_X1   g149(.A1(new_n518), .A2(G65), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT77), .Z(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n573), .A2(new_n574), .A3(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  AOI22_X1  g155(.A1(G87), .A2(new_n533), .B1(new_n534), .B2(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n542), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  NAND3_X1  g158(.A1(new_n511), .A2(new_n513), .A3(G61), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(KEYINPUT78), .B1(new_n534), .B2(G48), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n528), .B1(new_n584), .B2(new_n585), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n533), .A2(G86), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n588), .A2(new_n591), .ZN(G305));
  INV_X1    g167(.A(G47), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n593), .A2(new_n557), .B1(new_n532), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT79), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n542), .A2(G60), .ZN(new_n597));
  AND2_X1   g172(.A1(G72), .A2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n596), .A2(new_n599), .ZN(G290));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  OR3_X1    g176(.A1(new_n532), .A2(KEYINPUT10), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n514), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n534), .A2(G54), .B1(new_n605), .B2(G651), .ZN(new_n606));
  OAI21_X1  g181(.A(KEYINPUT10), .B1(new_n532), .B2(new_n601), .ZN(new_n607));
  AND3_X1   g182(.A1(new_n602), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(new_n610), .B2(G171), .ZN(G284));
  OAI21_X1  g187(.A(new_n611), .B1(new_n610), .B2(G171), .ZN(G321));
  NOR2_X1   g188(.A1(G168), .A2(new_n610), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(KEYINPUT80), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(G299), .B2(new_n610), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n615), .B1(new_n614), .B2(new_n617), .ZN(G297));
  OAI21_X1  g193(.A(new_n615), .B1(new_n614), .B2(new_n617), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n608), .B1(new_n620), .B2(G860), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT81), .Z(G148));
  NAND2_X1  g197(.A1(new_n564), .A2(new_n610), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n609), .A2(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(new_n610), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g201(.A1(new_n469), .A2(new_n471), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n627), .A2(new_n461), .A3(new_n463), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT12), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(G2100), .Z(new_n631));
  NAND2_X1  g206(.A1(new_n489), .A2(G123), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n487), .A2(G135), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n634), .A2(KEYINPUT82), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(KEYINPUT82), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n635), .B(new_n636), .C1(G111), .C2(new_n470), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n632), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n631), .A2(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT86), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2427), .B(G2430), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(KEYINPUT14), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT85), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n646), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G1341), .B(G1348), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT84), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n651), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(G14), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT87), .Z(new_n660));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(KEYINPUT17), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n662), .B(new_n664), .C1(new_n660), .C2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n661), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n667), .A2(new_n659), .A3(new_n663), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT18), .Z(new_n669));
  NAND3_X1  g244(.A1(new_n660), .A2(new_n665), .A3(new_n663), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n666), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2096), .B(G2100), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(new_n676), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n678), .A2(new_n680), .A3(new_n682), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n685), .B(new_n686), .C1(new_n684), .C2(new_n683), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  INV_X1    g265(.A(G1981), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G1986), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n689), .B(new_n693), .Z(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G229));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G22), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G166), .B2(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(G1971), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(G16), .A2(G23), .ZN(new_n701));
  INV_X1    g276(.A(G288), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(G16), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT33), .B(G1976), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(G6), .A2(G16), .ZN(new_n706));
  INV_X1    g281(.A(G305), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(G16), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT32), .B(G1981), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n700), .A2(new_n705), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT34), .ZN(new_n712));
  OR2_X1    g287(.A1(G16), .A2(G24), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G290), .B2(new_n696), .ZN(new_n714));
  INV_X1    g289(.A(G1986), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n714), .A2(new_n715), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n489), .A2(G119), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n487), .A2(G131), .ZN(new_n720));
  OR2_X1    g295(.A1(G95), .A2(G2105), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n721), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G29), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT88), .ZN(new_n726));
  OR2_X1    g301(.A1(G25), .A2(G29), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT35), .B(G1991), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n726), .B1(new_n725), .B2(new_n727), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n729), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n732), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n730), .B1(new_n734), .B2(new_n728), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n717), .B(new_n718), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n712), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(KEYINPUT89), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT89), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n737), .A2(new_n741), .A3(new_n738), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n740), .B(new_n742), .C1(new_n738), .C2(new_n737), .ZN(new_n743));
  NOR2_X1   g318(.A1(G5), .A2(G16), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G171), .B2(G16), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G1961), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT96), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(G160), .A2(G29), .ZN(new_n749));
  INV_X1    g324(.A(G29), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT24), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(G34), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(KEYINPUT93), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(G34), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(KEYINPUT93), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n749), .B1(KEYINPUT94), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(KEYINPUT94), .B2(new_n756), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n748), .B1(new_n758), .B2(G2084), .ZN(new_n759));
  NOR2_X1   g334(.A1(G29), .A2(G35), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G162), .B2(G29), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT29), .B(G2090), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n627), .A2(G105), .ZN(new_n764));
  NAND3_X1  g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT26), .ZN(new_n766));
  AOI211_X1 g341(.A(new_n764), .B(new_n766), .C1(new_n487), .C2(G141), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n489), .A2(G129), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(G29), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G29), .B2(G32), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT27), .B(G1996), .Z(new_n774));
  AOI211_X1 g349(.A(new_n759), .B(new_n763), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT23), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n696), .A2(G20), .ZN(new_n777));
  AOI22_X1  g352(.A1(G299), .A2(G16), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n776), .B2(new_n777), .ZN(new_n779));
  INV_X1    g354(.A(G1956), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT30), .B(G28), .Z(new_n782));
  OAI221_X1 g357(.A(new_n781), .B1(G29), .B2(new_n782), .C1(G1961), .C2(new_n745), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n638), .A2(new_n750), .ZN(new_n784));
  NOR2_X1   g359(.A1(G16), .A2(G19), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n565), .B2(G16), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT90), .B(G1341), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G2072), .ZN(new_n789));
  OR2_X1    g364(.A1(G29), .A2(G33), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n487), .A2(G139), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT25), .Z(new_n793));
  AND2_X1   g368(.A1(new_n461), .A2(new_n463), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n794), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n791), .B(new_n793), .C1(new_n470), .C2(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n790), .B1(new_n796), .B2(new_n750), .ZN(new_n797));
  OAI221_X1 g372(.A(new_n788), .B1(new_n747), .B2(new_n746), .C1(new_n789), .C2(new_n797), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n783), .A2(new_n784), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n750), .A2(G26), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n489), .A2(G128), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT91), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n470), .A2(G116), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n487), .A2(G140), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n489), .A2(KEYINPUT91), .A3(G128), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n803), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n800), .B1(new_n810), .B2(new_n750), .ZN(new_n811));
  MUX2_X1   g386(.A(new_n800), .B(new_n811), .S(KEYINPUT28), .Z(new_n812));
  XOR2_X1   g387(.A(KEYINPUT92), .B(G2067), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(G168), .A2(G16), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G16), .B2(G21), .ZN(new_n816));
  INV_X1    g391(.A(G1966), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n758), .A2(G2084), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n696), .A2(G4), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n608), .B2(new_n696), .ZN(new_n820));
  INV_X1    g395(.A(G1348), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n818), .B(new_n822), .C1(new_n773), .C2(new_n774), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n789), .B2(new_n797), .ZN(new_n824));
  AND4_X1   g399(.A1(new_n775), .A2(new_n799), .A3(new_n814), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n750), .A2(G27), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G164), .B2(new_n750), .ZN(new_n827));
  INV_X1    g402(.A(G2078), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT31), .B(G11), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n743), .A2(new_n825), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n816), .A2(new_n817), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT95), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n831), .A2(new_n833), .ZN(G311));
  INV_X1    g409(.A(G311), .ZN(G150));
  XOR2_X1   g410(.A(KEYINPUT97), .B(G860), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n542), .A2(G67), .ZN(new_n837));
  NAND2_X1  g412(.A1(G80), .A2(G543), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n528), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G55), .ZN(new_n840));
  INV_X1    g415(.A(G93), .ZN(new_n841));
  OAI22_X1  g416(.A1(new_n840), .A2(new_n557), .B1(new_n532), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n836), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT37), .Z(new_n844));
  NOR2_X1   g419(.A1(new_n839), .A2(new_n842), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n564), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT39), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n608), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n847), .B(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n844), .B1(new_n850), .B2(new_n836), .ZN(G145));
  NAND2_X1  g426(.A1(new_n489), .A2(G130), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n487), .A2(G142), .ZN(new_n853));
  OR2_X1    g428(.A1(G106), .A2(G2105), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n854), .B(G2104), .C1(G118), .C2(new_n470), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n770), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n770), .A2(new_n856), .ZN(new_n858));
  OR3_X1    g433(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT98), .ZN(new_n859));
  OAI21_X1  g434(.A(KEYINPUT98), .B1(new_n857), .B2(new_n858), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n809), .B(new_n723), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n796), .B(new_n508), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n862), .A2(new_n863), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n861), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n864), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n867), .A2(new_n860), .A3(new_n859), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n638), .B(G160), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(G162), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n629), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(G37), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n872), .A2(new_n866), .A3(new_n868), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g453(.A(G290), .B(G288), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(G303), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(G305), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT42), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n883));
  OR3_X1    g458(.A1(G299), .A2(new_n883), .A3(new_n608), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n883), .B1(G299), .B2(new_n608), .ZN(new_n885));
  NAND2_X1  g460(.A1(G299), .A2(new_n608), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n884), .A2(new_n885), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n884), .A2(KEYINPUT101), .A3(new_n885), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n886), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n889), .B1(new_n894), .B2(new_n888), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n846), .B(new_n624), .Z(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n887), .B(KEYINPUT100), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n897), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n882), .B(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(G868), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(G868), .B2(new_n845), .ZN(G295));
  OAI21_X1  g477(.A(new_n901), .B1(G868), .B2(new_n845), .ZN(G331));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n880), .B(new_n707), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n906));
  NAND2_X1  g481(.A1(G171), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n846), .B(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(G286), .B1(new_n906), .B2(G171), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n908), .B(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n898), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n908), .B(new_n909), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(new_n888), .B2(new_n894), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n887), .A2(new_n888), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT104), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n905), .B(new_n913), .C1(new_n915), .C2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n911), .A2(new_n887), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n920), .B(new_n881), .C1(new_n895), .C2(new_n911), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n918), .A2(new_n919), .A3(new_n875), .A4(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n911), .A2(new_n895), .ZN(new_n923));
  INV_X1    g498(.A(new_n887), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n914), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n905), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(new_n875), .A3(new_n921), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n922), .A2(KEYINPUT103), .B1(new_n927), .B2(KEYINPUT43), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n927), .A2(KEYINPUT103), .A3(KEYINPUT43), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n904), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n927), .A2(new_n919), .ZN(new_n931));
  AND4_X1   g506(.A1(KEYINPUT43), .A2(new_n918), .A3(new_n875), .A4(new_n921), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT44), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(G397));
  XOR2_X1   g509(.A(KEYINPUT105), .B(G1384), .Z(new_n935));
  NAND2_X1  g510(.A1(new_n508), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n467), .A2(G40), .A3(new_n472), .A4(new_n476), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n769), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G1996), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n809), .B(G2067), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n945), .B2(new_n941), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n941), .A2(new_n943), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n769), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT108), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n723), .B(new_n730), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n941), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(G290), .A2(G1986), .A3(new_n941), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n941), .A2(new_n596), .A3(new_n715), .A4(new_n599), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT107), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n530), .A2(G48), .A3(G543), .A4(new_n531), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n530), .A2(G86), .A3(new_n531), .A4(new_n518), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n587), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(G1981), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT111), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n588), .A2(new_n591), .A3(new_n691), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n963), .A2(new_n967), .A3(G1981), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT49), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n940), .ZN(new_n972));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n973), .A3(new_n508), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n974), .A2(G8), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n965), .A2(new_n966), .A3(KEYINPUT49), .A4(new_n968), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n971), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G1976), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT52), .B1(G288), .B2(new_n978), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n975), .B(new_n979), .C1(new_n978), .C2(G288), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n974), .A2(G8), .ZN(new_n981));
  NOR2_X1   g556(.A1(G288), .A2(new_n978), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT52), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n977), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT113), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n977), .A2(new_n980), .A3(new_n986), .A4(new_n983), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n935), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n508), .A2(KEYINPUT109), .A3(KEYINPUT45), .A4(new_n935), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n508), .A2(new_n973), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n940), .B1(new_n994), .B2(new_n938), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n993), .A2(KEYINPUT110), .A3(new_n995), .ZN(new_n999));
  AOI21_X1  g574(.A(G1971), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n940), .B1(new_n994), .B2(KEYINPUT50), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT112), .ZN(new_n1002));
  INV_X1    g577(.A(G2090), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n508), .A2(new_n1004), .A3(new_n973), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1004), .B1(new_n508), .B2(new_n973), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1006), .B1(new_n1007), .B2(new_n940), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .A4(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(G8), .B1(new_n1000), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G303), .A2(G8), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(G2090), .ZN(new_n1018));
  OAI211_X1 g593(.A(G8), .B(new_n1014), .C1(new_n1000), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G2084), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1001), .A2(new_n1020), .A3(new_n1005), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n940), .B1(new_n994), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n508), .A2(new_n973), .A3(new_n937), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1966), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(G8), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(G286), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n988), .A2(new_n1016), .A3(new_n1019), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT63), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(G8), .B1(new_n1000), .B2(new_n1018), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n984), .B1(new_n1031), .B2(new_n1015), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1032), .A2(KEYINPUT63), .A3(new_n1019), .A4(new_n1027), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1019), .A2(new_n984), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n977), .A2(new_n978), .A3(new_n702), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n981), .B1(new_n1037), .B2(new_n966), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1034), .A2(new_n1036), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n1041));
  NOR2_X1   g616(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(G299), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1043), .B1(G299), .B2(new_n1041), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT56), .B(G2072), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n993), .A2(new_n995), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1002), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1049), .A2(new_n1050), .A3(new_n780), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n1049), .B2(new_n780), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1046), .B(new_n1048), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1017), .ZN(new_n1054));
  OAI22_X1  g629(.A1(new_n1054), .A2(G1348), .B1(G2067), .B2(new_n974), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(new_n608), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1048), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1046), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1059), .A2(KEYINPUT61), .A3(new_n1053), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1062), .B(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT60), .ZN(new_n1065));
  OR2_X1    g640(.A1(new_n1055), .A2(new_n608), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1055), .A2(new_n608), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1065), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  XOR2_X1   g644(.A(KEYINPUT58), .B(G1341), .Z(new_n1070));
  NAND2_X1  g645(.A1(new_n974), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n996), .B2(G1996), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n565), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1073), .B(new_n1074), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1055), .A2(KEYINPUT60), .A3(new_n609), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1059), .A2(new_n1053), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1069), .B(new_n1077), .C1(new_n1078), .C2(KEYINPUT61), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1061), .B1(new_n1064), .B2(new_n1079), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n985), .A2(new_n987), .ZN(new_n1081));
  INV_X1    g656(.A(G8), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n993), .A2(KEYINPUT110), .A3(new_n995), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT110), .B1(new_n993), .B2(new_n995), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n699), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1082), .B1(new_n1085), .B2(new_n1009), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1019), .B1(new_n1014), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT122), .B1(new_n1081), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n988), .A2(new_n1016), .A3(new_n1089), .A4(new_n1019), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(G286), .A2(KEYINPUT117), .A3(G8), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1026), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT117), .B1(G286), .B2(G8), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT51), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n1096));
  NAND2_X1  g671(.A1(G286), .A2(G8), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1026), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT118), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1026), .A2(new_n1100), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1095), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(G8), .B(G286), .C1(new_n1021), .C2(new_n1025), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(G171), .B(KEYINPUT54), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n972), .A2(KEYINPUT119), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n940), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(new_n939), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(G2078), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1106), .A2(KEYINPUT120), .A3(new_n939), .A4(new_n1108), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1111), .A2(new_n993), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  XOR2_X1   g690(.A(new_n1115), .B(KEYINPUT121), .Z(new_n1116));
  NOR2_X1   g691(.A1(new_n1054), .A2(G1961), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n998), .A2(new_n828), .A3(new_n999), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1117), .B1(new_n1118), .B2(new_n1112), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1105), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1023), .A2(new_n1024), .A3(new_n1113), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1121), .B1(new_n1105), .B2(new_n1123), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1091), .A2(new_n1104), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1040), .B1(new_n1080), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1104), .A2(KEYINPUT62), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT124), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1102), .A2(new_n1130), .A3(new_n1103), .ZN(new_n1131));
  AOI21_X1  g706(.A(G301), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1091), .A2(new_n1129), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1129), .B1(new_n1091), .B2(new_n1133), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1128), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n960), .B1(new_n1126), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n724), .A2(new_n731), .ZN(new_n1138));
  OAI22_X1  g713(.A1(new_n950), .A2(new_n1138), .B1(G2067), .B2(new_n809), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(new_n941), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n956), .B(KEYINPUT48), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n951), .A2(new_n953), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n945), .A2(new_n941), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n942), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1144), .B(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT47), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n947), .B(KEYINPUT46), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1147), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1140), .B(new_n1142), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT126), .B1(new_n1137), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1127), .B(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1091), .A2(new_n1133), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT123), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1091), .A2(new_n1133), .A3(new_n1129), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1154), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g733(.A(new_n1035), .B(new_n1038), .C1(new_n1030), .C2(new_n1033), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1062), .B(KEYINPUT116), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT61), .B1(new_n1059), .B2(new_n1053), .ZN(new_n1161));
  NOR4_X1   g736(.A1(new_n1161), .A2(new_n1068), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1060), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1091), .A2(new_n1104), .A3(new_n1124), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1159), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n959), .B1(new_n1158), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1151), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1152), .A2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g745(.A1(new_n657), .A2(G319), .A3(new_n673), .A4(new_n694), .ZN(new_n1172));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n1173));
  OR2_X1    g747(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g748(.A1(new_n1174), .A2(new_n877), .ZN(new_n1175));
  INV_X1    g749(.A(new_n1175), .ZN(new_n1176));
  AND2_X1   g750(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1177));
  INV_X1    g751(.A(new_n1177), .ZN(new_n1178));
  OAI211_X1 g752(.A(new_n1176), .B(new_n1178), .C1(new_n928), .C2(new_n929), .ZN(G225));
  INV_X1    g753(.A(G225), .ZN(G308));
endmodule


