

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  XNOR2_X1 U553 ( .A(KEYINPUT70), .B(n587), .ZN(n1012) );
  XOR2_X1 U554 ( .A(n767), .B(KEYINPUT32), .Z(n518) );
  BUF_X1 U555 ( .A(n984), .Z(n519) );
  XOR2_X1 U556 ( .A(KEYINPUT17), .B(n520), .Z(n984) );
  OR2_X2 U557 ( .A1(n718), .A2(n717), .ZN(n760) );
  NOR2_X1 U558 ( .A1(n778), .A2(n799), .ZN(n784) );
  NOR2_X1 U559 ( .A1(G651), .A2(n637), .ZN(n640) );
  AND2_X1 U560 ( .A1(G138), .A2(n984), .ZN(n527) );
  OR2_X1 U561 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U562 ( .A(n528), .B(KEYINPUT85), .ZN(G164) );
  INV_X1 U563 ( .A(G2104), .ZN(n521) );
  NOR2_X2 U564 ( .A1(G2105), .A2(n521), .ZN(n983) );
  NAND2_X1 U565 ( .A1(G102), .A2(n983), .ZN(n525) );
  AND2_X1 U566 ( .A1(n521), .A2(G2105), .ZN(n979) );
  NAND2_X1 U567 ( .A1(G126), .A2(n979), .ZN(n523) );
  AND2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n980) );
  NAND2_X1 U569 ( .A1(G114), .A2(n980), .ZN(n522) );
  AND2_X1 U570 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U571 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U572 ( .A(KEYINPUT72), .B(KEYINPUT7), .ZN(n542) );
  NOR2_X1 U573 ( .A1(G651), .A2(G543), .ZN(n641) );
  NAND2_X1 U574 ( .A1(n641), .A2(G89), .ZN(n529) );
  XNOR2_X1 U575 ( .A(n529), .B(KEYINPUT4), .ZN(n531) );
  XOR2_X1 U576 ( .A(KEYINPUT0), .B(G543), .Z(n637) );
  INV_X1 U577 ( .A(G651), .ZN(n533) );
  NOR2_X2 U578 ( .A1(n637), .A2(n533), .ZN(n645) );
  NAND2_X1 U579 ( .A1(G76), .A2(n645), .ZN(n530) );
  NAND2_X1 U580 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U581 ( .A(n532), .B(KEYINPUT5), .ZN(n540) );
  XNOR2_X1 U582 ( .A(KEYINPUT71), .B(KEYINPUT6), .ZN(n538) );
  NOR2_X1 U583 ( .A1(G543), .A2(n533), .ZN(n534) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n534), .Z(n642) );
  NAND2_X1 U585 ( .A1(G63), .A2(n642), .ZN(n536) );
  NAND2_X1 U586 ( .A1(G51), .A2(n640), .ZN(n535) );
  NAND2_X1 U587 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U588 ( .A(n538), .B(n537), .ZN(n539) );
  NAND2_X1 U589 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U590 ( .A(n542), .B(n541), .ZN(G168) );
  XOR2_X1 U591 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U592 ( .A1(G91), .A2(n641), .ZN(n544) );
  NAND2_X1 U593 ( .A1(G65), .A2(n642), .ZN(n543) );
  NAND2_X1 U594 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U595 ( .A1(G78), .A2(n645), .ZN(n546) );
  NAND2_X1 U596 ( .A1(G53), .A2(n640), .ZN(n545) );
  NAND2_X1 U597 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U598 ( .A1(n548), .A2(n547), .ZN(G299) );
  XOR2_X1 U599 ( .A(G2446), .B(G2451), .Z(n550) );
  XNOR2_X1 U600 ( .A(G1348), .B(G2454), .ZN(n549) );
  XNOR2_X1 U601 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U602 ( .A(n551), .B(G2435), .Z(n553) );
  XNOR2_X1 U603 ( .A(G1341), .B(G2443), .ZN(n552) );
  XNOR2_X1 U604 ( .A(n553), .B(n552), .ZN(n557) );
  XOR2_X1 U605 ( .A(KEYINPUT96), .B(G2430), .Z(n555) );
  XNOR2_X1 U606 ( .A(G2427), .B(G2438), .ZN(n554) );
  XNOR2_X1 U607 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U608 ( .A(n557), .B(n556), .Z(n558) );
  AND2_X1 U609 ( .A1(G14), .A2(n558), .ZN(G401) );
  INV_X1 U610 ( .A(G57), .ZN(G237) );
  INV_X1 U611 ( .A(G132), .ZN(G219) );
  INV_X1 U612 ( .A(G82), .ZN(G220) );
  NAND2_X1 U613 ( .A1(G64), .A2(n642), .ZN(n560) );
  NAND2_X1 U614 ( .A1(G52), .A2(n640), .ZN(n559) );
  NAND2_X1 U615 ( .A1(n560), .A2(n559), .ZN(n565) );
  NAND2_X1 U616 ( .A1(G90), .A2(n641), .ZN(n562) );
  NAND2_X1 U617 ( .A1(G77), .A2(n645), .ZN(n561) );
  NAND2_X1 U618 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U619 ( .A(KEYINPUT9), .B(n563), .Z(n564) );
  NOR2_X1 U620 ( .A1(n565), .A2(n564), .ZN(G171) );
  NAND2_X1 U621 ( .A1(G94), .A2(G452), .ZN(n566) );
  XNOR2_X1 U622 ( .A(n566), .B(KEYINPUT67), .ZN(G173) );
  NAND2_X1 U623 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U624 ( .A(n567), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U625 ( .A(G223), .ZN(n825) );
  NAND2_X1 U626 ( .A1(n825), .A2(G567), .ZN(n568) );
  XOR2_X1 U627 ( .A(KEYINPUT11), .B(n568), .Z(G234) );
  XOR2_X1 U628 ( .A(KEYINPUT68), .B(KEYINPUT14), .Z(n570) );
  NAND2_X1 U629 ( .A1(G56), .A2(n642), .ZN(n569) );
  XNOR2_X1 U630 ( .A(n570), .B(n569), .ZN(n576) );
  NAND2_X1 U631 ( .A1(n641), .A2(G81), .ZN(n571) );
  XNOR2_X1 U632 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U633 ( .A1(G68), .A2(n645), .ZN(n572) );
  NAND2_X1 U634 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT13), .B(n574), .Z(n575) );
  NOR2_X1 U636 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n640), .A2(G43), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n578), .A2(n577), .ZN(n1010) );
  INV_X1 U639 ( .A(G860), .ZN(n593) );
  OR2_X1 U640 ( .A1(n1010), .A2(n593), .ZN(G153) );
  INV_X1 U641 ( .A(G171), .ZN(G301) );
  NAND2_X1 U642 ( .A1(G54), .A2(n640), .ZN(n585) );
  NAND2_X1 U643 ( .A1(G92), .A2(n641), .ZN(n580) );
  NAND2_X1 U644 ( .A1(G66), .A2(n642), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U646 ( .A1(G79), .A2(n645), .ZN(n581) );
  XNOR2_X1 U647 ( .A(KEYINPUT69), .B(n581), .ZN(n582) );
  NOR2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(n586), .B(KEYINPUT15), .ZN(n587) );
  INV_X1 U651 ( .A(G868), .ZN(n662) );
  AND2_X1 U652 ( .A1(n1012), .A2(n662), .ZN(n589) );
  NOR2_X1 U653 ( .A1(n662), .A2(G301), .ZN(n588) );
  NOR2_X1 U654 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U655 ( .A1(G299), .A2(n662), .ZN(n591) );
  NAND2_X1 U656 ( .A1(G868), .A2(G286), .ZN(n590) );
  NAND2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U658 ( .A(KEYINPUT73), .B(n592), .Z(G297) );
  NAND2_X1 U659 ( .A1(n593), .A2(G559), .ZN(n594) );
  NAND2_X1 U660 ( .A1(n594), .A2(n1012), .ZN(n595) );
  XNOR2_X1 U661 ( .A(n595), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U662 ( .A1(G868), .A2(n1010), .ZN(n596) );
  XNOR2_X1 U663 ( .A(KEYINPUT74), .B(n596), .ZN(n599) );
  NAND2_X1 U664 ( .A1(G868), .A2(n1012), .ZN(n597) );
  NOR2_X1 U665 ( .A1(G559), .A2(n597), .ZN(n598) );
  NOR2_X1 U666 ( .A1(n599), .A2(n598), .ZN(G282) );
  NAND2_X1 U667 ( .A1(G123), .A2(n979), .ZN(n600) );
  XOR2_X1 U668 ( .A(KEYINPUT75), .B(n600), .Z(n601) );
  XNOR2_X1 U669 ( .A(n601), .B(KEYINPUT18), .ZN(n603) );
  NAND2_X1 U670 ( .A1(G111), .A2(n980), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U672 ( .A1(G99), .A2(n983), .ZN(n605) );
  NAND2_X1 U673 ( .A1(G135), .A2(n519), .ZN(n604) );
  NAND2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U675 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U676 ( .A(KEYINPUT76), .B(n608), .ZN(n1005) );
  XNOR2_X1 U677 ( .A(G2096), .B(n1005), .ZN(n610) );
  INV_X1 U678 ( .A(G2100), .ZN(n609) );
  NAND2_X1 U679 ( .A1(n610), .A2(n609), .ZN(G156) );
  NAND2_X1 U680 ( .A1(G67), .A2(n642), .ZN(n612) );
  NAND2_X1 U681 ( .A1(G55), .A2(n640), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U683 ( .A1(G93), .A2(n641), .ZN(n614) );
  NAND2_X1 U684 ( .A1(G80), .A2(n645), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U686 ( .A1(n616), .A2(n615), .ZN(n661) );
  NAND2_X1 U687 ( .A1(n1012), .A2(G559), .ZN(n617) );
  XNOR2_X1 U688 ( .A(n617), .B(n1010), .ZN(n652) );
  XOR2_X1 U689 ( .A(n652), .B(KEYINPUT77), .Z(n618) );
  NOR2_X1 U690 ( .A1(G860), .A2(n618), .ZN(n619) );
  XOR2_X1 U691 ( .A(KEYINPUT78), .B(n619), .Z(n620) );
  XOR2_X1 U692 ( .A(n661), .B(n620), .Z(G145) );
  NAND2_X1 U693 ( .A1(G88), .A2(n641), .ZN(n622) );
  NAND2_X1 U694 ( .A1(G75), .A2(n645), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U696 ( .A1(G62), .A2(n642), .ZN(n624) );
  NAND2_X1 U697 ( .A1(G50), .A2(n640), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U699 ( .A1(n626), .A2(n625), .ZN(G166) );
  NAND2_X1 U700 ( .A1(G85), .A2(n641), .ZN(n628) );
  NAND2_X1 U701 ( .A1(G72), .A2(n645), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U703 ( .A(KEYINPUT66), .B(n629), .Z(n633) );
  NAND2_X1 U704 ( .A1(G60), .A2(n642), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G47), .A2(n640), .ZN(n630) );
  AND2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n633), .A2(n632), .ZN(G290) );
  NAND2_X1 U708 ( .A1(G49), .A2(n640), .ZN(n635) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U711 ( .A1(n642), .A2(n636), .ZN(n639) );
  NAND2_X1 U712 ( .A1(n637), .A2(G87), .ZN(n638) );
  NAND2_X1 U713 ( .A1(n639), .A2(n638), .ZN(G288) );
  NAND2_X1 U714 ( .A1(n640), .A2(G48), .ZN(n650) );
  NAND2_X1 U715 ( .A1(G86), .A2(n641), .ZN(n644) );
  NAND2_X1 U716 ( .A1(G61), .A2(n642), .ZN(n643) );
  NAND2_X1 U717 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U718 ( .A1(n645), .A2(G73), .ZN(n646) );
  XOR2_X1 U719 ( .A(KEYINPUT2), .B(n646), .Z(n647) );
  NOR2_X1 U720 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U722 ( .A(KEYINPUT79), .B(n651), .Z(G305) );
  XNOR2_X1 U723 ( .A(KEYINPUT81), .B(n652), .ZN(n659) );
  XNOR2_X1 U724 ( .A(n661), .B(KEYINPUT19), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n653), .B(KEYINPUT80), .ZN(n654) );
  XNOR2_X1 U726 ( .A(G166), .B(n654), .ZN(n657) );
  XOR2_X1 U727 ( .A(G299), .B(G288), .Z(n655) );
  XNOR2_X1 U728 ( .A(G290), .B(n655), .ZN(n656) );
  XNOR2_X1 U729 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U730 ( .A(n658), .B(G305), .ZN(n1009) );
  XNOR2_X1 U731 ( .A(n659), .B(n1009), .ZN(n660) );
  NAND2_X1 U732 ( .A1(n660), .A2(G868), .ZN(n664) );
  NAND2_X1 U733 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U734 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U735 ( .A(KEYINPUT82), .B(n665), .Z(G295) );
  NAND2_X1 U736 ( .A1(G2078), .A2(G2084), .ZN(n666) );
  XOR2_X1 U737 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U738 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U739 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U740 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U741 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U742 ( .A1(G220), .A2(G219), .ZN(n670) );
  XOR2_X1 U743 ( .A(KEYINPUT22), .B(n670), .Z(n671) );
  NOR2_X1 U744 ( .A1(G218), .A2(n671), .ZN(n672) );
  XOR2_X1 U745 ( .A(KEYINPUT83), .B(n672), .Z(n673) );
  NAND2_X1 U746 ( .A1(G96), .A2(n673), .ZN(n956) );
  NAND2_X1 U747 ( .A1(G2106), .A2(n956), .ZN(n678) );
  NAND2_X1 U748 ( .A1(G120), .A2(G69), .ZN(n674) );
  NOR2_X1 U749 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U750 ( .A1(n675), .A2(G108), .ZN(n676) );
  XNOR2_X1 U751 ( .A(n676), .B(KEYINPUT84), .ZN(n957) );
  NAND2_X1 U752 ( .A1(n957), .A2(G567), .ZN(n677) );
  NAND2_X1 U753 ( .A1(n678), .A2(n677), .ZN(n1016) );
  NAND2_X1 U754 ( .A1(G483), .A2(G661), .ZN(n679) );
  NOR2_X1 U755 ( .A1(n1016), .A2(n679), .ZN(n828) );
  NAND2_X1 U756 ( .A1(n828), .A2(G36), .ZN(G176) );
  NAND2_X1 U757 ( .A1(n980), .A2(G113), .ZN(n682) );
  NAND2_X1 U758 ( .A1(G101), .A2(n983), .ZN(n680) );
  XOR2_X1 U759 ( .A(KEYINPUT23), .B(n680), .Z(n681) );
  NAND2_X1 U760 ( .A1(n682), .A2(n681), .ZN(n686) );
  NAND2_X1 U761 ( .A1(G125), .A2(n979), .ZN(n684) );
  NAND2_X1 U762 ( .A1(G137), .A2(n519), .ZN(n683) );
  NAND2_X1 U763 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U764 ( .A1(n686), .A2(n685), .ZN(G160) );
  XOR2_X1 U765 ( .A(G166), .B(KEYINPUT86), .Z(G303) );
  XNOR2_X1 U766 ( .A(G1986), .B(G290), .ZN(n930) );
  NOR2_X1 U767 ( .A1(G1384), .A2(G164), .ZN(n687) );
  XNOR2_X1 U768 ( .A(n687), .B(KEYINPUT64), .ZN(n715) );
  NAND2_X1 U769 ( .A1(G160), .A2(G40), .ZN(n717) );
  NOR2_X1 U770 ( .A1(n715), .A2(n717), .ZN(n820) );
  NAND2_X1 U771 ( .A1(n930), .A2(n820), .ZN(n807) );
  NAND2_X1 U772 ( .A1(G95), .A2(n983), .ZN(n689) );
  NAND2_X1 U773 ( .A1(G131), .A2(n519), .ZN(n688) );
  NAND2_X1 U774 ( .A1(n689), .A2(n688), .ZN(n693) );
  NAND2_X1 U775 ( .A1(G119), .A2(n979), .ZN(n691) );
  NAND2_X1 U776 ( .A1(G107), .A2(n980), .ZN(n690) );
  NAND2_X1 U777 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U778 ( .A1(n693), .A2(n692), .ZN(n999) );
  INV_X1 U779 ( .A(G1991), .ZN(n809) );
  NOR2_X1 U780 ( .A1(n999), .A2(n809), .ZN(n703) );
  XOR2_X1 U781 ( .A(KEYINPUT38), .B(KEYINPUT88), .Z(n695) );
  NAND2_X1 U782 ( .A1(G105), .A2(n983), .ZN(n694) );
  XNOR2_X1 U783 ( .A(n695), .B(n694), .ZN(n699) );
  NAND2_X1 U784 ( .A1(G129), .A2(n979), .ZN(n697) );
  NAND2_X1 U785 ( .A1(G117), .A2(n980), .ZN(n696) );
  NAND2_X1 U786 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U787 ( .A1(n699), .A2(n698), .ZN(n701) );
  NAND2_X1 U788 ( .A1(n519), .A2(G141), .ZN(n700) );
  NAND2_X1 U789 ( .A1(n701), .A2(n700), .ZN(n992) );
  AND2_X1 U790 ( .A1(n992), .A2(G1996), .ZN(n702) );
  NOR2_X1 U791 ( .A1(n703), .A2(n702), .ZN(n840) );
  INV_X1 U792 ( .A(n840), .ZN(n704) );
  NAND2_X1 U793 ( .A1(n704), .A2(n820), .ZN(n808) );
  NAND2_X1 U794 ( .A1(G104), .A2(n983), .ZN(n706) );
  NAND2_X1 U795 ( .A1(G140), .A2(n519), .ZN(n705) );
  NAND2_X1 U796 ( .A1(n706), .A2(n705), .ZN(n708) );
  XOR2_X1 U797 ( .A(KEYINPUT34), .B(KEYINPUT87), .Z(n707) );
  XNOR2_X1 U798 ( .A(n708), .B(n707), .ZN(n713) );
  NAND2_X1 U799 ( .A1(G128), .A2(n979), .ZN(n710) );
  NAND2_X1 U800 ( .A1(G116), .A2(n980), .ZN(n709) );
  NAND2_X1 U801 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U802 ( .A(KEYINPUT35), .B(n711), .Z(n712) );
  NOR2_X1 U803 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U804 ( .A(KEYINPUT36), .B(n714), .ZN(n1006) );
  XNOR2_X1 U805 ( .A(G2067), .B(KEYINPUT37), .ZN(n817) );
  NOR2_X1 U806 ( .A1(n1006), .A2(n817), .ZN(n850) );
  NAND2_X1 U807 ( .A1(n820), .A2(n850), .ZN(n815) );
  NAND2_X1 U808 ( .A1(n808), .A2(n815), .ZN(n805) );
  INV_X1 U809 ( .A(n715), .ZN(n718) );
  NOR2_X2 U810 ( .A1(n718), .A2(n717), .ZN(n744) );
  NAND2_X1 U811 ( .A1(n744), .A2(G2072), .ZN(n716) );
  XOR2_X1 U812 ( .A(KEYINPUT27), .B(n716), .Z(n720) );
  NAND2_X1 U813 ( .A1(G1956), .A2(n760), .ZN(n719) );
  NAND2_X1 U814 ( .A1(n720), .A2(n719), .ZN(n737) );
  NAND2_X1 U815 ( .A1(G299), .A2(n737), .ZN(n721) );
  XOR2_X1 U816 ( .A(KEYINPUT28), .B(n721), .Z(n742) );
  INV_X1 U817 ( .A(G2067), .ZN(n900) );
  NOR2_X2 U818 ( .A1(n760), .A2(n900), .ZN(n722) );
  XNOR2_X1 U819 ( .A(n722), .B(KEYINPUT90), .ZN(n724) );
  AND2_X1 U820 ( .A1(n760), .A2(G1348), .ZN(n723) );
  OR2_X1 U821 ( .A1(n724), .A2(n723), .ZN(n732) );
  NAND2_X1 U822 ( .A1(n744), .A2(G1996), .ZN(n726) );
  XNOR2_X1 U823 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n725) );
  XNOR2_X1 U824 ( .A(n726), .B(n725), .ZN(n730) );
  NAND2_X1 U825 ( .A1(n760), .A2(G1341), .ZN(n728) );
  INV_X1 U826 ( .A(n1010), .ZN(n727) );
  NAND2_X1 U827 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X2 U828 ( .A1(n730), .A2(n729), .ZN(n734) );
  NAND2_X1 U829 ( .A1(n734), .A2(n1012), .ZN(n731) );
  NAND2_X1 U830 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U831 ( .A(n733), .B(KEYINPUT91), .ZN(n736) );
  NOR2_X1 U832 ( .A1(n1012), .A2(n734), .ZN(n735) );
  NOR2_X1 U833 ( .A1(n736), .A2(n735), .ZN(n739) );
  NOR2_X1 U834 ( .A1(G299), .A2(n737), .ZN(n738) );
  NOR2_X1 U835 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U836 ( .A(n740), .B(KEYINPUT92), .ZN(n741) );
  NOR2_X1 U837 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U838 ( .A(n743), .B(KEYINPUT29), .ZN(n748) );
  OR2_X1 U839 ( .A1(n744), .A2(G1961), .ZN(n746) );
  XNOR2_X1 U840 ( .A(G2078), .B(KEYINPUT25), .ZN(n904) );
  NAND2_X1 U841 ( .A1(n744), .A2(n904), .ZN(n745) );
  NAND2_X1 U842 ( .A1(n746), .A2(n745), .ZN(n754) );
  NAND2_X1 U843 ( .A1(G171), .A2(n754), .ZN(n747) );
  NAND2_X1 U844 ( .A1(n748), .A2(n747), .ZN(n759) );
  NAND2_X1 U845 ( .A1(n760), .A2(G8), .ZN(n799) );
  NOR2_X1 U846 ( .A1(n799), .A2(G1966), .ZN(n749) );
  XNOR2_X1 U847 ( .A(n749), .B(KEYINPUT89), .ZN(n771) );
  INV_X1 U848 ( .A(G8), .ZN(n750) );
  NOR2_X1 U849 ( .A1(G2084), .A2(n760), .ZN(n769) );
  NOR2_X1 U850 ( .A1(n750), .A2(n769), .ZN(n751) );
  AND2_X1 U851 ( .A1(n771), .A2(n751), .ZN(n752) );
  XOR2_X1 U852 ( .A(n752), .B(KEYINPUT30), .Z(n753) );
  NOR2_X1 U853 ( .A1(G168), .A2(n753), .ZN(n756) );
  NOR2_X1 U854 ( .A1(G171), .A2(n754), .ZN(n755) );
  NOR2_X1 U855 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U856 ( .A(KEYINPUT31), .B(n757), .Z(n758) );
  NAND2_X1 U857 ( .A1(n759), .A2(n758), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n768), .A2(G286), .ZN(n765) );
  NOR2_X1 U859 ( .A1(G1971), .A2(n799), .ZN(n762) );
  NOR2_X1 U860 ( .A1(G2090), .A2(n760), .ZN(n761) );
  NOR2_X1 U861 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U862 ( .A1(n763), .A2(G303), .ZN(n764) );
  NAND2_X1 U863 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U864 ( .A1(n766), .A2(G8), .ZN(n767) );
  INV_X1 U865 ( .A(n768), .ZN(n773) );
  NAND2_X1 U866 ( .A1(G8), .A2(n769), .ZN(n770) );
  NAND2_X1 U867 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U868 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X2 U869 ( .A1(n518), .A2(n774), .ZN(n794) );
  NOR2_X1 U870 ( .A1(G303), .A2(G1971), .ZN(n775) );
  NOR2_X1 U871 ( .A1(G1976), .A2(G288), .ZN(n942) );
  NOR2_X1 U872 ( .A1(n775), .A2(n942), .ZN(n776) );
  XNOR2_X1 U873 ( .A(n776), .B(KEYINPUT93), .ZN(n777) );
  NOR2_X1 U874 ( .A1(n794), .A2(n777), .ZN(n778) );
  NAND2_X1 U875 ( .A1(G1976), .A2(G288), .ZN(n945) );
  INV_X1 U876 ( .A(KEYINPUT33), .ZN(n786) );
  INV_X1 U877 ( .A(n799), .ZN(n792) );
  NAND2_X1 U878 ( .A1(n792), .A2(n942), .ZN(n779) );
  NOR2_X1 U879 ( .A1(n786), .A2(n779), .ZN(n780) );
  XOR2_X1 U880 ( .A(n780), .B(KEYINPUT94), .Z(n785) );
  AND2_X1 U881 ( .A1(n945), .A2(n785), .ZN(n782) );
  XNOR2_X1 U882 ( .A(G1981), .B(G305), .ZN(n927) );
  INV_X1 U883 ( .A(n927), .ZN(n781) );
  AND2_X1 U884 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U885 ( .A1(n784), .A2(n783), .ZN(n790) );
  INV_X1 U886 ( .A(n785), .ZN(n787) );
  OR2_X1 U887 ( .A1(n787), .A2(n786), .ZN(n788) );
  OR2_X1 U888 ( .A1(n927), .A2(n788), .ZN(n789) );
  NAND2_X1 U889 ( .A1(n790), .A2(n789), .ZN(n803) );
  NOR2_X1 U890 ( .A1(G1981), .A2(G305), .ZN(n791) );
  XNOR2_X1 U891 ( .A(KEYINPUT24), .B(n791), .ZN(n793) );
  NAND2_X1 U892 ( .A1(n793), .A2(n792), .ZN(n801) );
  INV_X1 U893 ( .A(n794), .ZN(n797) );
  NOR2_X1 U894 ( .A1(G2090), .A2(G303), .ZN(n795) );
  NAND2_X1 U895 ( .A1(G8), .A2(n795), .ZN(n796) );
  NAND2_X1 U896 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U897 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U898 ( .A1(n801), .A2(n800), .ZN(n802) );
  NOR2_X1 U899 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U900 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n823) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n992), .ZN(n843) );
  INV_X1 U903 ( .A(n808), .ZN(n812) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n810) );
  AND2_X1 U905 ( .A1(n809), .A2(n999), .ZN(n839) );
  NOR2_X1 U906 ( .A1(n810), .A2(n839), .ZN(n811) );
  NOR2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U908 ( .A1(n843), .A2(n813), .ZN(n814) );
  XNOR2_X1 U909 ( .A(n814), .B(KEYINPUT39), .ZN(n816) );
  NAND2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n1006), .A2(n817), .ZN(n852) );
  NAND2_X1 U912 ( .A1(n818), .A2(n852), .ZN(n819) );
  XOR2_X1 U913 ( .A(KEYINPUT95), .B(n819), .Z(n821) );
  NAND2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U916 ( .A(n824), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U917 ( .A1(n825), .A2(G2106), .ZN(n826) );
  XOR2_X1 U918 ( .A(KEYINPUT97), .B(n826), .Z(G217) );
  AND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U920 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G1), .A2(G3), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U923 ( .A(n830), .B(KEYINPUT98), .ZN(G188) );
  XNOR2_X1 U924 ( .A(G69), .B(KEYINPUT99), .ZN(G235) );
  NAND2_X1 U926 ( .A1(G124), .A2(n979), .ZN(n831) );
  XOR2_X1 U927 ( .A(KEYINPUT105), .B(n831), .Z(n832) );
  XNOR2_X1 U928 ( .A(n832), .B(KEYINPUT44), .ZN(n834) );
  NAND2_X1 U929 ( .A1(G112), .A2(n980), .ZN(n833) );
  NAND2_X1 U930 ( .A1(n834), .A2(n833), .ZN(n838) );
  NAND2_X1 U931 ( .A1(G100), .A2(n983), .ZN(n836) );
  NAND2_X1 U932 ( .A1(G136), .A2(n519), .ZN(n835) );
  NAND2_X1 U933 ( .A1(n836), .A2(n835), .ZN(n837) );
  NOR2_X1 U934 ( .A1(n838), .A2(n837), .ZN(G162) );
  XNOR2_X1 U935 ( .A(KEYINPUT55), .B(KEYINPUT112), .ZN(n918) );
  NOR2_X1 U936 ( .A1(n839), .A2(n1005), .ZN(n848) );
  XNOR2_X1 U937 ( .A(G160), .B(G2084), .ZN(n841) );
  NAND2_X1 U938 ( .A1(n841), .A2(n840), .ZN(n846) );
  XOR2_X1 U939 ( .A(G2090), .B(G162), .Z(n842) );
  NOR2_X1 U940 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U941 ( .A(n844), .B(KEYINPUT51), .ZN(n845) );
  NOR2_X1 U942 ( .A1(n846), .A2(n845), .ZN(n847) );
  NAND2_X1 U943 ( .A1(n848), .A2(n847), .ZN(n849) );
  NOR2_X1 U944 ( .A1(n850), .A2(n849), .ZN(n851) );
  XNOR2_X1 U945 ( .A(n851), .B(KEYINPUT110), .ZN(n853) );
  NAND2_X1 U946 ( .A1(n853), .A2(n852), .ZN(n854) );
  XOR2_X1 U947 ( .A(KEYINPUT111), .B(n854), .Z(n867) );
  NAND2_X1 U948 ( .A1(G103), .A2(n983), .ZN(n856) );
  NAND2_X1 U949 ( .A1(G139), .A2(n519), .ZN(n855) );
  NAND2_X1 U950 ( .A1(n856), .A2(n855), .ZN(n862) );
  NAND2_X1 U951 ( .A1(G127), .A2(n979), .ZN(n858) );
  NAND2_X1 U952 ( .A1(G115), .A2(n980), .ZN(n857) );
  NAND2_X1 U953 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U954 ( .A(KEYINPUT107), .B(n859), .ZN(n860) );
  XNOR2_X1 U955 ( .A(KEYINPUT47), .B(n860), .ZN(n861) );
  NOR2_X1 U956 ( .A1(n862), .A2(n861), .ZN(n991) );
  XOR2_X1 U957 ( .A(G2072), .B(n991), .Z(n864) );
  XOR2_X1 U958 ( .A(G164), .B(G2078), .Z(n863) );
  NOR2_X1 U959 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U960 ( .A(KEYINPUT50), .B(n865), .Z(n866) );
  NOR2_X1 U961 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U962 ( .A(KEYINPUT52), .B(n868), .Z(n869) );
  NOR2_X1 U963 ( .A1(n918), .A2(n869), .ZN(n870) );
  XNOR2_X1 U964 ( .A(KEYINPUT113), .B(n870), .ZN(n871) );
  NAND2_X1 U965 ( .A1(n871), .A2(G29), .ZN(n925) );
  XNOR2_X1 U966 ( .A(G1986), .B(G24), .ZN(n877) );
  XNOR2_X1 U967 ( .A(G1971), .B(G22), .ZN(n872) );
  XNOR2_X1 U968 ( .A(n872), .B(KEYINPUT124), .ZN(n874) );
  XNOR2_X1 U969 ( .A(G23), .B(G1976), .ZN(n873) );
  NOR2_X1 U970 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U971 ( .A(KEYINPUT125), .B(n875), .ZN(n876) );
  NOR2_X1 U972 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U973 ( .A(KEYINPUT126), .B(n878), .ZN(n879) );
  XNOR2_X1 U974 ( .A(n879), .B(KEYINPUT58), .ZN(n893) );
  XOR2_X1 U975 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n889) );
  XNOR2_X1 U976 ( .A(G1956), .B(G20), .ZN(n881) );
  XNOR2_X1 U977 ( .A(G6), .B(G1981), .ZN(n880) );
  NOR2_X1 U978 ( .A1(n881), .A2(n880), .ZN(n887) );
  XOR2_X1 U979 ( .A(G4), .B(KEYINPUT122), .Z(n883) );
  XNOR2_X1 U980 ( .A(G1348), .B(KEYINPUT59), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n885) );
  XNOR2_X1 U982 ( .A(G1341), .B(G19), .ZN(n884) );
  NOR2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n886) );
  NAND2_X1 U984 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U985 ( .A(n889), .B(n888), .ZN(n891) );
  XNOR2_X1 U986 ( .A(G21), .B(G1966), .ZN(n890) );
  NOR2_X1 U987 ( .A1(n891), .A2(n890), .ZN(n892) );
  NAND2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n895) );
  XNOR2_X1 U989 ( .A(G5), .B(G1961), .ZN(n894) );
  NOR2_X1 U990 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U991 ( .A(KEYINPUT61), .B(n896), .Z(n897) );
  NOR2_X1 U992 ( .A1(G16), .A2(n897), .ZN(n923) );
  XOR2_X1 U993 ( .A(KEYINPUT115), .B(G34), .Z(n899) );
  XNOR2_X1 U994 ( .A(G2084), .B(KEYINPUT54), .ZN(n898) );
  XNOR2_X1 U995 ( .A(n899), .B(n898), .ZN(n916) );
  XOR2_X1 U996 ( .A(G2090), .B(G35), .Z(n914) );
  XNOR2_X1 U997 ( .A(G26), .B(n900), .ZN(n901) );
  NAND2_X1 U998 ( .A1(n901), .A2(G28), .ZN(n910) );
  XNOR2_X1 U999 ( .A(G1996), .B(G32), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(G33), .B(G2072), .ZN(n902) );
  NOR2_X1 U1001 ( .A1(n903), .A2(n902), .ZN(n908) );
  XOR2_X1 U1002 ( .A(n904), .B(G27), .Z(n906) );
  XNOR2_X1 U1003 ( .A(G1991), .B(G25), .ZN(n905) );
  NOR2_X1 U1004 ( .A1(n906), .A2(n905), .ZN(n907) );
  NAND2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1007 ( .A(KEYINPUT53), .B(n911), .Z(n912) );
  XNOR2_X1 U1008 ( .A(n912), .B(KEYINPUT114), .ZN(n913) );
  NAND2_X1 U1009 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1011 ( .A(n918), .B(n917), .ZN(n920) );
  INV_X1 U1012 ( .A(G29), .ZN(n919) );
  NAND2_X1 U1013 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1014 ( .A1(n921), .A2(G11), .ZN(n922) );
  NOR2_X1 U1015 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1016 ( .A1(n925), .A2(n924), .ZN(n954) );
  XOR2_X1 U1017 ( .A(KEYINPUT56), .B(G16), .Z(n952) );
  XOR2_X1 U1018 ( .A(G168), .B(G1966), .Z(n926) );
  NOR2_X1 U1019 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1020 ( .A(KEYINPUT57), .B(n928), .Z(n941) );
  XNOR2_X1 U1021 ( .A(G1956), .B(G299), .ZN(n929) );
  NOR2_X1 U1022 ( .A1(n930), .A2(n929), .ZN(n932) );
  XOR2_X1 U1023 ( .A(G1341), .B(n1010), .Z(n931) );
  NAND2_X1 U1024 ( .A1(n932), .A2(n931), .ZN(n939) );
  XNOR2_X1 U1025 ( .A(G171), .B(G1961), .ZN(n933) );
  XNOR2_X1 U1026 ( .A(n933), .B(KEYINPUT117), .ZN(n936) );
  XOR2_X1 U1027 ( .A(G1348), .B(KEYINPUT116), .Z(n934) );
  XNOR2_X1 U1028 ( .A(n1012), .B(n934), .ZN(n935) );
  NOR2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1030 ( .A(KEYINPUT118), .B(n937), .Z(n938) );
  NOR2_X1 U1031 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1032 ( .A1(n941), .A2(n940), .ZN(n949) );
  XOR2_X1 U1033 ( .A(n942), .B(KEYINPUT119), .Z(n944) );
  XNOR2_X1 U1034 ( .A(G303), .B(G1971), .ZN(n943) );
  NOR2_X1 U1035 ( .A1(n944), .A2(n943), .ZN(n946) );
  NAND2_X1 U1036 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1037 ( .A(KEYINPUT120), .B(n947), .ZN(n948) );
  NOR2_X1 U1038 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1039 ( .A(KEYINPUT121), .B(n950), .Z(n951) );
  NOR2_X1 U1040 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1041 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1042 ( .A(n955), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1043 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1044 ( .A(G120), .ZN(G236) );
  INV_X1 U1045 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1046 ( .A1(n957), .A2(n956), .ZN(G325) );
  INV_X1 U1047 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1048 ( .A(G1966), .B(G2474), .ZN(n967) );
  XOR2_X1 U1049 ( .A(KEYINPUT104), .B(G1986), .Z(n959) );
  XNOR2_X1 U1050 ( .A(G1971), .B(G1981), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(n959), .B(n958), .ZN(n963) );
  XOR2_X1 U1052 ( .A(KEYINPUT41), .B(G1991), .Z(n961) );
  XNOR2_X1 U1053 ( .A(G1996), .B(G1976), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(n961), .B(n960), .ZN(n962) );
  XOR2_X1 U1055 ( .A(n963), .B(n962), .Z(n965) );
  XNOR2_X1 U1056 ( .A(G1961), .B(G1956), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(n965), .B(n964), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(n967), .B(n966), .ZN(G229) );
  XNOR2_X1 U1059 ( .A(G2078), .B(G2072), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(n968), .B(G2100), .ZN(n978) );
  XOR2_X1 U1061 ( .A(KEYINPUT42), .B(G2678), .Z(n970) );
  XNOR2_X1 U1062 ( .A(KEYINPUT43), .B(KEYINPUT103), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(n970), .B(n969), .ZN(n974) );
  XOR2_X1 U1064 ( .A(KEYINPUT102), .B(G2096), .Z(n972) );
  XNOR2_X1 U1065 ( .A(G2090), .B(KEYINPUT101), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(n972), .B(n971), .ZN(n973) );
  XOR2_X1 U1067 ( .A(n974), .B(n973), .Z(n976) );
  XNOR2_X1 U1068 ( .A(G2067), .B(G2084), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(n976), .B(n975), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(n978), .B(n977), .ZN(G227) );
  NAND2_X1 U1071 ( .A1(G130), .A2(n979), .ZN(n982) );
  NAND2_X1 U1072 ( .A1(G118), .A2(n980), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n990) );
  NAND2_X1 U1074 ( .A1(G106), .A2(n983), .ZN(n986) );
  NAND2_X1 U1075 ( .A1(G142), .A2(n519), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1077 ( .A(KEYINPUT45), .B(n987), .Z(n988) );
  XNOR2_X1 U1078 ( .A(KEYINPUT106), .B(n988), .ZN(n989) );
  NOR2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n1003) );
  XOR2_X1 U1080 ( .A(G162), .B(n991), .Z(n994) );
  XOR2_X1 U1081 ( .A(G160), .B(n992), .Z(n993) );
  XNOR2_X1 U1082 ( .A(n994), .B(n993), .ZN(n998) );
  XOR2_X1 U1083 ( .A(KEYINPUT46), .B(KEYINPUT108), .Z(n996) );
  XNOR2_X1 U1084 ( .A(KEYINPUT109), .B(KEYINPUT48), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(n996), .B(n995), .ZN(n997) );
  XOR2_X1 U1086 ( .A(n998), .B(n997), .Z(n1001) );
  XNOR2_X1 U1087 ( .A(G164), .B(n999), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(n1001), .B(n1000), .ZN(n1002) );
  XOR2_X1 U1089 ( .A(n1003), .B(n1002), .Z(n1004) );
  XNOR2_X1 U1090 ( .A(n1005), .B(n1004), .ZN(n1007) );
  XOR2_X1 U1091 ( .A(n1007), .B(n1006), .Z(n1008) );
  NOR2_X1 U1092 ( .A1(G37), .A2(n1008), .ZN(G395) );
  XNOR2_X1 U1093 ( .A(n1009), .B(G301), .ZN(n1011) );
  XNOR2_X1 U1094 ( .A(n1011), .B(n1010), .ZN(n1013) );
  XNOR2_X1 U1095 ( .A(n1013), .B(n1012), .ZN(n1014) );
  XNOR2_X1 U1096 ( .A(n1014), .B(G286), .ZN(n1015) );
  NOR2_X1 U1097 ( .A1(G37), .A2(n1015), .ZN(G397) );
  XOR2_X1 U1098 ( .A(KEYINPUT100), .B(n1016), .Z(G319) );
  NOR2_X1 U1099 ( .A1(G229), .A2(G227), .ZN(n1017) );
  XNOR2_X1 U1100 ( .A(KEYINPUT49), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1101 ( .A1(G401), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1102 ( .A1(G395), .A2(G397), .ZN(n1019) );
  AND2_X1 U1103 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1104 ( .A1(n1021), .A2(G319), .ZN(G225) );
  INV_X1 U1105 ( .A(G225), .ZN(G308) );
  INV_X1 U1106 ( .A(G108), .ZN(G238) );
endmodule

