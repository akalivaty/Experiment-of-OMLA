//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1307, new_n1308, new_n1309,
    new_n1310, new_n1311, new_n1312, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT65), .B(G20), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(new_n201), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G50), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI22_X1  g0029(.A1(new_n226), .A2(new_n229), .B1(new_n210), .B2(new_n211), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n217), .B1(new_n221), .B2(new_n223), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT66), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G244), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G1), .A3(G13), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(G274), .ZN(new_n254));
  OAI22_X1  g0054(.A1(new_n249), .A2(new_n253), .B1(new_n254), .B2(new_n252), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(G232), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(G238), .A3(G1698), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n258), .B(new_n259), .C1(new_n207), .C2(new_n256), .ZN(new_n260));
  AND2_X1   g0060(.A1(G1), .A2(G13), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT68), .ZN(new_n262));
  AND3_X1   g0062(.A1(new_n261), .A2(new_n262), .A3(new_n250), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n262), .B1(new_n261), .B2(new_n250), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n255), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G200), .ZN(new_n268));
  NAND3_X1  g0068(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n219), .ZN(new_n270));
  INV_X1    g0070(.A(G77), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT8), .B(G58), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  OAI22_X1  g0074(.A1(new_n271), .A2(new_n218), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT65), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G20), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(new_n278), .A3(G33), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT15), .B(G87), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n270), .B1(new_n275), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G77), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n270), .B1(new_n210), .B2(G20), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(G77), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT70), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n282), .A2(KEYINPUT70), .A3(new_n286), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n266), .A2(G190), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n268), .A2(new_n289), .A3(new_n290), .A4(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n260), .A2(new_n265), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  INV_X1    g0094(.A(new_n255), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT71), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT71), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n266), .A2(new_n298), .A3(new_n294), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n289), .A2(new_n290), .ZN(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n267), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n292), .B1(new_n300), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT72), .ZN(new_n306));
  INV_X1    g0106(.A(new_n270), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(G1), .B2(new_n211), .ZN(new_n308));
  INV_X1    g0108(.A(G58), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT8), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT8), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G58), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT69), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n272), .A2(KEYINPUT69), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n308), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n313), .A2(new_n314), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n272), .A2(KEYINPUT69), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n283), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT7), .ZN(new_n324));
  AND2_X1   g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  NOR2_X1   g0125(.A1(KEYINPUT3), .A2(G33), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n324), .B1(new_n327), .B2(new_n218), .ZN(new_n328));
  NOR4_X1   g0128(.A1(new_n325), .A2(new_n326), .A3(KEYINPUT7), .A4(G20), .ZN(new_n329));
  INV_X1    g0129(.A(G68), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AND2_X1   g0131(.A1(G58), .A2(G68), .ZN(new_n332));
  OAI21_X1  g0132(.A(G20), .B1(new_n332), .B2(new_n201), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n273), .A2(G159), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n323), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT3), .ZN(new_n337));
  INV_X1    g0137(.A(G33), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(KEYINPUT3), .A2(G33), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(new_n211), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n330), .B1(new_n341), .B2(KEYINPUT7), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n327), .A2(new_n218), .A3(new_n324), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n335), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n307), .B1(new_n344), .B2(KEYINPUT16), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n321), .B1(new_n336), .B2(new_n345), .ZN(new_n346));
  OAI211_X1 g0146(.A(G223), .B(new_n257), .C1(new_n325), .C2(new_n326), .ZN(new_n347));
  OAI211_X1 g0147(.A(G226), .B(G1698), .C1(new_n325), .C2(new_n326), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G87), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n265), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n251), .A2(new_n252), .ZN(new_n352));
  INV_X1    g0152(.A(new_n252), .ZN(new_n353));
  INV_X1    g0153(.A(G274), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n261), .B2(new_n250), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n352), .A2(G232), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n351), .A2(G179), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n302), .B1(new_n351), .B2(new_n356), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR3_X1   g0159(.A1(new_n346), .A2(new_n359), .A3(KEYINPUT18), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT18), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n317), .A2(new_n320), .ZN(new_n362));
  INV_X1    g0162(.A(new_n335), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n325), .A2(new_n326), .A3(G20), .ZN(new_n364));
  OAI21_X1  g0164(.A(G68), .B1(new_n364), .B2(new_n324), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n327), .A2(new_n218), .A3(new_n324), .ZN(new_n366));
  OAI211_X1 g0166(.A(KEYINPUT16), .B(new_n363), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n270), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n276), .A2(new_n278), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT7), .B1(new_n369), .B2(new_n256), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n327), .A2(new_n324), .A3(new_n211), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(G68), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n322), .B1(new_n372), .B2(new_n363), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n362), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n351), .A2(G179), .A3(new_n356), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n351), .A2(new_n356), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(new_n302), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n361), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n360), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(G200), .B1(new_n351), .B2(new_n356), .ZN(new_n380));
  INV_X1    g0180(.A(G190), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n380), .B1(new_n381), .B2(new_n376), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT17), .B1(new_n374), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n351), .A2(new_n381), .A3(new_n356), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n376), .B2(G200), .ZN(new_n385));
  XOR2_X1   g0185(.A(KEYINPUT74), .B(KEYINPUT17), .Z(new_n386));
  NAND3_X1  g0186(.A1(new_n346), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT72), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n389), .B(new_n292), .C1(new_n300), .C2(new_n304), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n306), .A2(new_n379), .A3(new_n388), .A4(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n283), .A2(G50), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n285), .B2(G50), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n315), .A2(new_n316), .A3(G33), .A4(new_n218), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n273), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT9), .B(new_n393), .C1(new_n396), .C2(new_n307), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT9), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n307), .B1(new_n394), .B2(new_n395), .ZN(new_n399));
  INV_X1    g0199(.A(new_n393), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n254), .A2(new_n252), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(G226), .B2(new_n352), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n265), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n256), .A2(G222), .A3(new_n257), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n256), .A2(G223), .A3(G1698), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n327), .A2(G77), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n405), .B1(new_n409), .B2(KEYINPUT67), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT67), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n406), .A2(new_n407), .A3(new_n411), .A4(new_n408), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n404), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G200), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n397), .B(new_n401), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n410), .A2(new_n412), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n403), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(new_n381), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT10), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n397), .A2(new_n401), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n417), .A2(G200), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT10), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n413), .A2(G190), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n420), .A2(new_n421), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n413), .A2(new_n294), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n393), .B1(new_n396), .B2(new_n307), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n426), .B(new_n427), .C1(G169), .C2(new_n413), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n273), .A2(G50), .B1(G20), .B2(new_n330), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n279), .B2(new_n271), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n431), .A2(new_n270), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n432), .A2(KEYINPUT11), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(KEYINPUT11), .ZN(new_n434));
  OR3_X1    g0234(.A1(new_n283), .A2(KEYINPUT12), .A3(G68), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT12), .B1(new_n283), .B2(G68), .ZN(new_n436));
  AOI22_X1  g0236(.A1(G68), .A2(new_n285), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n433), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n256), .A2(G232), .A3(G1698), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n256), .A2(G226), .A3(new_n257), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G97), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n265), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n402), .B1(G238), .B2(new_n352), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT13), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n446), .B1(new_n444), .B2(new_n445), .ZN(new_n448));
  OAI21_X1  g0248(.A(G169), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n444), .A2(new_n445), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT13), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI22_X1  g0253(.A1(new_n449), .A2(KEYINPUT14), .B1(new_n453), .B2(new_n294), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT14), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(new_n453), .B2(G169), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n439), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n453), .A2(G200), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n451), .A2(G190), .A3(new_n452), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n438), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n391), .A2(new_n429), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G45), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(G1), .ZN(new_n465));
  AND2_X1   g0265(.A1(KEYINPUT5), .A2(G41), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(G264), .A3(new_n251), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT83), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT83), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n468), .A2(new_n471), .A3(G264), .A4(new_n251), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(G250), .B(new_n257), .C1(new_n325), .C2(new_n326), .ZN(new_n474));
  OAI211_X1 g0274(.A(G257), .B(G1698), .C1(new_n325), .C2(new_n326), .ZN(new_n475));
  XOR2_X1   g0275(.A(KEYINPUT82), .B(G294), .Z(new_n476));
  OAI211_X1 g0276(.A(new_n474), .B(new_n475), .C1(new_n476), .C2(new_n338), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n265), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n254), .A2(new_n468), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n473), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n414), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n478), .A2(new_n381), .A3(new_n480), .A4(new_n469), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT23), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n369), .A2(new_n485), .A3(new_n207), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT80), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G116), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n487), .B1(new_n488), .B2(G20), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n211), .A2(KEYINPUT80), .A3(G33), .A4(G116), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n486), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n276), .B(new_n278), .C1(new_n325), .C2(new_n326), .ZN(new_n494));
  INV_X1    g0294(.A(G87), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT22), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT22), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n218), .A2(new_n256), .A3(new_n497), .A4(G87), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT24), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n493), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n500), .B1(new_n493), .B2(new_n499), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n270), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n283), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT25), .B1(new_n504), .B2(new_n207), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(KEYINPUT25), .A3(new_n207), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n210), .A2(G33), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n283), .A2(new_n508), .A3(new_n219), .A4(new_n269), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n506), .A2(new_n507), .B1(new_n510), .B2(G107), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n484), .A2(new_n503), .A3(new_n511), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n328), .A2(new_n329), .A3(new_n207), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n207), .A2(KEYINPUT6), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n206), .A2(KEYINPUT75), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT75), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G97), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n514), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G97), .A2(G107), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT6), .B1(new_n208), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n369), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n274), .A2(new_n271), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n270), .B1(new_n513), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n283), .A2(G97), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(new_n510), .B2(G97), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT77), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT6), .ZN(new_n529));
  AND2_X1   g0329(.A1(G97), .A2(G107), .ZN(new_n530));
  NOR2_X1   g0330(.A1(G97), .A2(G107), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g0332(.A(KEYINPUT75), .B(G97), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n532), .B1(new_n533), .B2(new_n514), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n522), .B1(new_n534), .B2(new_n369), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n370), .A2(G107), .A3(new_n371), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n307), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT77), .ZN(new_n538));
  INV_X1    g0338(.A(new_n527), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n468), .A2(G257), .A3(new_n251), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT76), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT76), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n468), .A2(new_n543), .A3(G257), .A4(new_n251), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n479), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(G244), .B(new_n257), .C1(new_n325), .C2(new_n326), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT4), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n256), .A2(KEYINPUT4), .A3(G244), .A4(new_n257), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G283), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n256), .A2(G250), .A3(G1698), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n548), .A2(new_n549), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n265), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n545), .A2(new_n553), .A3(G179), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n302), .B1(new_n545), .B2(new_n553), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n528), .A2(new_n540), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n280), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(new_n283), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT19), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n279), .B2(new_n533), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n276), .B(new_n278), .C1(new_n559), .C2(new_n442), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n515), .A2(new_n517), .A3(new_n495), .A4(new_n207), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n218), .A2(new_n256), .A3(G68), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n560), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n558), .B1(new_n565), .B2(new_n270), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n510), .A2(G87), .ZN(new_n567));
  OAI211_X1 g0367(.A(G244), .B(G1698), .C1(new_n325), .C2(new_n326), .ZN(new_n568));
  OAI211_X1 g0368(.A(G238), .B(new_n257), .C1(new_n325), .C2(new_n326), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n569), .A3(new_n488), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n265), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n355), .A2(new_n465), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n210), .A2(G45), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n251), .A2(G250), .A3(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n571), .A2(new_n575), .A3(G190), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n566), .A2(new_n567), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n571), .A2(new_n575), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G200), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n571), .A2(new_n575), .A3(new_n294), .ZN(new_n580));
  AOI21_X1  g0380(.A(G169), .B1(new_n571), .B2(new_n575), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n510), .A2(new_n557), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n566), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n577), .A2(new_n579), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n545), .A2(new_n553), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G200), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n537), .A2(new_n539), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n587), .B(new_n588), .C1(new_n381), .C2(new_n586), .ZN(new_n589));
  AND4_X1   g0389(.A1(new_n512), .A2(new_n556), .A3(new_n585), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n493), .A2(new_n499), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT24), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n493), .A2(new_n499), .A3(new_n500), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n307), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n511), .ZN(new_n595));
  OAI21_X1  g0395(.A(KEYINPUT81), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n478), .A2(new_n480), .A3(new_n469), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n597), .A2(new_n302), .B1(new_n481), .B2(new_n294), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT81), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n503), .A2(new_n599), .A3(new_n511), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n596), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(G257), .B(new_n257), .C1(new_n325), .C2(new_n326), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT78), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n327), .A2(G303), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n256), .A2(G264), .A3(G1698), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n602), .A2(new_n603), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n265), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n468), .A2(new_n251), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n479), .B1(new_n610), .B2(G270), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n302), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(G116), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n504), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n509), .B2(new_n613), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n269), .A2(new_n219), .B1(G20), .B2(new_n613), .ZN(new_n616));
  AOI21_X1  g0416(.A(G33), .B1(new_n515), .B2(new_n517), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n276), .A2(new_n278), .A3(new_n550), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT20), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(KEYINPUT20), .B(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n615), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n623), .A2(KEYINPUT79), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT79), .ZN(new_n625));
  AOI211_X1 g0425(.A(new_n625), .B(new_n615), .C1(new_n621), .C2(new_n622), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n612), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT21), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n609), .A2(G179), .A3(new_n611), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n624), .B2(new_n626), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n612), .B(KEYINPUT21), .C1(new_n624), .C2(new_n626), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n624), .A2(new_n626), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n609), .A2(new_n611), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(G200), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n609), .A2(G190), .A3(new_n611), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n590), .A2(new_n601), .A3(new_n633), .A4(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n463), .A2(new_n639), .ZN(G372));
  OAI21_X1  g0440(.A(KEYINPUT18), .B1(new_n346), .B2(new_n359), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n374), .A2(new_n361), .A3(new_n377), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n641), .A2(KEYINPUT84), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT84), .B1(new_n641), .B2(new_n642), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n460), .ZN(new_n646));
  INV_X1    g0446(.A(new_n304), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n297), .A2(new_n299), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n457), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n645), .B1(new_n650), .B2(new_n388), .ZN(new_n651));
  INV_X1    g0451(.A(new_n425), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n428), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n586), .A2(G169), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n545), .A2(new_n553), .A3(G179), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n588), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n582), .A2(new_n584), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n579), .A2(new_n566), .A3(new_n567), .A4(new_n576), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n657), .A2(new_n658), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n659), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n538), .B1(new_n537), .B2(new_n539), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n525), .A2(KEYINPUT77), .A3(new_n527), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n663), .A2(new_n664), .B1(new_n655), .B2(new_n656), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n658), .B1(new_n665), .B2(new_n585), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n598), .B1(new_n594), .B2(new_n595), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n629), .A2(new_n668), .A3(new_n631), .A4(new_n632), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n512), .A2(new_n585), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n556), .A2(new_n589), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n654), .B1(new_n463), .B2(new_n674), .ZN(G369));
  NAND3_X1  g0475(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n218), .A2(new_n210), .A3(G13), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  OR3_X1    g0483(.A1(new_n676), .A2(new_n634), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n638), .ZN(new_n685));
  OAI22_X1  g0485(.A1(new_n676), .A2(new_n685), .B1(new_n634), .B2(new_n683), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G330), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n596), .A2(new_n600), .A3(new_n682), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n601), .A2(new_n690), .A3(new_n512), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT85), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n601), .A2(new_n690), .A3(KEYINPUT85), .A4(new_n512), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n596), .A2(new_n598), .A3(new_n600), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n682), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n689), .A2(new_n698), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n668), .A2(new_n682), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n633), .A2(new_n682), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n693), .A2(new_n694), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n699), .A2(new_n700), .A3(new_n702), .ZN(G399));
  NOR2_X1   g0503(.A1(new_n214), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G1), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n533), .A2(new_n495), .A3(new_n207), .A4(new_n613), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n706), .A2(new_n707), .B1(new_n223), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n696), .A2(new_n676), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n512), .A2(new_n556), .A3(new_n585), .A4(new_n589), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n685), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n710), .A2(new_n712), .A3(new_n683), .ZN(new_n713));
  INV_X1    g0513(.A(new_n586), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n572), .A2(new_n574), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n570), .B2(new_n265), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n716), .A2(new_n473), .A3(new_n478), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n630), .A2(new_n714), .A3(new_n717), .A4(KEYINPUT30), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n470), .A2(new_n472), .B1(new_n477), .B2(new_n265), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n720), .A2(new_n545), .A3(new_n553), .A4(new_n716), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n609), .A2(G179), .A3(new_n611), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n716), .A2(G179), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n635), .A2(new_n724), .A3(new_n586), .A4(new_n481), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n718), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n726), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT31), .B1(new_n726), .B2(new_n682), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n688), .B1(new_n713), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n632), .A2(new_n631), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n601), .A2(new_n732), .A3(new_n629), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n556), .A2(new_n589), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT87), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT87), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n556), .A2(new_n736), .A3(new_n589), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n733), .A2(new_n670), .A3(new_n735), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n659), .A2(new_n660), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n556), .A2(new_n739), .A3(KEYINPUT26), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n659), .B(KEYINPUT86), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n658), .B1(new_n585), .B2(new_n657), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(KEYINPUT88), .A3(KEYINPUT29), .A4(new_n683), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT29), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n746), .B(new_n682), .C1(new_n738), .C2(new_n743), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT88), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n682), .B1(new_n667), .B2(new_n672), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n748), .B1(new_n749), .B2(KEYINPUT29), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n731), .B(new_n745), .C1(new_n747), .C2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n709), .B1(new_n752), .B2(G1), .ZN(G364));
  NOR2_X1   g0553(.A1(new_n369), .A2(new_n213), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n706), .B1(G45), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n219), .B1(G20), .B2(new_n302), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n214), .A2(new_n327), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT89), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G355), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(G116), .B2(new_n215), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n214), .A2(new_n256), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G45), .B2(new_n223), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(G45), .B2(new_n247), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n760), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n414), .A2(G179), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(G20), .A3(G190), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n495), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n381), .A2(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n369), .B1(new_n773), .B2(G179), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n327), .B(new_n771), .C1(G97), .C2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n369), .A2(G179), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n414), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n381), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n775), .B1(new_n330), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT90), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n776), .A2(G190), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n776), .A2(new_n773), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n782), .A2(new_n271), .B1(new_n784), .B2(new_n309), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n779), .B1(new_n780), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(KEYINPUT92), .B1(new_n218), .B2(G190), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT92), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n369), .A2(new_n788), .A3(new_n381), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n790), .A2(G179), .A3(new_n414), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n207), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n786), .B(new_n794), .C1(new_n780), .C2(new_n785), .ZN(new_n795));
  AND3_X1   g0595(.A1(new_n777), .A2(KEYINPUT91), .A3(G190), .ZN(new_n796));
  AOI21_X1  g0596(.A(KEYINPUT91), .B1(new_n777), .B2(G190), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n795), .B1(G50), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT93), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n294), .A2(new_n414), .ZN(new_n802));
  OR3_X1    g0602(.A1(new_n790), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n801), .B1(new_n790), .B2(new_n802), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G159), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT32), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n805), .B(KEYINPUT94), .Z(new_n809));
  INV_X1    g0609(.A(G329), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G311), .ZN(new_n812));
  INV_X1    g0612(.A(G322), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n782), .A2(new_n812), .B1(new_n784), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G303), .ZN(new_n815));
  INV_X1    g0615(.A(new_n774), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n327), .B1(new_n815), .B2(new_n770), .C1(new_n816), .C2(new_n476), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G283), .ZN(new_n819));
  XOR2_X1   g0619(.A(KEYINPUT33), .B(G317), .Z(new_n820));
  OAI221_X1 g0620(.A(new_n818), .B1(new_n819), .B2(new_n792), .C1(new_n778), .C2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G326), .B2(new_n799), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n800), .A2(new_n808), .B1(new_n811), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n759), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n755), .B(new_n768), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n687), .B2(new_n758), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT95), .Z(new_n827));
  INV_X1    g0627(.A(new_n689), .ZN(new_n828));
  INV_X1    g0628(.A(new_n755), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n687), .A2(new_n688), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G396));
  NAND4_X1  g0634(.A1(new_n648), .A2(new_n303), .A3(new_n301), .A4(new_n682), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT98), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT98), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n647), .A2(new_n837), .A3(new_n648), .A4(new_n682), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n301), .A2(new_n682), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n649), .A2(new_n292), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n749), .B(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n755), .B1(new_n843), .B2(new_n731), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n731), .B2(new_n843), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n824), .A2(new_n757), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n755), .B1(G77), .B2(new_n846), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n781), .A2(G159), .B1(new_n783), .B2(G143), .ZN(new_n848));
  INV_X1    g0648(.A(G150), .ZN(new_n849));
  INV_X1    g0649(.A(G137), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n848), .B1(new_n849), .B2(new_n778), .C1(new_n798), .C2(new_n850), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT34), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n791), .A2(G68), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n202), .B2(new_n770), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT97), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n854), .A2(KEYINPUT97), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n327), .B1(new_n774), .B2(G58), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n852), .A2(new_n855), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G132), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n809), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n809), .A2(new_n812), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n792), .A2(new_n495), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT96), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n783), .A2(G294), .B1(G97), .B2(new_n774), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n770), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n256), .B1(new_n866), .B2(G107), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n867), .B1(new_n778), .B2(new_n819), .C1(new_n613), .C2(new_n782), .ZN(new_n868));
  INV_X1    g0668(.A(new_n864), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(KEYINPUT96), .B2(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n865), .B(new_n870), .C1(new_n815), .C2(new_n798), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n858), .A2(new_n860), .B1(new_n861), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n847), .B1(new_n872), .B2(new_n759), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n757), .B2(new_n842), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n845), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(G384));
  OAI21_X1  g0676(.A(new_n745), .B1(new_n747), .B2(new_n750), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n462), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n654), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT103), .Z(new_n880));
  NAND2_X1  g0680(.A1(new_n645), .A2(new_n680), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n711), .B1(new_n633), .B2(new_n668), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT26), .B1(new_n556), .B2(new_n739), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(new_n659), .A3(new_n661), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n842), .B(new_n683), .C1(new_n882), .C2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n649), .A2(new_n682), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n457), .B(new_n460), .C1(new_n438), .C2(new_n683), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n449), .A2(KEYINPUT14), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n453), .A2(new_n455), .A3(G169), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n890), .B(new_n891), .C1(new_n294), .C2(new_n453), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n439), .B(new_n682), .C1(new_n646), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n346), .A2(new_n385), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n374), .A2(new_n377), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n346), .A2(new_n680), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(KEYINPUT37), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n344), .A2(new_n322), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n362), .B1(new_n368), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n680), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n903), .A2(new_n377), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n897), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n899), .A2(new_n901), .B1(new_n907), .B2(KEYINPUT37), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n905), .B1(new_n379), .B2(new_n388), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n896), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n905), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n346), .A2(new_n385), .A3(new_n386), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT17), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n346), .B2(new_n385), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n641), .A2(new_n642), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n907), .A2(KEYINPUT37), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n374), .A2(new_n904), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT37), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n898), .A2(new_n897), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n917), .A2(new_n922), .A3(KEYINPUT38), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n910), .A2(KEYINPUT100), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT100), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n925), .B(new_n896), .C1(new_n908), .C2(new_n909), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n881), .B1(new_n895), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n892), .A2(new_n439), .A3(new_n683), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n924), .A2(KEYINPUT39), .A3(new_n926), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n920), .B1(new_n919), .B2(KEYINPUT101), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n899), .A2(new_n932), .A3(new_n919), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT101), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT37), .B1(new_n900), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n898), .A2(new_n897), .A3(new_n919), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT102), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n912), .B2(new_n914), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n383), .A2(KEYINPUT102), .A3(new_n387), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n940), .B(new_n941), .C1(new_n643), .C2(new_n644), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n938), .B1(new_n942), .B2(new_n900), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n931), .B(new_n923), .C1(new_n943), .C2(KEYINPUT38), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n929), .B1(new_n930), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n928), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n880), .B(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT40), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n670), .A2(new_n671), .A3(new_n638), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n950), .A2(new_n733), .A3(new_n682), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n727), .A2(new_n728), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n842), .B(new_n894), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n949), .B1(new_n927), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n923), .B1(new_n943), .B2(KEYINPUT38), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n713), .A2(new_n729), .B1(new_n841), .B2(new_n839), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n955), .A2(KEYINPUT40), .A3(new_n894), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n729), .B1(new_n639), .B2(new_n682), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n462), .A2(new_n959), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n958), .A2(new_n960), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n961), .A2(new_n962), .A3(new_n688), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n948), .A2(new_n963), .B1(new_n210), .B2(new_n754), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n948), .B2(new_n963), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n223), .A2(new_n271), .A3(new_n332), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n202), .A2(G68), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n210), .B(G13), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n534), .A2(KEYINPUT35), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n534), .A2(KEYINPUT35), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n969), .A2(G116), .A3(new_n220), .A4(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(KEYINPUT99), .B(KEYINPUT36), .Z(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  OR3_X1    g0773(.A1(new_n965), .A2(new_n968), .A3(new_n973), .ZN(G367));
  OAI21_X1  g0774(.A(new_n682), .B1(new_n537), .B2(new_n539), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n735), .A2(new_n737), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n657), .A2(new_n682), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n979), .A2(new_n702), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT42), .Z(new_n981));
  OAI21_X1  g0781(.A(new_n556), .B1(new_n979), .B2(new_n601), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n981), .B1(new_n683), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n566), .A2(new_n567), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n682), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n585), .A2(new_n985), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n659), .A2(new_n985), .ZN(new_n987));
  XNOR2_X1  g0787(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n983), .A2(new_n986), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n986), .A2(new_n987), .ZN(new_n990));
  MUX2_X1   g0790(.A(new_n988), .B(KEYINPUT43), .S(new_n990), .Z(new_n991));
  OAI21_X1  g0791(.A(new_n989), .B1(new_n983), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n699), .A2(new_n979), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n992), .B(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n754), .A2(G45), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(G1), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT107), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n704), .B(KEYINPUT41), .Z(new_n999));
  NAND3_X1  g0799(.A1(new_n702), .A2(new_n700), .A3(new_n978), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT45), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n702), .A2(new_n700), .ZN(new_n1004));
  AOI21_X1  g0804(.A(KEYINPUT44), .B1(new_n1004), .B2(new_n979), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT44), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1006), .B(new_n978), .C1(new_n702), .C2(new_n700), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n1002), .A2(new_n1003), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n699), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n699), .B1(new_n1005), .B2(new_n1007), .C1(new_n1003), .C2(new_n1002), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n695), .B(new_n697), .C1(new_n633), .C2(new_n682), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n702), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n689), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n828), .A2(new_n1012), .A3(new_n702), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n751), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1010), .A2(new_n1011), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(KEYINPUT105), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT105), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1010), .A2(new_n1011), .A3(new_n1019), .A4(new_n1016), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n999), .B1(new_n1021), .B2(new_n752), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n998), .B1(new_n1022), .B2(KEYINPUT106), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT106), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1024), .B(new_n999), .C1(new_n1021), .C2(new_n752), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n994), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n765), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n760), .B1(new_n215), .B2(new_n280), .C1(new_n236), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT108), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1030), .A2(new_n1031), .A3(new_n829), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n758), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n792), .A2(new_n533), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n770), .A2(new_n613), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n256), .B1(new_n1035), .B2(KEYINPUT46), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(KEYINPUT46), .B2(new_n1035), .C1(new_n778), .C2(new_n476), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n782), .A2(new_n819), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n784), .A2(new_n815), .B1(new_n816), .B2(new_n207), .ZN(new_n1039));
  NOR4_X1   g0839(.A1(new_n1034), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(G317), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1040), .B1(new_n812), .B2(new_n798), .C1(new_n1041), .C2(new_n805), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n784), .A2(new_n849), .B1(new_n816), .B2(new_n330), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n799), .B2(G143), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(KEYINPUT109), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n327), .B1(new_n866), .B2(G58), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n778), .B2(new_n806), .C1(new_n202), .C2(new_n782), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(G77), .B2(new_n791), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1045), .B(new_n1048), .C1(new_n850), .C2(new_n805), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1044), .A2(KEYINPUT109), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1042), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT47), .Z(new_n1052));
  OAI221_X1 g0852(.A(new_n1032), .B1(new_n1033), .B2(new_n990), .C1(new_n1052), .C2(new_n824), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1026), .A2(new_n1053), .ZN(G387));
  XNOR2_X1  g0854(.A(new_n707), .B(KEYINPUT110), .ZN(new_n1055));
  OR3_X1    g0855(.A1(new_n272), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1056));
  OAI21_X1  g0856(.A(KEYINPUT50), .B1(new_n272), .B2(G50), .ZN(new_n1057));
  AOI21_X1  g0857(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n765), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1060), .A2(KEYINPUT111), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(KEYINPUT111), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(new_n464), .C2(new_n240), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n762), .A2(new_n707), .B1(new_n207), .B2(new_n214), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n829), .B1(new_n1065), .B2(new_n760), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT112), .Z(new_n1067));
  INV_X1    g0867(.A(new_n805), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(G150), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n866), .A2(G77), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n256), .B(new_n1070), .C1(new_n782), .C2(new_n330), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n816), .A2(new_n280), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G50), .B2(new_n783), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1074), .A2(KEYINPUT113), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n318), .A2(new_n319), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n778), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1071), .B(new_n1075), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n799), .A2(G159), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1074), .A2(KEYINPUT113), .B1(G97), .B2(new_n791), .ZN(new_n1080));
  AND4_X1   g0880(.A1(new_n1069), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n781), .A2(G303), .B1(new_n783), .B2(G317), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n812), .B2(new_n778), .C1(new_n798), .C2(new_n813), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT48), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n476), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(G283), .A2(new_n774), .B1(new_n1087), .B2(new_n866), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1085), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1090), .A2(KEYINPUT49), .ZN(new_n1091));
  INV_X1    g0891(.A(G326), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n327), .B1(new_n613), .B2(new_n792), .C1(new_n805), .C2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n1090), .B2(KEYINPUT49), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1081), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1067), .B1(new_n1095), .B2(new_n824), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n698), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(new_n1097), .B2(new_n758), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(new_n1099), .B2(new_n997), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n752), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n704), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1099), .A2(new_n752), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1100), .B1(new_n1102), .B2(new_n1103), .ZN(G393));
  NAND2_X1  g0904(.A1(new_n244), .A2(new_n765), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1105), .B(new_n760), .C1(new_n215), .C2(new_n533), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT114), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n829), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n1107), .B2(new_n1106), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n327), .B1(new_n866), .B2(G68), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1110), .B1(new_n816), .B2(new_n271), .C1(new_n782), .C2(new_n272), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1111), .B(new_n862), .C1(G50), .C2(new_n1077), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n798), .A2(new_n849), .B1(new_n806), .B2(new_n784), .ZN(new_n1113));
  XOR2_X1   g0913(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1068), .A2(G143), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1112), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n256), .B(new_n793), .C1(G283), .C2(new_n866), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n781), .A2(G294), .B1(G116), .B2(new_n774), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n815), .B2(new_n778), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT116), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1121), .B(new_n1124), .C1(new_n813), .C2(new_n805), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n798), .A2(new_n1041), .B1(new_n812), .B2(new_n784), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT52), .Z(new_n1127));
  NOR2_X1   g0927(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1120), .B1(new_n1129), .B2(KEYINPUT117), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(KEYINPUT117), .B2(new_n1129), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1109), .B1(new_n1131), .B2(new_n759), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n1033), .B2(new_n978), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1133), .B1(new_n1134), .B2(new_n998), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n705), .B1(new_n1134), .B2(new_n1101), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1135), .B1(new_n1021), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(G390));
  AOI21_X1  g0938(.A(new_n682), .B1(new_n738), .B2(new_n743), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n886), .B1(new_n1139), .B2(new_n842), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n889), .A2(new_n893), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n929), .B(new_n955), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1141), .B1(new_n885), .B2(new_n887), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n929), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n930), .B(new_n944), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n730), .A2(new_n842), .A3(new_n894), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1142), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1146), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n959), .A2(G330), .A3(new_n842), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n1141), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n1152), .A2(new_n1146), .A3(new_n1140), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1152), .A2(new_n1146), .B1(new_n885), .B2(new_n887), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n462), .A2(new_n959), .A3(G330), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n878), .A2(new_n654), .A3(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n705), .B1(new_n1150), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n730), .A2(new_n842), .A3(new_n894), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n1147), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1156), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n653), .B(new_n1164), .C1(new_n877), .C2(new_n462), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n894), .B1(new_n730), .B2(new_n842), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n888), .B1(new_n1161), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1152), .A2(new_n1146), .A3(new_n1140), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1163), .A2(KEYINPUT118), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(KEYINPUT118), .B1(new_n1163), .B2(new_n1170), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1159), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n755), .B1(new_n1076), .B2(new_n846), .ZN(new_n1174));
  XOR2_X1   g0974(.A(KEYINPUT54), .B(G143), .Z(new_n1175));
  AOI22_X1  g0975(.A1(new_n781), .A2(new_n1175), .B1(G159), .B2(new_n774), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n850), .B2(new_n778), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT119), .Z(new_n1178));
  NOR2_X1   g0978(.A1(new_n770), .A2(new_n849), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT53), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n327), .B1(new_n783), .B2(G132), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(new_n792), .C2(new_n202), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G128), .B2(new_n799), .ZN(new_n1183));
  INV_X1    g0983(.A(G125), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1178), .B(new_n1183), .C1(new_n809), .C2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(G294), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n853), .B1(new_n809), .B2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT120), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n256), .B(new_n771), .C1(G77), .C2(new_n774), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n533), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n781), .A2(new_n1190), .B1(new_n783), .B2(G116), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n207), .B2(new_n778), .C1(new_n819), .C2(new_n798), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1185), .B1(new_n1188), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT121), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n824), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1174), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n930), .A2(new_n944), .A3(new_n756), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT122), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1198), .A2(KEYINPUT122), .A3(new_n1199), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1150), .A2(new_n997), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1173), .A2(new_n1204), .ZN(G378));
  INV_X1    g1005(.A(KEYINPUT125), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n427), .A2(new_n904), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n429), .A2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n429), .A2(new_n1207), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  OR3_X1    g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1211), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n924), .A2(new_n926), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n959), .A2(new_n842), .A3(new_n894), .ZN(new_n1217));
  AOI21_X1  g1017(.A(KEYINPUT40), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n923), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n942), .A2(new_n900), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n938), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1219), .B1(new_n1222), .B2(new_n896), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n959), .A2(KEYINPUT40), .A3(new_n842), .A4(new_n894), .ZN(new_n1224));
  OAI21_X1  g1024(.A(G330), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1215), .B1(new_n1218), .B2(new_n1225), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n954), .A2(new_n1214), .A3(new_n957), .A4(G330), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1226), .A2(new_n946), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n946), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1206), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1224), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n688), .B1(new_n1231), .B2(new_n955), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1214), .B1(new_n1232), .B2(new_n954), .ZN(new_n1233));
  AND4_X1   g1033(.A1(G330), .A2(new_n954), .A3(new_n957), .A4(new_n1214), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n947), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1226), .A2(new_n946), .A3(new_n1227), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(KEYINPUT125), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1230), .A2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1165), .B1(new_n1163), .B2(new_n1170), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT57), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1239), .A2(new_n1241), .A3(KEYINPUT57), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n704), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1240), .A2(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1214), .A2(new_n757), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n755), .B1(G50), .B2(new_n846), .ZN(new_n1246));
  INV_X1    g1046(.A(G41), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n791), .A2(G58), .ZN(new_n1248));
  AND4_X1   g1048(.A1(new_n1247), .A2(new_n1248), .A3(new_n327), .A4(new_n1070), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n809), .B2(new_n819), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT124), .Z(new_n1251));
  AOI22_X1  g1051(.A1(new_n781), .A2(new_n557), .B1(G68), .B2(new_n774), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n207), .B2(new_n784), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G97), .B2(new_n1077), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1251), .B(new_n1254), .C1(new_n613), .C2(new_n798), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT58), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(G33), .A2(G41), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT123), .ZN(new_n1260));
  AOI211_X1 g1060(.A(G50), .B(new_n1260), .C1(new_n1247), .C2(new_n327), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n774), .A2(G150), .B1(new_n866), .B2(new_n1175), .ZN(new_n1262));
  INV_X1    g1062(.A(G128), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n1262), .B1(new_n784), .B2(new_n1263), .C1(new_n782), .C2(new_n850), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(G132), .B2(new_n1077), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1184), .B2(new_n798), .ZN(new_n1266));
  OR2_X1    g1066(.A1(new_n1266), .A2(KEYINPUT59), .ZN(new_n1267));
  INV_X1    g1067(.A(G124), .ZN(new_n1268));
  OAI221_X1 g1068(.A(new_n1260), .B1(new_n806), .B2(new_n792), .C1(new_n805), .C2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n1266), .B2(KEYINPUT59), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1261), .B1(new_n1267), .B2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1257), .A2(new_n1258), .A3(new_n1271), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n1245), .B(new_n1246), .C1(new_n1272), .C2(new_n759), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n1238), .B2(new_n997), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1244), .A2(new_n1274), .ZN(G375));
  NAND2_X1  g1075(.A1(new_n1169), .A2(new_n997), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n755), .B1(G68), .B2(new_n846), .ZN(new_n1277));
  AOI211_X1 g1077(.A(new_n256), .B(new_n1072), .C1(G97), .C2(new_n866), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n781), .A2(G107), .B1(new_n783), .B2(G283), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1278), .B(new_n1279), .C1(new_n613), .C2(new_n778), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(G77), .B2(new_n791), .ZN(new_n1281));
  OAI221_X1 g1081(.A(new_n1281), .B1(new_n1186), .B2(new_n798), .C1(new_n815), .C2(new_n809), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1077), .A2(new_n1175), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n256), .B1(new_n770), .B2(new_n806), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1284), .B1(G50), .B2(new_n774), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n781), .A2(G150), .B1(new_n783), .B2(G137), .ZN(new_n1286));
  AND4_X1   g1086(.A1(new_n1248), .A2(new_n1283), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1287));
  OAI221_X1 g1087(.A(new_n1287), .B1(new_n859), .B2(new_n798), .C1(new_n809), .C2(new_n1263), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1282), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1277), .B1(new_n1289), .B2(new_n759), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1290), .B1(new_n757), .B2(new_n894), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1276), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n999), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1294), .A2(new_n1170), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1293), .A2(new_n1296), .ZN(G381));
  INV_X1    g1097(.A(new_n1204), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT118), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n1150), .B2(new_n1158), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1163), .A2(KEYINPUT118), .A3(new_n1170), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1298), .B1(new_n1302), .B2(new_n1159), .ZN(new_n1303));
  NOR4_X1   g1103(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n1304), .A3(new_n1137), .ZN(new_n1305));
  OR3_X1    g1105(.A1(G387), .A2(G375), .A3(new_n1305), .ZN(G407));
  NAND4_X1  g1106(.A1(new_n1244), .A2(new_n681), .A3(new_n1303), .A4(new_n1274), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1307), .A2(G213), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(G407), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(KEYINPUT126), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT126), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(G407), .A2(new_n1311), .A3(new_n1308), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(G409));
  OAI211_X1 g1113(.A(G378), .B(new_n1274), .C1(new_n1240), .C2(new_n1243), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1228), .A2(new_n1229), .A3(new_n1206), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT125), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1295), .B(new_n1239), .C1(new_n1315), .C2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1273), .B1(new_n1241), .B2(new_n997), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1303), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1314), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n681), .A2(G213), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT60), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1324), .B1(new_n1294), .B2(new_n1170), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1324), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n704), .ZN(new_n1327));
  NOR3_X1   g1127(.A1(new_n1325), .A2(new_n1327), .A3(KEYINPUT127), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT127), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1330));
  OAI21_X1  g1130(.A(KEYINPUT60), .B1(new_n1158), .B2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n705), .B1(new_n1294), .B2(new_n1324), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1329), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1293), .B1(new_n1328), .B2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n875), .ZN(new_n1335));
  OAI21_X1  g1135(.A(KEYINPUT127), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1331), .A2(new_n1329), .A3(new_n1332), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1338), .A2(G384), .A3(new_n1293), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n681), .A2(G213), .A3(G2897), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1335), .A2(new_n1339), .A3(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1340), .ZN(new_n1342));
  AOI21_X1  g1142(.A(G384), .B1(new_n1338), .B2(new_n1293), .ZN(new_n1343));
  AOI211_X1 g1143(.A(new_n875), .B(new_n1292), .C1(new_n1336), .C2(new_n1337), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1342), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1323), .A2(new_n1341), .A3(new_n1345), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1321), .A2(new_n1347), .A3(new_n1322), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(KEYINPUT62), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT61), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT62), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1321), .A2(new_n1347), .A3(new_n1351), .A4(new_n1322), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1346), .A2(new_n1349), .A3(new_n1350), .A4(new_n1352), .ZN(new_n1353));
  XNOR2_X1  g1153(.A(G393), .B(new_n833), .ZN(new_n1354));
  XNOR2_X1  g1154(.A(new_n1354), .B(new_n1137), .ZN(new_n1355));
  AND3_X1   g1155(.A1(new_n1026), .A2(new_n1053), .A3(new_n1355), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1355), .B1(new_n1026), .B2(new_n1053), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1353), .A2(new_n1359), .ZN(new_n1360));
  AND2_X1   g1160(.A1(new_n1345), .A2(new_n1341), .ZN(new_n1361));
  AOI21_X1  g1161(.A(KEYINPUT61), .B1(new_n1361), .B2(new_n1323), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT63), .ZN(new_n1363));
  OR2_X1    g1163(.A1(new_n1348), .A2(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1348), .A2(new_n1363), .ZN(new_n1365));
  NAND4_X1  g1165(.A1(new_n1362), .A2(new_n1364), .A3(new_n1358), .A4(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1360), .A2(new_n1366), .ZN(G405));
  OAI21_X1  g1167(.A(new_n1347), .B1(new_n1356), .B2(new_n1357), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1355), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(G387), .A2(new_n1369), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1026), .A2(new_n1355), .A3(new_n1053), .ZN(new_n1371));
  INV_X1    g1171(.A(new_n1347), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1370), .A2(new_n1371), .A3(new_n1372), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1368), .A2(new_n1373), .ZN(new_n1374));
  AOI21_X1  g1174(.A(G378), .B1(new_n1244), .B2(new_n1274), .ZN(new_n1375));
  INV_X1    g1175(.A(new_n1314), .ZN(new_n1376));
  NOR2_X1   g1176(.A1(new_n1375), .A2(new_n1376), .ZN(new_n1377));
  INV_X1    g1177(.A(new_n1377), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1374), .A2(new_n1378), .ZN(new_n1379));
  NAND3_X1  g1179(.A1(new_n1368), .A2(new_n1373), .A3(new_n1377), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1379), .A2(new_n1380), .ZN(G402));
endmodule


