//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G131), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  AOI21_X1  g004(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n187), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT17), .ZN(new_n193));
  INV_X1    g007(.A(G237), .ZN(new_n194));
  INV_X1    g008(.A(G953), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G214), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G131), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT64), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G131), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n198), .A2(new_n203), .A3(new_n189), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n192), .A2(new_n193), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n198), .A2(new_n189), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT17), .A3(new_n187), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT79), .A2(G125), .ZN(new_n209));
  INV_X1    g023(.A(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(KEYINPUT79), .A2(G125), .A3(G140), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT80), .ZN(new_n214));
  INV_X1    g028(.A(G125), .ZN(new_n215));
  NOR3_X1   g029(.A1(new_n215), .A2(KEYINPUT16), .A3(G140), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n213), .A2(KEYINPUT16), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n210), .A2(G125), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT80), .B1(new_n218), .B2(KEYINPUT16), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n217), .A2(KEYINPUT81), .A3(G146), .A4(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n212), .ZN(new_n221));
  AOI21_X1  g035(.A(G140), .B1(KEYINPUT79), .B2(G125), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT16), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n216), .A2(new_n214), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n223), .A2(G146), .A3(new_n224), .A4(new_n219), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT81), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n220), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT82), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n223), .A2(new_n219), .A3(new_n224), .ZN(new_n230));
  INV_X1    g044(.A(G146), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(new_n229), .A3(new_n231), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n208), .B(new_n228), .C1(new_n232), .C2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n206), .A2(KEYINPUT18), .A3(G131), .ZN(new_n236));
  XNOR2_X1  g050(.A(G125), .B(G140), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n231), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n238), .B1(new_n213), .B2(new_n231), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT18), .A2(G131), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n198), .A2(new_n189), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n236), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(G113), .B(G122), .ZN(new_n243));
  INV_X1    g057(.A(G104), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n245), .B(KEYINPUT94), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n235), .A2(new_n242), .A3(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n237), .A2(KEYINPUT19), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT19), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(new_n211), .B2(new_n212), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n231), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT93), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n192), .A2(new_n204), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n225), .A3(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n252), .A2(new_n253), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n242), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n245), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(G475), .B1(new_n248), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G902), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n261), .A2(KEYINPUT20), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT20), .B1(new_n261), .B2(new_n262), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n248), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n245), .B1(new_n235), .B2(new_n242), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n262), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT95), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI211_X1 g084(.A(KEYINPUT95), .B(new_n262), .C1(new_n266), .C2(new_n267), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(G475), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n197), .A2(G128), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT13), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G128), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G143), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n273), .A2(new_n274), .ZN(new_n279));
  OAI21_X1  g093(.A(G134), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G134), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n273), .A2(new_n277), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(G116), .B(G122), .ZN(new_n283));
  INV_X1    g097(.A(G107), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n283), .A2(new_n284), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n280), .B(new_n282), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G116), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT14), .B1(new_n288), .B2(G122), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n283), .B1(KEYINPUT14), .B2(new_n284), .ZN(new_n291));
  INV_X1    g105(.A(new_n282), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n281), .B1(new_n273), .B2(new_n277), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n290), .B(new_n291), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  XOR2_X1   g109(.A(KEYINPUT75), .B(G217), .Z(new_n296));
  XOR2_X1   g110(.A(KEYINPUT9), .B(G234), .Z(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(new_n195), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n295), .B(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n262), .ZN(new_n300));
  INV_X1    g114(.A(G478), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n301), .A2(KEYINPUT15), .ZN(new_n302));
  XOR2_X1   g116(.A(new_n300), .B(new_n302), .Z(new_n303));
  AND3_X1   g117(.A1(new_n265), .A2(new_n272), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT87), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n195), .A2(G227), .ZN(new_n306));
  XOR2_X1   g120(.A(new_n306), .B(KEYINPUT83), .Z(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(G110), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(new_n210), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT11), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n310), .B1(new_n281), .B2(G137), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n281), .A2(G137), .ZN(new_n312));
  INV_X1    g126(.A(G137), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT11), .A3(G134), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G131), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n203), .A2(new_n312), .A3(new_n311), .A4(new_n314), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT86), .B1(new_n284), .B2(G104), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT86), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n244), .A3(G107), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n284), .A2(G104), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G101), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n244), .B2(G107), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n284), .A2(KEYINPUT3), .A3(G104), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G101), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n244), .A2(G107), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n324), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n276), .A2(KEYINPUT1), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n231), .A2(G143), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n197), .A2(G146), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n197), .A2(KEYINPUT1), .A3(G146), .ZN(new_n337));
  XNOR2_X1  g151(.A(G143), .B(G146), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n336), .B(new_n337), .C1(G128), .C2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n331), .A3(new_n324), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n318), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT12), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n343), .B(new_n344), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n284), .A2(KEYINPUT3), .A3(G104), .ZN(new_n346));
  AOI21_X1  g160(.A(KEYINPUT3), .B1(new_n284), .B2(G104), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n330), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G101), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(KEYINPUT4), .A3(new_n331), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT0), .A4(G128), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT0), .B(G128), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n351), .B1(new_n338), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT67), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n351), .B(KEYINPUT67), .C1(new_n338), .C2(new_n352), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n350), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT84), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n329), .B1(new_n328), .B2(new_n330), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n326), .A2(new_n327), .B1(new_n244), .B2(G107), .ZN(new_n362));
  NOR4_X1   g176(.A1(new_n362), .A2(KEYINPUT84), .A3(KEYINPUT4), .A4(new_n329), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT85), .B1(new_n357), .B2(new_n364), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n355), .A2(new_n356), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n348), .A2(new_n360), .A3(G101), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT84), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n359), .A2(new_n358), .A3(new_n360), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n366), .A2(new_n370), .A3(new_n371), .A4(new_n350), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n365), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n318), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n341), .B(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n373), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n345), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n373), .A2(new_n377), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n318), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n376), .B1(new_n365), .B2(new_n372), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n309), .B1(new_n382), .B2(new_n374), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n309), .A2(new_n379), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n305), .B(G469), .C1(new_n384), .C2(G902), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n382), .A2(new_n374), .ZN(new_n386));
  AOI211_X1 g200(.A(new_n318), .B(new_n376), .C1(new_n365), .C2(new_n372), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n309), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n383), .A2(new_n345), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G469), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT88), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(KEYINPUT88), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n390), .A2(new_n262), .A3(new_n392), .A4(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n381), .A2(new_n383), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n343), .B(KEYINPUT12), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n309), .B1(new_n387), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(new_n398), .A3(G469), .ZN(new_n399));
  NAND2_X1  g213(.A1(G469), .A2(G902), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(KEYINPUT87), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n385), .A2(new_n395), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n297), .A2(new_n262), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n403), .A2(G221), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G952), .ZN(new_n406));
  AOI211_X1 g220(.A(G953), .B(new_n406), .C1(G234), .C2(G237), .ZN(new_n407));
  INV_X1    g221(.A(G234), .ZN(new_n408));
  OAI211_X1 g222(.A(G902), .B(G953), .C1(new_n408), .C2(new_n194), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n409), .B(KEYINPUT96), .Z(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT21), .B(G898), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n407), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G214), .B1(G237), .B2(G902), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT66), .ZN(new_n416));
  OR2_X1    g230(.A1(KEYINPUT2), .A2(G113), .ZN(new_n417));
  NAND2_X1  g231(.A1(KEYINPUT2), .A2(G113), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G119), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G116), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n288), .A2(G119), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n416), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G116), .B(G119), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n425), .A2(KEYINPUT66), .A3(new_n417), .A4(new_n418), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n421), .A2(new_n422), .B1(new_n417), .B2(new_n418), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n430), .B(new_n350), .C1(new_n361), .C2(new_n363), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n288), .A2(KEYINPUT5), .A3(G119), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n432), .B1(new_n425), .B2(KEYINPUT5), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n424), .A2(new_n426), .B1(new_n433), .B2(G113), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n434), .A2(new_n332), .A3(KEYINPUT89), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT89), .B1(new_n434), .B2(new_n332), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n431), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XOR2_X1   g251(.A(G110), .B(G122), .Z(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n438), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n431), .B(new_n440), .C1(new_n435), .C2(new_n436), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(KEYINPUT6), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n437), .A2(new_n443), .A3(new_n438), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n445));
  AOI21_X1  g259(.A(G128), .B1(new_n334), .B2(new_n335), .ZN(new_n446));
  INV_X1    g260(.A(new_n337), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n215), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n353), .A2(G125), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n195), .A2(G224), .ZN(new_n452));
  XOR2_X1   g266(.A(new_n451), .B(new_n452), .Z(new_n453));
  NAND3_X1  g267(.A1(new_n442), .A2(new_n444), .A3(new_n453), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n449), .A2(KEYINPUT90), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n449), .A2(KEYINPUT90), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n450), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n452), .A2(KEYINPUT7), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n451), .A2(new_n458), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n457), .A2(new_n458), .B1(KEYINPUT91), .B2(new_n459), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n438), .B(KEYINPUT8), .Z(new_n461));
  AND2_X1   g275(.A1(new_n434), .A2(new_n332), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n434), .A2(new_n332), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n459), .A2(KEYINPUT91), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n460), .A2(new_n464), .A3(new_n441), .A4(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n454), .A2(new_n262), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(G210), .B1(G237), .B2(G902), .ZN(new_n468));
  XOR2_X1   g282(.A(new_n468), .B(KEYINPUT92), .Z(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n454), .A2(new_n262), .A3(new_n468), .A4(new_n466), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n415), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND4_X1   g286(.A1(new_n304), .A2(new_n402), .A3(new_n405), .A4(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n313), .A2(G134), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n281), .A2(G137), .ZN(new_n475));
  OAI21_X1  g289(.A(G131), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n315), .B2(new_n187), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT68), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n317), .A2(KEYINPUT68), .A3(new_n476), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(new_n339), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n355), .A2(new_n318), .A3(new_n356), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT69), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n483), .B1(new_n427), .B2(new_n429), .ZN(new_n484));
  AOI211_X1 g298(.A(KEYINPUT69), .B(new_n428), .C1(new_n424), .C2(new_n426), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n481), .B(new_n482), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT73), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT28), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n487), .B1(new_n486), .B2(new_n488), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT26), .B(G101), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n188), .A2(G210), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT65), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n497), .B1(new_n448), .B2(new_n477), .ZN(new_n498));
  INV_X1    g312(.A(new_n353), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n318), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n339), .A2(KEYINPUT65), .A3(new_n317), .A4(new_n476), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n502), .A2(new_n430), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n430), .A2(KEYINPUT69), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n427), .A2(new_n483), .A3(new_n429), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n506), .A2(KEYINPUT70), .A3(new_n482), .A4(new_n481), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT70), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n486), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n503), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n491), .B(new_n496), .C1(new_n488), .C2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT29), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n507), .A2(new_n509), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n502), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n481), .A2(KEYINPUT30), .A3(new_n482), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n516), .A3(new_n430), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n496), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n511), .A2(new_n512), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT74), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n481), .A2(new_n482), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n504), .A3(new_n505), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n488), .B1(new_n513), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n490), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n519), .A2(new_n512), .ZN(new_n531));
  AOI21_X1  g345(.A(G902), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n511), .A2(KEYINPUT74), .A3(new_n512), .A4(new_n520), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n523), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G472), .ZN(new_n535));
  NOR2_X1   g349(.A1(G472), .A2(G902), .ZN(new_n536));
  INV_X1    g350(.A(new_n503), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n488), .B1(new_n513), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n519), .B1(new_n538), .B2(new_n529), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n513), .A2(new_n517), .A3(new_n496), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT31), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n513), .A2(new_n517), .A3(new_n496), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT72), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT72), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n513), .A2(new_n546), .A3(new_n517), .A4(new_n496), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n541), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n536), .B1(new_n543), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT32), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT32), .B(new_n536), .C1(new_n543), .C2(new_n548), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n535), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n296), .B1(new_n408), .B2(G902), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n228), .B1(new_n234), .B2(new_n232), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT23), .B1(new_n276), .B2(G119), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT77), .B1(new_n276), .B2(G119), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n557), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n560), .A2(KEYINPUT78), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(KEYINPUT78), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(G110), .A3(new_n562), .ZN(new_n563));
  XOR2_X1   g377(.A(KEYINPUT24), .B(G110), .Z(new_n564));
  XNOR2_X1  g378(.A(G119), .B(G128), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XOR2_X1   g380(.A(new_n566), .B(KEYINPUT76), .Z(new_n567));
  NAND3_X1  g381(.A1(new_n555), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  OAI22_X1  g382(.A1(new_n560), .A2(G110), .B1(new_n565), .B2(new_n564), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(new_n225), .A3(new_n238), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n195), .A2(G221), .A3(G234), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT22), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(G137), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n568), .A2(new_n574), .A3(new_n570), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n262), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT25), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n576), .A2(KEYINPUT25), .A3(new_n262), .A4(new_n577), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n554), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n576), .A2(new_n577), .ZN(new_n583));
  AOI21_X1  g397(.A(G902), .B1(new_n296), .B2(new_n408), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n473), .A2(new_n553), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G101), .ZN(G3));
  XNOR2_X1  g402(.A(new_n299), .B(KEYINPUT33), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n301), .A2(G902), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n300), .A2(new_n301), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n272), .B2(new_n265), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n468), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n467), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n471), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n414), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n595), .A2(new_n412), .A3(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n402), .A2(new_n405), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n545), .A2(new_n547), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT31), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n491), .B1(new_n510), .B2(new_n488), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n604), .A2(new_n519), .B1(new_n540), .B2(new_n541), .ZN(new_n605));
  AOI21_X1  g419(.A(G902), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(G472), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n586), .B(new_n549), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n600), .A2(new_n601), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT34), .B(G104), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G6));
  NAND2_X1  g426(.A1(new_n265), .A2(new_n272), .ZN(new_n613));
  NOR4_X1   g427(.A1(new_n599), .A2(new_n303), .A3(new_n613), .A4(new_n412), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(new_n609), .A3(new_n601), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(new_n284), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT97), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n617), .B(KEYINPUT35), .Z(G9));
  OAI21_X1  g432(.A(new_n262), .B1(new_n543), .B2(new_n548), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(G472), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT36), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n574), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(new_n622), .B(KEYINPUT98), .Z(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n571), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n623), .A2(new_n568), .A3(new_n570), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n625), .A2(new_n584), .A3(new_n626), .ZN(new_n627));
  OR2_X1    g441(.A1(new_n582), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n473), .A2(new_n549), .A3(new_n620), .A4(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n629), .B(KEYINPUT37), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G110), .ZN(G12));
  INV_X1    g445(.A(new_n414), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n597), .B2(new_n471), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n402), .A2(new_n405), .A3(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n265), .A2(new_n272), .ZN(new_n635));
  INV_X1    g449(.A(G900), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n410), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(KEYINPUT99), .Z(new_n638));
  INV_X1    g452(.A(new_n407), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n303), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n553), .A2(new_n634), .A3(new_n628), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G128), .ZN(G30));
  XOR2_X1   g458(.A(new_n640), .B(KEYINPUT39), .Z(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n601), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT40), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n601), .A2(new_n649), .A3(new_n646), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n582), .A2(new_n627), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n303), .B1(new_n265), .B2(new_n272), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n470), .A2(new_n471), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT38), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n551), .A2(new_n552), .ZN(new_n660));
  INV_X1    g474(.A(new_n602), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n496), .B1(new_n513), .B2(new_n525), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n262), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G472), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n659), .A2(new_n665), .A3(new_n414), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n651), .A2(KEYINPUT100), .A3(new_n652), .A4(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT100), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n648), .A2(new_n652), .A3(new_n650), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n659), .A2(new_n665), .A3(new_n414), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(new_n197), .ZN(G45));
  NAND2_X1  g487(.A1(new_n594), .A2(new_n640), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n553), .A2(new_n634), .A3(new_n675), .A4(new_n628), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  AOI211_X1 g491(.A(G902), .B(new_n393), .C1(new_n388), .C2(new_n389), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n390), .A2(new_n262), .ZN(new_n679));
  AOI22_X1  g493(.A1(new_n678), .A2(new_n392), .B1(new_n679), .B2(G469), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT101), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n681), .A3(new_n405), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n679), .A2(G469), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n405), .A3(new_n395), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT101), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n600), .A2(new_n686), .A3(new_n553), .A4(new_n586), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT41), .B(G113), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  NAND4_X1  g503(.A1(new_n686), .A2(new_n614), .A3(new_n553), .A4(new_n586), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G116), .ZN(G18));
  AOI21_X1  g505(.A(new_n652), .B1(new_n660), .B2(new_n535), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(new_n684), .B2(new_n599), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n680), .A2(KEYINPUT102), .A3(new_n405), .A4(new_n633), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n692), .A2(new_n304), .A3(new_n413), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G119), .ZN(G21));
  OAI21_X1  g512(.A(KEYINPUT104), .B1(new_n654), .B2(new_n599), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n633), .A2(new_n653), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  OR3_X1    g516(.A1(new_n582), .A2(KEYINPUT103), .A3(new_n585), .ZN(new_n703));
  OAI21_X1  g517(.A(KEYINPUT103), .B1(new_n582), .B2(new_n585), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n519), .B1(new_n526), .B2(new_n529), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n603), .A2(new_n542), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n536), .ZN(new_n707));
  AND4_X1   g521(.A1(new_n620), .A2(new_n703), .A3(new_n704), .A4(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n702), .A2(new_n708), .A3(new_n413), .A4(new_n686), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G122), .ZN(G24));
  AOI22_X1  g524(.A1(new_n536), .A2(new_n706), .B1(new_n619), .B2(G472), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT105), .B1(new_n711), .B2(new_n628), .ZN(new_n712));
  AND4_X1   g526(.A1(KEYINPUT105), .A2(new_n707), .A3(new_n620), .A4(new_n628), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n675), .B(new_n696), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G125), .ZN(G27));
  XOR2_X1   g529(.A(new_n400), .B(KEYINPUT106), .Z(new_n716));
  NAND3_X1  g530(.A1(new_n395), .A2(new_n399), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n404), .A2(new_n632), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n717), .A2(new_n655), .A3(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n553), .A2(new_n586), .A3(new_n675), .A4(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT42), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n703), .A2(new_n704), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n660), .B2(new_n535), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n717), .A2(new_n655), .A3(new_n718), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n724), .A2(new_n674), .A3(new_n721), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n720), .A2(new_n721), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT107), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n199), .ZN(G33));
  NAND4_X1  g542(.A1(new_n553), .A2(new_n586), .A3(new_n642), .A4(new_n719), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G134), .ZN(G36));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n384), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(G469), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(KEYINPUT46), .A3(new_n716), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n733), .A2(new_n716), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT46), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n733), .A2(KEYINPUT108), .A3(KEYINPUT46), .A4(new_n716), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n736), .A2(new_n739), .A3(new_n395), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n405), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n645), .ZN(new_n743));
  INV_X1    g557(.A(new_n593), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n635), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n635), .A2(KEYINPUT43), .A3(new_n744), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n620), .A2(new_n549), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n749), .A2(KEYINPUT44), .A3(new_n750), .A4(new_n628), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n655), .A2(new_n414), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n749), .A2(new_n750), .A3(new_n628), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n743), .A2(new_n753), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G137), .ZN(G39));
  NAND2_X1  g573(.A1(new_n742), .A2(KEYINPUT47), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n553), .A2(new_n586), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n741), .A2(new_n762), .A3(new_n405), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n674), .A2(new_n754), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n760), .A2(new_n761), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G140), .ZN(G42));
  INV_X1    g580(.A(new_n722), .ZN(new_n767));
  INV_X1    g581(.A(new_n745), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n718), .A3(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n769), .A2(KEYINPUT110), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n657), .A2(new_n658), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n769), .B2(KEYINPUT110), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n683), .A2(new_n395), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT49), .ZN(new_n774));
  OR4_X1    g588(.A1(new_n665), .A2(new_n770), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n639), .B1(new_n747), .B2(new_n748), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n708), .A3(new_n632), .ZN(new_n777));
  INV_X1    g591(.A(new_n684), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n771), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n780));
  OR3_X1    g594(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n780), .B1(new_n777), .B2(new_n779), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n707), .A2(new_n620), .A3(new_n628), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT105), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n707), .A2(new_n620), .A3(new_n628), .A4(KEYINPUT105), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n754), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n778), .A3(new_n789), .A4(new_n776), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n586), .A2(new_n407), .ZN(new_n791));
  NOR4_X1   g605(.A1(new_n665), .A2(new_n684), .A3(new_n754), .A4(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n635), .A3(new_n593), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n783), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n741), .A2(new_n762), .A3(new_n405), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n762), .B1(new_n741), .B2(new_n405), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT116), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n760), .A2(new_n798), .A3(new_n763), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n773), .A2(new_n405), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n797), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n776), .A2(new_n708), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(new_n789), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n794), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n805), .A2(KEYINPUT51), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n803), .A2(new_n696), .ZN(new_n808));
  AOI211_X1 g622(.A(new_n406), .B(G953), .C1(new_n792), .C2(new_n594), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n723), .A2(new_n778), .A3(new_n776), .A4(new_n789), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n810), .A2(KEYINPUT48), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(KEYINPUT48), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n809), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n783), .A2(new_n790), .A3(new_n793), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n801), .B1(new_n795), .B2(new_n796), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n815), .B1(new_n816), .B2(new_n804), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n813), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n806), .A2(new_n807), .A3(new_n808), .A4(new_n818), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n818), .B(new_n808), .C1(new_n805), .C2(KEYINPUT51), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT117), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n404), .B1(new_n638), .B2(new_n639), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n717), .A2(new_n652), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n717), .A2(new_n652), .A3(KEYINPUT113), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n665), .A3(new_n702), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n714), .A2(new_n831), .A3(new_n643), .A4(new_n676), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT52), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n402), .A2(new_n405), .A3(new_n472), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n609), .A2(new_n834), .A3(new_n594), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n587), .A2(KEYINPUT111), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT111), .B1(new_n587), .B2(new_n835), .ZN(new_n838));
  XOR2_X1   g652(.A(new_n303), .B(KEYINPUT112), .Z(new_n839));
  NAND4_X1  g653(.A1(new_n609), .A2(new_n834), .A3(new_n635), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n629), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n837), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  AOI211_X1 g656(.A(new_n674), .B(new_n724), .C1(new_n786), .C2(new_n787), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n754), .A2(new_n839), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n641), .A2(new_n652), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n553), .A2(new_n844), .A3(new_n601), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n729), .A2(new_n846), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n726), .A2(new_n843), .A3(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n697), .A2(new_n687), .A3(new_n690), .A4(new_n709), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n842), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n833), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n720), .A2(new_n721), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n723), .A2(new_n725), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n788), .A2(new_n675), .A3(new_n719), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n729), .A3(new_n857), .A4(new_n846), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n587), .A2(new_n835), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT111), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n629), .A2(new_n840), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n862), .A3(new_n836), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n858), .A2(new_n863), .A3(new_n849), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT52), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n832), .B(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT53), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n824), .B1(new_n853), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n852), .B1(new_n833), .B2(new_n851), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT114), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n823), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n864), .A2(new_n866), .A3(KEYINPUT53), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n869), .A2(new_n872), .A3(new_n823), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT115), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT114), .B1(new_n869), .B2(new_n872), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n867), .A2(new_n824), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT54), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n869), .A2(new_n872), .A3(new_n823), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n822), .B1(new_n874), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(G952), .A2(G953), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n775), .B1(new_n881), .B2(new_n882), .ZN(G75));
  NAND2_X1  g697(.A1(new_n442), .A2(new_n444), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(new_n453), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT55), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n262), .B1(new_n869), .B2(new_n872), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(G210), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n195), .A2(G952), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n886), .A2(new_n889), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n887), .B2(new_n469), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(G51));
  XOR2_X1   g708(.A(new_n716), .B(KEYINPUT57), .Z(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT54), .B1(new_n853), .B2(new_n867), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n896), .B1(new_n897), .B2(new_n879), .ZN(new_n898));
  INV_X1    g712(.A(new_n390), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT118), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n823), .B1(new_n869), .B2(new_n872), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n895), .B1(new_n873), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n903), .A3(new_n390), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n887), .A2(G469), .A3(new_n732), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n900), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n891), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(G54));
  NAND3_X1  g722(.A1(new_n887), .A2(KEYINPUT58), .A3(G475), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n248), .A2(new_n260), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n909), .A2(new_n911), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n912), .A2(new_n913), .A3(new_n891), .ZN(G60));
  NAND2_X1  g728(.A1(G478), .A2(G902), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT59), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n589), .B(KEYINPUT119), .Z(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n916), .B(new_n918), .C1(new_n873), .C2(new_n901), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n907), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n874), .A2(new_n880), .A3(new_n916), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n920), .B1(new_n921), .B2(new_n917), .ZN(G63));
  NAND2_X1  g736(.A1(new_n869), .A2(new_n872), .ZN(new_n923));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT60), .Z(new_n925));
  AOI21_X1  g739(.A(new_n583), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT120), .B1(new_n926), .B2(new_n891), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT120), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n625), .A2(new_n626), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n928), .B1(new_n930), .B2(KEYINPUT121), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n930), .A2(KEYINPUT121), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n923), .A2(new_n925), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n927), .A2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(G66));
  INV_X1    g750(.A(G224), .ZN(new_n937));
  OAI21_X1  g751(.A(G953), .B1(new_n411), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n863), .A2(new_n849), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n938), .B1(new_n939), .B2(G953), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n884), .B1(G898), .B2(new_n195), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT122), .Z(new_n942));
  XNOR2_X1  g756(.A(new_n940), .B(new_n942), .ZN(G69));
  NAND2_X1  g757(.A1(new_n515), .A2(new_n516), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n249), .A2(new_n251), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n944), .B(new_n945), .Z(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n636), .B2(G953), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n758), .A2(new_n765), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n743), .A2(new_n702), .A3(new_n723), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n714), .A2(new_n643), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n676), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n951), .A2(new_n726), .ZN(new_n952));
  AND4_X1   g766(.A1(new_n729), .A2(new_n948), .A3(new_n949), .A4(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n947), .B1(new_n953), .B2(G953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n950), .A2(new_n676), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n955), .A2(KEYINPUT62), .A3(new_n671), .A4(new_n667), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n672), .B2(new_n951), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n594), .B1(new_n839), .B2(new_n635), .ZN(new_n960));
  AOI211_X1 g774(.A(new_n754), .B(new_n647), .C1(KEYINPUT123), .C2(new_n960), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n960), .A2(KEYINPUT123), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n961), .A2(new_n553), .A3(new_n586), .A4(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT124), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n959), .A2(new_n948), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n966), .A2(new_n195), .A3(new_n946), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n954), .A2(KEYINPUT125), .A3(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n946), .A2(KEYINPUT125), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n969), .A2(G227), .ZN(new_n970));
  OAI21_X1  g784(.A(G953), .B1(new_n970), .B2(new_n636), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n968), .B(new_n971), .ZN(G72));
  INV_X1    g786(.A(new_n518), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n953), .A2(new_n939), .ZN(new_n974));
  XNOR2_X1  g788(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n607), .A2(new_n262), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n973), .B(new_n519), .C1(new_n974), .C2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n959), .A2(new_n939), .A3(new_n948), .A4(new_n965), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n977), .ZN(new_n982));
  AND4_X1   g796(.A1(new_n980), .A2(new_n982), .A3(new_n518), .A4(new_n496), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n519), .B1(new_n981), .B2(new_n977), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n980), .B1(new_n984), .B2(new_n518), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n979), .B(new_n907), .C1(new_n983), .C2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n602), .A2(new_n520), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n977), .B(new_n987), .C1(new_n875), .C2(new_n876), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n986), .A2(new_n989), .ZN(G57));
endmodule


