

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581;

  XNOR2_X1 U323 ( .A(n379), .B(n378), .ZN(n547) );
  XNOR2_X1 U324 ( .A(n447), .B(KEYINPUT38), .ZN(n494) );
  XOR2_X1 U325 ( .A(n309), .B(n308), .Z(n520) );
  XNOR2_X1 U326 ( .A(n414), .B(n413), .ZN(n513) );
  XNOR2_X1 U327 ( .A(KEYINPUT94), .B(n440), .ZN(n533) );
  XOR2_X1 U328 ( .A(n368), .B(KEYINPUT9), .Z(n291) );
  XNOR2_X1 U329 ( .A(n458), .B(n457), .ZN(n459) );
  NAND2_X1 U330 ( .A1(n444), .A2(n443), .ZN(n477) );
  XOR2_X1 U331 ( .A(G36GAT), .B(n374), .Z(n405) );
  XNOR2_X1 U332 ( .A(n405), .B(n377), .ZN(n378) );
  NOR2_X1 U333 ( .A1(n572), .A2(n445), .ZN(n446) );
  NOR2_X1 U334 ( .A1(n560), .A2(n415), .ZN(n535) );
  NOR2_X1 U335 ( .A1(n520), .A2(n470), .ZN(n555) );
  INV_X1 U336 ( .A(G43GAT), .ZN(n448) );
  XNOR2_X1 U337 ( .A(n471), .B(G176GAT), .ZN(n472) );
  XNOR2_X1 U338 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U339 ( .A(n473), .B(n472), .ZN(G1349GAT) );
  XNOR2_X1 U340 ( .A(n451), .B(n450), .ZN(G1330GAT) );
  XOR2_X1 U341 ( .A(G176GAT), .B(G127GAT), .Z(n293) );
  XNOR2_X1 U342 ( .A(G15GAT), .B(G183GAT), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n293), .B(n292), .ZN(n309) );
  XOR2_X1 U344 ( .A(G71GAT), .B(G120GAT), .Z(n295) );
  XNOR2_X1 U345 ( .A(G134GAT), .B(G99GAT), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U347 ( .A(n296), .B(G190GAT), .Z(n298) );
  XOR2_X1 U348 ( .A(G113GAT), .B(KEYINPUT0), .Z(n422) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(n422), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U351 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n300) );
  NAND2_X1 U352 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U354 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U355 ( .A(KEYINPUT87), .B(KEYINPUT17), .Z(n304) );
  XNOR2_X1 U356 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U358 ( .A(G169GAT), .B(n305), .Z(n414) );
  XNOR2_X1 U359 ( .A(n414), .B(KEYINPUT86), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U361 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n311) );
  XNOR2_X1 U362 ( .A(G8GAT), .B(KEYINPUT69), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n329) );
  XOR2_X1 U364 ( .A(G113GAT), .B(G29GAT), .Z(n313) );
  XNOR2_X1 U365 ( .A(G50GAT), .B(G36GAT), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U367 ( .A(G1GAT), .B(G141GAT), .Z(n315) );
  XNOR2_X1 U368 ( .A(G169GAT), .B(G197GAT), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U370 ( .A(n317), .B(n316), .Z(n327) );
  XOR2_X1 U371 ( .A(KEYINPUT68), .B(KEYINPUT73), .Z(n319) );
  XNOR2_X1 U372 ( .A(KEYINPUT71), .B(KEYINPUT70), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n325) );
  XOR2_X1 U374 ( .A(G43GAT), .B(KEYINPUT7), .Z(n321) );
  XNOR2_X1 U375 ( .A(KEYINPUT8), .B(KEYINPUT72), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n368) );
  XOR2_X1 U377 ( .A(G15GAT), .B(G22GAT), .Z(n347) );
  XOR2_X1 U378 ( .A(n368), .B(n347), .Z(n323) );
  NAND2_X1 U379 ( .A1(G229GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U383 ( .A(n329), .B(n328), .Z(n536) );
  INV_X1 U384 ( .A(n536), .ZN(n563) );
  XNOR2_X1 U385 ( .A(G120GAT), .B(G148GAT), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n330), .B(G57GAT), .ZN(n421) );
  XNOR2_X1 U387 ( .A(G99GAT), .B(G106GAT), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n331), .B(KEYINPUT76), .ZN(n376) );
  XNOR2_X1 U389 ( .A(n421), .B(n376), .ZN(n344) );
  XOR2_X1 U390 ( .A(G71GAT), .B(KEYINPUT13), .Z(n346) );
  XOR2_X1 U391 ( .A(G176GAT), .B(G64GAT), .Z(n401) );
  XOR2_X1 U392 ( .A(n346), .B(n401), .Z(n333) );
  NAND2_X1 U393 ( .A1(G230GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U394 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U395 ( .A(KEYINPUT32), .B(KEYINPUT77), .Z(n335) );
  XNOR2_X1 U396 ( .A(KEYINPUT74), .B(KEYINPUT33), .ZN(n334) );
  XNOR2_X1 U397 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U398 ( .A(n337), .B(n336), .Z(n342) );
  XOR2_X1 U399 ( .A(KEYINPUT75), .B(G78GAT), .Z(n383) );
  XOR2_X1 U400 ( .A(KEYINPUT31), .B(G92GAT), .Z(n339) );
  XNOR2_X1 U401 ( .A(G204GAT), .B(G85GAT), .ZN(n338) );
  XNOR2_X1 U402 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n383), .B(n340), .ZN(n341) );
  XNOR2_X1 U404 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U405 ( .A(n344), .B(n343), .ZN(n566) );
  NAND2_X1 U406 ( .A1(n563), .A2(n566), .ZN(n345) );
  XOR2_X1 U407 ( .A(KEYINPUT78), .B(n345), .Z(n480) );
  XOR2_X1 U408 ( .A(G8GAT), .B(G183GAT), .Z(n402) );
  XOR2_X1 U409 ( .A(n346), .B(n402), .Z(n349) );
  XOR2_X1 U410 ( .A(G1GAT), .B(G127GAT), .Z(n430) );
  XNOR2_X1 U411 ( .A(n347), .B(n430), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n362) );
  XOR2_X1 U413 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n351) );
  NAND2_X1 U414 ( .A1(G231GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U415 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U416 ( .A(n352), .B(KEYINPUT12), .Z(n360) );
  XOR2_X1 U417 ( .A(G57GAT), .B(G78GAT), .Z(n354) );
  XNOR2_X1 U418 ( .A(G155GAT), .B(G211GAT), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U420 ( .A(KEYINPUT83), .B(KEYINPUT14), .Z(n356) );
  XNOR2_X1 U421 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n355) );
  XNOR2_X1 U422 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n362), .B(n361), .ZN(n572) );
  XOR2_X1 U426 ( .A(KEYINPUT79), .B(KEYINPUT10), .Z(n364) );
  XNOR2_X1 U427 ( .A(KEYINPUT11), .B(KEYINPUT67), .ZN(n363) );
  XNOR2_X1 U428 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U429 ( .A(n365), .B(KEYINPUT65), .Z(n367) );
  XOR2_X1 U430 ( .A(G50GAT), .B(G162GAT), .Z(n384) );
  XNOR2_X1 U431 ( .A(n384), .B(KEYINPUT81), .ZN(n366) );
  XNOR2_X1 U432 ( .A(n367), .B(n366), .ZN(n371) );
  NAND2_X1 U433 ( .A1(G232GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U434 ( .A(n291), .B(n369), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n371), .B(n370), .ZN(n379) );
  XOR2_X1 U436 ( .A(G92GAT), .B(KEYINPUT80), .Z(n373) );
  XNOR2_X1 U437 ( .A(G190GAT), .B(G218GAT), .ZN(n372) );
  XNOR2_X1 U438 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U439 ( .A(G29GAT), .B(G134GAT), .ZN(n375) );
  XNOR2_X1 U440 ( .A(n375), .B(G85GAT), .ZN(n434) );
  XOR2_X1 U441 ( .A(n434), .B(n376), .Z(n377) );
  XNOR2_X1 U442 ( .A(KEYINPUT82), .B(n547), .ZN(n554) );
  XOR2_X1 U443 ( .A(KEYINPUT36), .B(KEYINPUT107), .Z(n380) );
  XNOR2_X1 U444 ( .A(n554), .B(n380), .ZN(n576) );
  XOR2_X1 U445 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n382) );
  XNOR2_X1 U446 ( .A(KEYINPUT90), .B(KEYINPUT24), .ZN(n381) );
  XNOR2_X1 U447 ( .A(n382), .B(n381), .ZN(n388) );
  XOR2_X1 U448 ( .A(G106GAT), .B(G218GAT), .Z(n386) );
  XNOR2_X1 U449 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U450 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U451 ( .A(n388), .B(n387), .Z(n390) );
  NAND2_X1 U452 ( .A1(G228GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U454 ( .A(n391), .B(G148GAT), .Z(n395) );
  XOR2_X1 U455 ( .A(G204GAT), .B(G211GAT), .Z(n393) );
  XNOR2_X1 U456 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n392) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n406) );
  XNOR2_X1 U458 ( .A(G22GAT), .B(n406), .ZN(n394) );
  XNOR2_X1 U459 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U460 ( .A(KEYINPUT89), .B(KEYINPUT2), .Z(n397) );
  XNOR2_X1 U461 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U463 ( .A(G141GAT), .B(n398), .ZN(n426) );
  XNOR2_X1 U464 ( .A(n399), .B(n426), .ZN(n467) );
  NAND2_X1 U465 ( .A1(n467), .A2(n520), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n400), .B(KEYINPUT26), .ZN(n560) );
  XOR2_X1 U467 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n404) );
  XNOR2_X1 U468 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U469 ( .A(n404), .B(n403), .ZN(n410) );
  XOR2_X1 U470 ( .A(KEYINPUT98), .B(KEYINPUT95), .Z(n408) );
  XNOR2_X1 U471 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U472 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U473 ( .A(n410), .B(n409), .Z(n412) );
  NAND2_X1 U474 ( .A1(G226GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U476 ( .A(KEYINPUT27), .B(n513), .Z(n441) );
  INV_X1 U477 ( .A(n441), .ZN(n415) );
  XNOR2_X1 U478 ( .A(n535), .B(KEYINPUT99), .ZN(n420) );
  NOR2_X1 U479 ( .A1(n520), .A2(n513), .ZN(n416) );
  XNOR2_X1 U480 ( .A(n416), .B(KEYINPUT100), .ZN(n417) );
  NOR2_X1 U481 ( .A1(n467), .A2(n417), .ZN(n418) );
  XNOR2_X1 U482 ( .A(KEYINPUT25), .B(n418), .ZN(n419) );
  NAND2_X1 U483 ( .A1(n420), .A2(n419), .ZN(n439) );
  XOR2_X1 U484 ( .A(n422), .B(n421), .Z(n424) );
  NAND2_X1 U485 ( .A1(G225GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U486 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U487 ( .A(n426), .B(n425), .Z(n438) );
  XOR2_X1 U488 ( .A(KEYINPUT1), .B(KEYINPUT91), .Z(n428) );
  XNOR2_X1 U489 ( .A(KEYINPUT5), .B(KEYINPUT6), .ZN(n427) );
  XNOR2_X1 U490 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U491 ( .A(n429), .B(KEYINPUT93), .Z(n432) );
  XNOR2_X1 U492 ( .A(G162GAT), .B(n430), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U494 ( .A(n433), .B(KEYINPUT4), .Z(n436) );
  XNOR2_X1 U495 ( .A(n434), .B(KEYINPUT92), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n440) );
  NAND2_X1 U498 ( .A1(n439), .A2(n440), .ZN(n444) );
  XOR2_X1 U499 ( .A(n467), .B(KEYINPUT28), .Z(n517) );
  NAND2_X1 U500 ( .A1(n517), .A2(n441), .ZN(n442) );
  NOR2_X1 U501 ( .A1(n533), .A2(n442), .ZN(n522) );
  NAND2_X1 U502 ( .A1(n520), .A2(n522), .ZN(n443) );
  NAND2_X1 U503 ( .A1(n576), .A2(n477), .ZN(n445) );
  XOR2_X1 U504 ( .A(KEYINPUT37), .B(n446), .Z(n510) );
  NAND2_X1 U505 ( .A1(n480), .A2(n510), .ZN(n447) );
  NOR2_X1 U506 ( .A1(n520), .A2(n494), .ZN(n451) );
  XNOR2_X1 U507 ( .A(KEYINPUT40), .B(KEYINPUT108), .ZN(n449) );
  XNOR2_X1 U508 ( .A(KEYINPUT119), .B(KEYINPUT55), .ZN(n469) );
  XNOR2_X1 U509 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n452) );
  XOR2_X1 U510 ( .A(n566), .B(n452), .Z(n541) );
  INV_X1 U511 ( .A(n541), .ZN(n496) );
  NAND2_X1 U512 ( .A1(n496), .A2(n563), .ZN(n453) );
  XNOR2_X1 U513 ( .A(KEYINPUT46), .B(n453), .ZN(n454) );
  INV_X1 U514 ( .A(n572), .ZN(n544) );
  NAND2_X1 U515 ( .A1(n454), .A2(n544), .ZN(n455) );
  NOR2_X1 U516 ( .A1(n547), .A2(n455), .ZN(n456) );
  XOR2_X1 U517 ( .A(KEYINPUT47), .B(n456), .Z(n463) );
  NAND2_X1 U518 ( .A1(n576), .A2(n572), .ZN(n458) );
  XOR2_X1 U519 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n457) );
  NAND2_X1 U520 ( .A1(n459), .A2(n566), .ZN(n460) );
  NOR2_X1 U521 ( .A1(n563), .A2(n460), .ZN(n461) );
  XNOR2_X1 U522 ( .A(KEYINPUT114), .B(n461), .ZN(n462) );
  NOR2_X1 U523 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U524 ( .A(n464), .B(KEYINPUT48), .ZN(n532) );
  NOR2_X1 U525 ( .A1(n513), .A2(n532), .ZN(n465) );
  XNOR2_X1 U526 ( .A(n465), .B(KEYINPUT54), .ZN(n466) );
  NAND2_X1 U527 ( .A1(n466), .A2(n533), .ZN(n561) );
  NOR2_X1 U528 ( .A1(n561), .A2(n467), .ZN(n468) );
  XOR2_X1 U529 ( .A(n469), .B(n468), .Z(n470) );
  NAND2_X1 U530 ( .A1(n555), .A2(n496), .ZN(n473) );
  XOR2_X1 U531 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n471) );
  XOR2_X1 U532 ( .A(KEYINPUT103), .B(KEYINPUT34), .Z(n475) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(KEYINPUT104), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n475), .B(n474), .ZN(n483) );
  NOR2_X1 U535 ( .A1(n544), .A2(n554), .ZN(n476) );
  XNOR2_X1 U536 ( .A(KEYINPUT16), .B(n476), .ZN(n478) );
  NAND2_X1 U537 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n479), .B(KEYINPUT101), .ZN(n498) );
  NAND2_X1 U539 ( .A1(n480), .A2(n498), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n481), .B(KEYINPUT102), .ZN(n489) );
  NOR2_X1 U541 ( .A1(n489), .A2(n533), .ZN(n482) );
  XOR2_X1 U542 ( .A(n483), .B(n482), .Z(G1324GAT) );
  NOR2_X1 U543 ( .A1(n489), .A2(n513), .ZN(n484) );
  XOR2_X1 U544 ( .A(G8GAT), .B(n484), .Z(G1325GAT) );
  NOR2_X1 U545 ( .A1(n489), .A2(n520), .ZN(n488) );
  XOR2_X1 U546 ( .A(KEYINPUT105), .B(KEYINPUT35), .Z(n486) );
  XNOR2_X1 U547 ( .A(G15GAT), .B(KEYINPUT106), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(G1326GAT) );
  NOR2_X1 U550 ( .A1(n517), .A2(n489), .ZN(n490) );
  XOR2_X1 U551 ( .A(G22GAT), .B(n490), .Z(G1327GAT) );
  NOR2_X1 U552 ( .A1(n494), .A2(n533), .ZN(n492) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  NOR2_X1 U555 ( .A1(n494), .A2(n513), .ZN(n493) );
  XOR2_X1 U556 ( .A(G36GAT), .B(n493), .Z(G1329GAT) );
  NOR2_X1 U557 ( .A1(n517), .A2(n494), .ZN(n495) );
  XOR2_X1 U558 ( .A(G50GAT), .B(n495), .Z(G1331GAT) );
  NAND2_X1 U559 ( .A1(n496), .A2(n536), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n497), .B(KEYINPUT109), .ZN(n509) );
  NAND2_X1 U561 ( .A1(n509), .A2(n498), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n499), .B(KEYINPUT110), .ZN(n504) );
  NOR2_X1 U563 ( .A1(n504), .A2(n533), .ZN(n500) );
  XOR2_X1 U564 ( .A(G57GAT), .B(n500), .Z(n501) );
  XNOR2_X1 U565 ( .A(KEYINPUT42), .B(n501), .ZN(G1332GAT) );
  NOR2_X1 U566 ( .A1(n504), .A2(n513), .ZN(n502) );
  XOR2_X1 U567 ( .A(G64GAT), .B(n502), .Z(G1333GAT) );
  NOR2_X1 U568 ( .A1(n520), .A2(n504), .ZN(n503) );
  XOR2_X1 U569 ( .A(G71GAT), .B(n503), .Z(G1334GAT) );
  NOR2_X1 U570 ( .A1(n504), .A2(n517), .ZN(n508) );
  XOR2_X1 U571 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n506) );
  XNOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT112), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(G1335GAT) );
  NAND2_X1 U575 ( .A1(n510), .A2(n509), .ZN(n516) );
  NOR2_X1 U576 ( .A1(n533), .A2(n516), .ZN(n512) );
  XNOR2_X1 U577 ( .A(G85GAT), .B(KEYINPUT113), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(G1336GAT) );
  NOR2_X1 U579 ( .A1(n513), .A2(n516), .ZN(n514) );
  XOR2_X1 U580 ( .A(G92GAT), .B(n514), .Z(G1337GAT) );
  NOR2_X1 U581 ( .A1(n520), .A2(n516), .ZN(n515) );
  XOR2_X1 U582 ( .A(G99GAT), .B(n515), .Z(G1338GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n518) );
  XOR2_X1 U584 ( .A(KEYINPUT44), .B(n518), .Z(n519) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(n519), .ZN(G1339GAT) );
  NOR2_X1 U586 ( .A1(n520), .A2(n532), .ZN(n521) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n528) );
  NOR2_X1 U588 ( .A1(n536), .A2(n528), .ZN(n523) );
  XOR2_X1 U589 ( .A(G113GAT), .B(n523), .Z(G1340GAT) );
  NOR2_X1 U590 ( .A1(n541), .A2(n528), .ZN(n525) );
  XNOR2_X1 U591 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(G1341GAT) );
  NOR2_X1 U593 ( .A1(n544), .A2(n528), .ZN(n526) );
  XOR2_X1 U594 ( .A(KEYINPUT50), .B(n526), .Z(n527) );
  XNOR2_X1 U595 ( .A(G127GAT), .B(n527), .ZN(G1342GAT) );
  XOR2_X1 U596 ( .A(G134GAT), .B(KEYINPUT51), .Z(n531) );
  INV_X1 U597 ( .A(n528), .ZN(n529) );
  NAND2_X1 U598 ( .A1(n529), .A2(n554), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(G1343GAT) );
  NOR2_X1 U600 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n546) );
  NOR2_X1 U602 ( .A1(n536), .A2(n546), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(G1344GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n540) );
  XNOR2_X1 U606 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n543) );
  NOR2_X1 U608 ( .A1(n541), .A2(n546), .ZN(n542) );
  XOR2_X1 U609 ( .A(n543), .B(n542), .Z(G1345GAT) );
  NOR2_X1 U610 ( .A1(n544), .A2(n546), .ZN(n545) );
  XOR2_X1 U611 ( .A(G155GAT), .B(n545), .Z(G1346GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n550) );
  INV_X1 U613 ( .A(n546), .ZN(n548) );
  NAND2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(n551), .ZN(G1347GAT) );
  NAND2_X1 U617 ( .A1(n555), .A2(n563), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G169GAT), .B(n552), .ZN(G1348GAT) );
  NAND2_X1 U619 ( .A1(n572), .A2(n555), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(KEYINPUT58), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G190GAT), .B(n557), .ZN(G1351GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n559) );
  XNOR2_X1 U625 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n565) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U628 ( .A(n562), .B(KEYINPUT120), .Z(n567) );
  INV_X1 U629 ( .A(n567), .ZN(n577) );
  NAND2_X1 U630 ( .A1(n577), .A2(n563), .ZN(n564) );
  XOR2_X1 U631 ( .A(n565), .B(n564), .Z(G1352GAT) );
  NOR2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT122), .B(KEYINPUT61), .Z(n569) );
  XNOR2_X1 U634 ( .A(G204GAT), .B(KEYINPUT123), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1353GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n574) );
  NAND2_X1 U638 ( .A1(n577), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(n575), .ZN(G1354GAT) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT127), .B(KEYINPUT126), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(G1355GAT) );
endmodule

