//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1017,
    new_n1018, new_n1019, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062;
  INV_X1    g000(.A(KEYINPUT67), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT67), .A2(G953), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n189), .A2(G210), .A3(new_n190), .A4(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT69), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT26), .B(G101), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT67), .A2(G953), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT67), .A2(G953), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT69), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G210), .A4(new_n190), .ZN(new_n202));
  XOR2_X1   g016(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(new_n194), .ZN(new_n204));
  AND4_X1   g018(.A1(new_n193), .A2(new_n197), .A3(new_n202), .A4(new_n204), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n197), .A2(new_n204), .B1(new_n193), .B2(new_n202), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  AND2_X1   g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT64), .A3(new_n212), .ZN(new_n217));
  INV_X1    g031(.A(new_n216), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n212), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n215), .A2(new_n217), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT11), .ZN(new_n222));
  INV_X1    g036(.A(G134), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n222), .B1(new_n223), .B2(G137), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(G137), .ZN(new_n225));
  INV_X1    g039(.A(G137), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(KEYINPUT11), .A3(G134), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n224), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G131), .ZN(new_n229));
  INV_X1    g043(.A(G131), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n224), .A2(new_n227), .A3(new_n230), .A4(new_n225), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n221), .A2(new_n232), .ZN(new_n233));
  XOR2_X1   g047(.A(KEYINPUT2), .B(G113), .Z(new_n234));
  INV_X1    g048(.A(G116), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT66), .B1(new_n235), .B2(G119), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n237));
  INV_X1    g051(.A(G119), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n238), .A3(G116), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n238), .A2(G116), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n234), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n241), .B1(new_n236), .B2(new_n239), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(new_n234), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G128), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(KEYINPUT1), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n216), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n247), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n249), .B1(new_n216), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n223), .A2(G137), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n226), .A2(G134), .ZN(new_n253));
  OAI21_X1  g067(.A(G131), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(new_n231), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n233), .A2(new_n246), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n256), .B(KEYINPUT28), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT65), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT1), .B1(new_n210), .B2(G146), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n259), .A2(G128), .B1(new_n209), .B2(new_n211), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n248), .A2(new_n209), .A3(new_n211), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n231), .A2(new_n254), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n258), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n251), .A2(KEYINPUT65), .A3(new_n231), .A4(new_n254), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n264), .A2(new_n265), .B1(new_n232), .B2(new_n221), .ZN(new_n266));
  OR2_X1    g080(.A1(new_n266), .A2(new_n246), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n207), .B1(new_n257), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n256), .B2(new_n207), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n256), .A2(new_n207), .A3(new_n270), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n244), .B(new_n234), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n233), .A2(KEYINPUT30), .A3(new_n255), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n275), .B(new_n276), .C1(new_n266), .C2(KEYINPUT30), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT31), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n256), .A2(new_n207), .A3(new_n270), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n277), .B(KEYINPUT31), .C1(new_n279), .C2(new_n271), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n269), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(G472), .A2(G902), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(KEYINPUT32), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT32), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n277), .B1(new_n279), .B2(new_n271), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT31), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n268), .B1(new_n288), .B2(new_n280), .ZN(new_n289));
  INV_X1    g103(.A(new_n283), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n285), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT28), .ZN(new_n292));
  OR2_X1    g106(.A1(new_n256), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n256), .A2(new_n292), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n205), .A2(new_n206), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n233), .A2(new_n255), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n275), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n293), .A2(new_n294), .A3(new_n296), .A4(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n257), .A2(new_n267), .A3(new_n207), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n295), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n207), .B1(new_n277), .B2(new_n256), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n301), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G472), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n284), .A2(new_n291), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n284), .A2(new_n291), .A3(new_n306), .A4(KEYINPUT71), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT9), .B(G234), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT75), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n312), .B(new_n313), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n188), .A2(G217), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT92), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n314), .A2(KEYINPUT92), .A3(new_n315), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G122), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G116), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n235), .A2(G122), .ZN(new_n323));
  INV_X1    g137(.A(G107), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT90), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n324), .B1(new_n322), .B2(new_n323), .ZN(new_n328));
  OR3_X1    g142(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n327), .B1(new_n326), .B2(new_n328), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G128), .B(G143), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT13), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n210), .A2(G128), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n333), .B(G134), .C1(KEYINPUT13), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(new_n223), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n331), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n323), .A2(KEYINPUT91), .A3(KEYINPUT14), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT91), .B1(new_n323), .B2(KEYINPUT14), .ZN(new_n340));
  OAI221_X1 g154(.A(new_n322), .B1(KEYINPUT14), .B2(new_n323), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G107), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n332), .B(new_n223), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n325), .A3(new_n343), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n320), .A2(new_n337), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n320), .B1(new_n344), .B2(new_n337), .ZN(new_n346));
  OAI211_X1 g160(.A(KEYINPUT93), .B(new_n300), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G478), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(KEYINPUT15), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n337), .A2(new_n344), .ZN(new_n351));
  INV_X1    g165(.A(new_n320), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n320), .A2(new_n337), .A3(new_n344), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n349), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n355), .A2(KEYINPUT93), .A3(new_n300), .A4(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n350), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G140), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G125), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(KEYINPUT16), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n360), .A2(KEYINPUT72), .A3(G125), .ZN(new_n364));
  XNOR2_X1  g178(.A(G125), .B(G140), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n364), .B1(new_n365), .B2(KEYINPUT72), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT16), .ZN(new_n367));
  OAI211_X1 g181(.A(G146), .B(new_n363), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT73), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n364), .ZN(new_n371));
  INV_X1    g185(.A(G125), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G140), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n361), .A3(KEYINPUT72), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT16), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n376), .A2(KEYINPUT73), .A3(G146), .A4(new_n363), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n367), .B1(new_n371), .B2(new_n374), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n208), .B1(new_n378), .B2(new_n362), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n370), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n189), .A2(G214), .A3(new_n190), .A4(new_n191), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n381), .A2(new_n210), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(new_n210), .ZN(new_n383));
  OAI21_X1  g197(.A(G131), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT85), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n381), .A2(new_n210), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n200), .A2(G143), .A3(G214), .A4(new_n190), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT85), .A3(G131), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n380), .B1(new_n391), .B2(KEYINPUT17), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT85), .B1(new_n389), .B2(G131), .ZN(new_n393));
  AOI211_X1 g207(.A(new_n385), .B(new_n230), .C1(new_n387), .C2(new_n388), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT17), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n387), .A2(new_n388), .A3(new_n230), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT84), .A4(new_n230), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n395), .A2(new_n396), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n365), .A2(new_n208), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(new_n375), .B2(new_n208), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT18), .A2(G131), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n389), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n389), .A2(new_n404), .ZN(new_n407));
  OR2_X1    g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n392), .A2(new_n401), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G113), .B(G122), .ZN(new_n410));
  INV_X1    g224(.A(G104), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n410), .B(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(KEYINPUT89), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n300), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n370), .A2(new_n379), .A3(new_n377), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT17), .B1(new_n393), .B2(new_n394), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n386), .A2(new_n390), .A3(new_n399), .A4(new_n400), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n415), .B(new_n416), .C1(new_n417), .C2(KEYINPUT17), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n403), .B1(new_n406), .B2(new_n407), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n418), .A2(new_n419), .A3(new_n413), .ZN(new_n420));
  OAI21_X1  g234(.A(G475), .B1(new_n414), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n422));
  INV_X1    g236(.A(new_n412), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(new_n418), .B2(new_n419), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n419), .A2(new_n423), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n365), .A2(KEYINPUT86), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n375), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(KEYINPUT86), .A2(KEYINPUT19), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n427), .A2(KEYINPUT19), .B1(new_n365), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n208), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n430), .A2(new_n368), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n425), .B1(new_n417), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT87), .B1(new_n424), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n417), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n419), .A3(new_n423), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n435), .B(new_n436), .C1(new_n409), .C2(new_n423), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(G475), .A2(G902), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n422), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n399), .A2(new_n400), .ZN(new_n441));
  NOR4_X1   g255(.A1(new_n441), .A2(new_n393), .A3(new_n394), .A4(KEYINPUT17), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n415), .A2(new_n416), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n419), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n412), .ZN(new_n445));
  INV_X1    g259(.A(new_n439), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(KEYINPUT20), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n435), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT88), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT88), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n445), .A2(new_n450), .A3(new_n435), .A4(new_n447), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n359), .B(new_n421), .C1(new_n440), .C2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G234), .ZN(new_n455));
  OAI21_X1  g269(.A(G217), .B1(new_n455), .B2(G902), .ZN(new_n456));
  XOR2_X1   g270(.A(G119), .B(G128), .Z(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT24), .B(G110), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT23), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n238), .B2(G128), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n247), .A2(KEYINPUT23), .A3(G119), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n461), .B(new_n462), .C1(G119), .C2(new_n247), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n459), .B1(G110), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n380), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n457), .A2(new_n458), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n463), .B2(G110), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n368), .A2(new_n402), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n200), .A2(G221), .A3(G234), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT22), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(G137), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n472), .B(new_n226), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n465), .A2(new_n475), .A3(new_n468), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n474), .A2(new_n300), .A3(new_n476), .ZN(new_n477));
  AND2_X1   g291(.A1(KEYINPUT74), .A2(KEYINPUT25), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n456), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(KEYINPUT74), .A2(KEYINPUT25), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n474), .A2(new_n300), .A3(new_n476), .A4(new_n481), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n474), .A2(new_n476), .ZN(new_n483));
  AOI21_X1  g297(.A(G902), .B1(new_n455), .B2(G217), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n479), .A2(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G469), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT10), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n259), .A2(KEYINPUT77), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT77), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n209), .A2(new_n489), .A3(KEYINPUT1), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(G128), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n261), .B1(new_n491), .B2(new_n218), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT3), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n411), .B2(G107), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n324), .A2(KEYINPUT3), .A3(G104), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT76), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n497), .B1(new_n324), .B2(G104), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n411), .A2(KEYINPUT76), .A3(G107), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G101), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n496), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n324), .A2(G104), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n411), .A2(G107), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n487), .B1(new_n492), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT78), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g324(.A(KEYINPUT78), .B(new_n487), .C1(new_n492), .C2(new_n507), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n496), .A2(new_n500), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G101), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(KEYINPUT4), .A3(new_n502), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT4), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n513), .A2(new_n516), .A3(G101), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n221), .A3(new_n517), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n494), .A2(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n505), .B1(new_n519), .B2(new_n501), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(KEYINPUT10), .A3(new_n251), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n232), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n512), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT80), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(KEYINPUT12), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(KEYINPUT12), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT79), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n520), .B2(new_n251), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n247), .B1(new_n259), .B2(KEYINPUT77), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n216), .B1(new_n532), .B2(new_n490), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n520), .B1(new_n261), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n507), .A2(KEYINPUT79), .A3(new_n262), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n529), .B1(new_n536), .B2(new_n232), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n200), .A2(G227), .ZN(new_n539));
  XOR2_X1   g353(.A(G110), .B(G140), .Z(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n536), .A2(new_n232), .A3(new_n526), .ZN(new_n543));
  AND4_X1   g357(.A1(new_n524), .A2(new_n538), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT78), .B1(new_n534), .B2(new_n487), .ZN(new_n545));
  INV_X1    g359(.A(new_n511), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n518), .A2(new_n521), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n232), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n542), .B1(new_n549), .B2(new_n524), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n486), .B(new_n300), .C1(new_n544), .C2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n486), .A2(new_n300), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n524), .A2(new_n538), .A3(new_n543), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n541), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n549), .A2(new_n524), .A3(new_n542), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(G469), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n551), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n314), .A2(new_n300), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(G221), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G214), .B1(G237), .B2(G902), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n188), .A2(G952), .ZN(new_n563));
  NAND2_X1  g377(.A1(G234), .A2(G237), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n200), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(G902), .A3(new_n564), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT21), .B(G898), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n515), .A2(new_n275), .A3(new_n517), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n244), .A2(new_n234), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n240), .A2(KEYINPUT5), .A3(new_n242), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n238), .A2(G116), .ZN(new_n576));
  OAI21_X1  g390(.A(G113), .B1(new_n576), .B2(KEYINPUT5), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n520), .A2(new_n574), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(G110), .B(G122), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n573), .A2(new_n580), .A3(new_n582), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(KEYINPUT6), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n215), .A2(new_n217), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n218), .A2(new_n220), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G125), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n249), .B(new_n372), .C1(new_n216), .C2(new_n250), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G224), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(G953), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n592), .B(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT6), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n581), .A2(new_n596), .A3(new_n583), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n586), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n582), .B(KEYINPUT8), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n577), .B1(new_n244), .B2(KEYINPUT5), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n507), .A2(new_n600), .A3(new_n243), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n579), .A2(new_n574), .B1(new_n502), .B2(new_n506), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(KEYINPUT81), .A2(KEYINPUT7), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n591), .B(new_n604), .C1(new_n221), .C2(new_n372), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT7), .B1(new_n593), .B2(G953), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n606), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n590), .A2(new_n591), .A3(new_n608), .A4(new_n604), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n603), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(G902), .B1(new_n610), .B2(new_n585), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n598), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(G210), .B1(G237), .B2(G902), .ZN(new_n613));
  XOR2_X1   g427(.A(new_n613), .B(KEYINPUT83), .Z(new_n614));
  AOI21_X1  g428(.A(new_n612), .B1(KEYINPUT82), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(KEYINPUT82), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n598), .B2(new_n611), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n562), .B(new_n572), .C1(new_n615), .C2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n561), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n311), .A2(new_n454), .A3(new_n485), .A4(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT94), .B(G101), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT95), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n620), .B(new_n622), .ZN(G3));
  INV_X1    g437(.A(KEYINPUT33), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n354), .B2(KEYINPUT96), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n355), .B(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n348), .A2(G902), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n355), .A2(new_n300), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT97), .B(G478), .Z(new_n629));
  AOI22_X1  g443(.A1(new_n626), .A2(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n614), .B1(new_n598), .B2(new_n611), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n598), .A2(new_n611), .A3(new_n614), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n632), .A2(new_n562), .A3(new_n572), .A4(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n446), .B1(new_n433), .B2(new_n437), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n451), .B(new_n449), .C1(new_n635), .C2(new_n422), .ZN(new_n636));
  AOI211_X1 g450(.A(new_n630), .B(new_n634), .C1(new_n636), .C2(new_n421), .ZN(new_n637));
  OAI21_X1  g451(.A(G472), .B1(new_n289), .B2(G902), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n282), .A2(new_n283), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n485), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n561), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  AOI21_X1  g458(.A(new_n436), .B1(new_n445), .B2(new_n435), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n424), .A2(KEYINPUT87), .A3(new_n432), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n439), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n422), .ZN(new_n648));
  INV_X1    g462(.A(new_n633), .ZN(new_n649));
  INV_X1    g463(.A(new_n562), .ZN(new_n650));
  NOR4_X1   g464(.A1(new_n649), .A2(new_n631), .A3(new_n650), .A4(new_n571), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n635), .A2(KEYINPUT20), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n421), .A2(new_n358), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n648), .A2(new_n651), .A3(new_n652), .A4(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT98), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n641), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT35), .B(G107), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  NAND2_X1  g475(.A1(new_n479), .A2(new_n482), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n473), .A2(KEYINPUT36), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(new_n469), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n484), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n638), .A2(new_n639), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n454), .A2(new_n619), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  AOI211_X1 g486(.A(new_n561), .B(new_n667), .C1(new_n309), .C2(new_n310), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n565), .B(KEYINPUT99), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(G900), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n675), .B1(new_n676), .B2(new_n569), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  AND4_X1   g492(.A1(new_n648), .A2(new_n652), .A3(new_n653), .A4(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n632), .A2(new_n562), .A3(new_n633), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(KEYINPUT100), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n648), .A2(new_n652), .A3(new_n653), .A4(new_n678), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n683), .A2(new_n684), .A3(new_n680), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n673), .B1(new_n682), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  INV_X1    g501(.A(new_n561), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n677), .B(KEYINPUT39), .Z(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n690), .B(KEYINPUT40), .Z(new_n691));
  AOI21_X1  g505(.A(new_n207), .B1(new_n298), .B2(new_n256), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n274), .B2(new_n277), .ZN(new_n693));
  OAI21_X1  g507(.A(G472), .B1(new_n693), .B2(G902), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n284), .A2(new_n291), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT101), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n359), .B1(new_n636), .B2(new_n421), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n615), .A2(new_n617), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT38), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n700), .A2(new_n650), .A3(new_n666), .ZN(new_n701));
  AND4_X1   g515(.A1(new_n691), .A2(new_n697), .A3(new_n698), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n210), .ZN(G45));
  OAI21_X1  g517(.A(new_n421), .B1(new_n440), .B2(new_n452), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n626), .A2(new_n627), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n628), .A2(new_n629), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n704), .A2(new_n707), .A3(new_n678), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n667), .B1(new_n309), .B2(new_n310), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n709), .A2(new_n710), .A3(new_n688), .A4(new_n681), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  OAI21_X1  g526(.A(new_n300), .B1(new_n544), .B2(new_n550), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(G469), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n560), .A3(new_n551), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT102), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT102), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n714), .A2(new_n717), .A3(new_n560), .A4(new_n551), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n483), .A2(new_n484), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n662), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n309), .B2(new_n310), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n719), .A2(new_n722), .A3(new_n637), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT41), .B(G113), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  OAI211_X1 g539(.A(new_n722), .B(new_n719), .C1(new_n657), .C2(new_n658), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  NOR3_X1   g541(.A1(new_n715), .A2(new_n571), .A3(new_n680), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n710), .A2(new_n454), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  AOI211_X1 g544(.A(new_n359), .B(new_n680), .C1(new_n636), .C2(new_n421), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n288), .A2(new_n280), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n257), .A2(new_n298), .ZN(new_n733));
  INV_X1    g547(.A(new_n207), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n290), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n638), .A2(KEYINPUT103), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT103), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n738), .B(G472), .C1(new_n289), .C2(G902), .ZN(new_n739));
  AOI211_X1 g553(.A(new_n736), .B(new_n721), .C1(new_n737), .C2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n719), .A2(new_n731), .A3(new_n572), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  INV_X1    g556(.A(new_n736), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n282), .A2(new_n300), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n738), .B1(new_n744), .B2(G472), .ZN(new_n745));
  INV_X1    g559(.A(new_n739), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n666), .B(new_n743), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n551), .ZN(new_n748));
  INV_X1    g562(.A(new_n524), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n523), .B1(new_n512), .B2(new_n522), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n541), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n536), .A2(new_n232), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n537), .B1(new_n753), .B2(new_n526), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n524), .A3(new_n542), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n486), .B1(new_n756), .B2(new_n300), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n748), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n560), .A3(new_n681), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n708), .A2(new_n747), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n372), .ZN(G27));
  NAND2_X1  g575(.A1(new_n555), .A2(KEYINPUT104), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT104), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n554), .A2(new_n763), .A3(new_n541), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n762), .A2(G469), .A3(new_n556), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT105), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n551), .A2(new_n553), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n542), .B1(new_n754), .B2(new_n524), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n749), .A2(new_n750), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n768), .A2(new_n763), .B1(new_n769), .B2(new_n542), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT105), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n770), .A2(new_n771), .A3(G469), .A4(new_n762), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n766), .A2(new_n767), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n560), .A2(new_n562), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n615), .A2(new_n617), .A3(new_n774), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n773), .A2(KEYINPUT106), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT106), .B1(new_n773), .B2(new_n775), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n722), .B(new_n709), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT42), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n773), .A2(new_n775), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT106), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n773), .A2(KEYINPUT106), .A3(new_n775), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n307), .A2(new_n485), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n708), .A2(new_n779), .A3(new_n785), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n778), .A2(new_n779), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n230), .ZN(G33));
  INV_X1    g602(.A(KEYINPUT107), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n683), .B(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n784), .A2(new_n722), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT108), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G134), .ZN(G36));
  NAND2_X1  g607(.A1(new_n668), .A2(new_n666), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT110), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n707), .B(new_n421), .C1(new_n440), .C2(new_n452), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT109), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT43), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n796), .A2(new_n797), .A3(KEYINPUT43), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n795), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT44), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n802), .A2(new_n803), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n770), .A2(KEYINPUT45), .A3(new_n762), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT45), .B1(new_n555), .B2(new_n556), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n486), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n552), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n812), .A2(KEYINPUT46), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n551), .B1(new_n812), .B2(KEYINPUT46), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n560), .B(new_n689), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n699), .A2(new_n562), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n807), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n804), .A2(new_n805), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n806), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G137), .ZN(G39));
  OAI21_X1  g634(.A(new_n560), .B1(new_n813), .B2(new_n814), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT47), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT47), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n823), .B(new_n560), .C1(new_n813), .C2(new_n814), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n311), .A2(new_n708), .A3(new_n485), .A4(new_n816), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G140), .ZN(G42));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n758), .A2(new_n775), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n800), .A2(new_n675), .A3(new_n801), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n785), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n831), .B(KEYINPUT48), .Z(new_n832));
  NAND4_X1  g646(.A1(new_n696), .A2(new_n485), .A3(new_n566), .A4(new_n829), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n630), .B1(new_n636), .B2(new_n421), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n563), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n800), .A2(new_n675), .A3(new_n740), .A4(new_n801), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n759), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n832), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n830), .A2(new_n747), .ZN(new_n842));
  OR3_X1    g656(.A1(new_n833), .A2(new_n704), .A3(new_n707), .ZN(new_n843));
  INV_X1    g657(.A(new_n758), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n560), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n822), .B2(new_n824), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n837), .A2(new_n816), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n842), .B(new_n843), .C1(new_n846), .C2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n700), .A2(new_n650), .A3(new_n560), .A4(new_n758), .ZN(new_n852));
  OR3_X1    g666(.A1(new_n837), .A2(KEYINPUT117), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT117), .B1(new_n837), .B2(new_n852), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(KEYINPUT118), .B(KEYINPUT50), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n837), .A2(new_n852), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT50), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n841), .B1(new_n851), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n849), .B1(new_n860), .B2(KEYINPUT119), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n855), .A2(new_n856), .B1(KEYINPUT50), .B2(new_n858), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT119), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT51), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n828), .B1(new_n862), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n849), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n864), .B2(new_n865), .ZN(new_n870));
  INV_X1    g684(.A(new_n866), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n850), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n872), .A2(new_n861), .A3(KEYINPUT120), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n708), .A2(new_n747), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n776), .B2(new_n777), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT113), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n816), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n635), .A2(KEYINPUT20), .ZN(new_n880));
  AOI211_X1 g694(.A(new_n422), .B(new_n446), .C1(new_n433), .C2(new_n437), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n358), .B(KEYINPUT112), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n677), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n421), .A2(new_n879), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n673), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n875), .B(KEYINPUT113), .C1(new_n777), .C2(new_n776), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n878), .A2(new_n791), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n561), .A2(new_n640), .A3(new_n618), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n636), .A2(new_n883), .A3(new_n421), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n891), .B2(new_n834), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n892), .A2(new_n620), .A3(new_n670), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n716), .A2(new_n572), .A3(new_n718), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n485), .B(new_n743), .C1(new_n745), .C2(new_n746), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n759), .A2(new_n453), .A3(new_n571), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n896), .A2(new_n731), .B1(new_n897), .B2(new_n710), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n893), .A2(new_n898), .A3(new_n723), .A4(new_n726), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n888), .A2(new_n899), .A3(new_n787), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n875), .A2(new_n839), .ZN(new_n901));
  AND4_X1   g715(.A1(new_n560), .A2(new_n695), .A3(new_n667), .A4(new_n678), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n731), .A2(new_n902), .A3(new_n773), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n686), .A2(new_n711), .A3(new_n901), .A4(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT52), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n684), .B1(new_n683), .B2(new_n680), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n421), .A2(new_n358), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n880), .A2(new_n881), .A3(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(KEYINPUT100), .A3(new_n681), .A4(new_n678), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n760), .B1(new_n673), .B2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n912), .A2(KEYINPUT52), .A3(new_n711), .A4(new_n903), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n906), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT53), .B1(new_n900), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n741), .A2(new_n723), .A3(new_n729), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n882), .A2(KEYINPUT98), .A3(new_n651), .A4(new_n653), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n656), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n719), .A2(new_n722), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT115), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT115), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n898), .A2(new_n922), .A3(new_n726), .A4(new_n723), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n892), .A2(new_n620), .A3(KEYINPUT53), .A4(new_n670), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n888), .A2(new_n787), .A3(new_n925), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n906), .A2(KEYINPUT114), .A3(new_n913), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT114), .B1(new_n906), .B2(new_n913), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n924), .B(new_n926), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT116), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n915), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT54), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT114), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n914), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n906), .A2(new_n913), .A3(KEYINPUT114), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n936), .A2(KEYINPUT116), .A3(new_n924), .A4(new_n926), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n931), .A2(new_n932), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT53), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n900), .B2(new_n914), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n722), .B1(new_n776), .B2(new_n777), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n683), .B(KEYINPUT107), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n886), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n887), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT113), .B1(new_n784), .B2(new_n875), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n899), .ZN(new_n947));
  INV_X1    g761(.A(new_n787), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n949), .A2(KEYINPUT53), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n940), .B1(new_n936), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT54), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n938), .A2(new_n952), .ZN(new_n953));
  OAI22_X1  g767(.A1(new_n874), .A2(new_n953), .B1(G952), .B2(G953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n700), .A2(new_n485), .A3(new_n562), .A4(new_n560), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n758), .B(KEYINPUT49), .Z(new_n956));
  OR4_X1    g770(.A1(new_n697), .A2(new_n955), .A3(new_n956), .A4(new_n796), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n954), .A2(new_n957), .ZN(G75));
  INV_X1    g772(.A(new_n914), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n939), .B1(new_n949), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n787), .A2(new_n925), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n924), .A2(new_n946), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n934), .B2(new_n935), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n960), .B1(new_n963), .B2(KEYINPUT116), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n929), .A2(new_n930), .ZN(new_n965));
  OAI211_X1 g779(.A(G902), .B(new_n614), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT121), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n300), .B1(new_n931), .B2(new_n937), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n969), .A2(KEYINPUT121), .A3(new_n614), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n586), .A2(new_n597), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(new_n595), .Z(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT55), .ZN(new_n973));
  XNOR2_X1  g787(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n968), .A2(new_n970), .A3(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n200), .A2(G952), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(KEYINPUT56), .B1(new_n969), .B2(new_n614), .ZN(new_n979));
  INV_X1    g793(.A(new_n973), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n976), .A2(new_n981), .ZN(G51));
  INV_X1    g796(.A(KEYINPUT123), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n929), .A2(new_n930), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n984), .A2(new_n937), .A3(new_n960), .ZN(new_n985));
  AND4_X1   g799(.A1(new_n983), .A2(new_n985), .A3(G902), .A4(new_n811), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n983), .B1(new_n969), .B2(new_n811), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n552), .B(KEYINPUT57), .ZN(new_n989));
  AND4_X1   g803(.A1(new_n932), .A2(new_n984), .A3(new_n937), .A4(new_n960), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n932), .B1(new_n931), .B2(new_n937), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n756), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n977), .B1(new_n988), .B2(new_n993), .ZN(G54));
  AND2_X1   g808(.A1(KEYINPUT58), .A2(G475), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n969), .A2(new_n438), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n438), .B1(new_n969), .B2(new_n995), .ZN(new_n997));
  NOR3_X1   g811(.A1(new_n996), .A2(new_n997), .A3(new_n977), .ZN(G60));
  NAND2_X1  g812(.A1(G478), .A2(G902), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT59), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n626), .B1(new_n953), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n626), .A2(new_n1000), .ZN(new_n1002));
  INV_X1    g816(.A(new_n991), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1002), .B1(new_n1003), .B2(new_n938), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n1001), .A2(new_n1004), .A3(new_n977), .ZN(G63));
  INV_X1    g819(.A(KEYINPUT61), .ZN(new_n1006));
  NAND2_X1  g820(.A1(G217), .A2(G902), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT60), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1008), .B1(new_n931), .B2(new_n937), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n664), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n978), .B1(new_n1009), .B2(new_n483), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1006), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OR2_X1    g827(.A1(new_n1009), .A2(new_n483), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1014), .A2(KEYINPUT61), .A3(new_n978), .A4(new_n1010), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1013), .A2(new_n1015), .ZN(G66));
  OAI21_X1  g830(.A(G953), .B1(new_n570), .B2(new_n593), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1017), .B1(new_n947), .B2(new_n567), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n971), .B1(G898), .B2(new_n200), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1018), .B(new_n1019), .ZN(G69));
  INV_X1    g834(.A(KEYINPUT62), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n912), .A2(new_n711), .ZN(new_n1022));
  OR3_X1    g836(.A1(new_n702), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1021), .B1(new_n702), .B2(new_n1022), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n826), .ZN(new_n1026));
  AOI211_X1 g840(.A(new_n816), .B(new_n690), .C1(new_n835), .C2(new_n890), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1026), .B1(new_n722), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1025), .A2(new_n819), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n276), .B1(new_n266), .B2(KEYINPUT30), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n1030), .B(KEYINPUT124), .Z(new_n1031));
  XOR2_X1   g845(.A(new_n1031), .B(new_n429), .Z(new_n1032));
  NAND3_X1  g846(.A1(new_n1029), .A2(new_n200), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n731), .A2(new_n307), .A3(new_n485), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n791), .B1(new_n815), .B2(new_n1034), .ZN(new_n1035));
  NOR3_X1   g849(.A1(new_n1026), .A2(new_n1022), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1036), .A2(new_n948), .A3(new_n819), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(new_n200), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1032), .B1(new_n676), .B2(new_n567), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT125), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n200), .B1(G227), .B2(G900), .ZN(new_n1042));
  OAI211_X1 g856(.A(new_n1033), .B(new_n1040), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1042), .A2(new_n1041), .ZN(new_n1044));
  XNOR2_X1  g858(.A(new_n1043), .B(new_n1044), .ZN(G72));
  NAND2_X1  g859(.A1(G472), .A2(G902), .ZN(new_n1046));
  XOR2_X1   g860(.A(new_n1046), .B(KEYINPUT63), .Z(new_n1047));
  OAI21_X1  g861(.A(new_n1047), .B1(new_n1037), .B2(new_n899), .ZN(new_n1048));
  AND3_X1   g862(.A1(new_n277), .A2(new_n256), .A3(new_n734), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n977), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g864(.A1(new_n1025), .A2(new_n819), .A3(new_n947), .A4(new_n1028), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1051), .A2(new_n1047), .ZN(new_n1052));
  INV_X1    g866(.A(KEYINPUT126), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n734), .B1(new_n277), .B2(new_n256), .ZN(new_n1054));
  AND3_X1   g868(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g869(.A(new_n1053), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n1050), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g871(.A(new_n304), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1058), .A2(new_n286), .ZN(new_n1059));
  NAND3_X1  g873(.A1(new_n951), .A2(new_n1047), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1060), .A2(KEYINPUT127), .ZN(new_n1061));
  OR2_X1    g875(.A1(new_n1060), .A2(KEYINPUT127), .ZN(new_n1062));
  AOI21_X1  g876(.A(new_n1057), .B1(new_n1061), .B2(new_n1062), .ZN(G57));
endmodule


