//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT81), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(KEYINPUT64), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n190), .B1(new_n194), .B2(G143), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT68), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n190), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G146), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n200), .B(new_n198), .C1(new_n201), .C2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT68), .ZN(new_n204));
  INV_X1    g018(.A(new_n195), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n189), .A2(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G128), .ZN(new_n208));
  AOI22_X1  g022(.A1(new_n199), .A2(new_n204), .B1(new_n205), .B2(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(G104), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n213), .A2(G107), .B1(KEYINPUT79), .B2(KEYINPUT3), .ZN(new_n214));
  OAI22_X1  g028(.A1(new_n213), .A2(G107), .B1(KEYINPUT79), .B2(KEYINPUT3), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n212), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  OR2_X1    g030(.A1(new_n216), .A2(G101), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n211), .A2(G104), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n213), .A2(G107), .ZN(new_n219));
  OAI21_X1  g033(.A(G101), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n188), .B1(new_n209), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n205), .A2(new_n208), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n196), .B1(new_n195), .B2(new_n198), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n203), .A2(KEYINPUT68), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n217), .A2(new_n220), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(KEYINPUT81), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT10), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n202), .B1(new_n191), .B2(new_n193), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT1), .ZN(new_n231));
  OAI21_X1  g045(.A(G128), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n206), .B1(new_n194), .B2(G143), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n234), .B1(new_n224), .B2(new_n225), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(KEYINPUT10), .A3(new_n227), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n216), .A2(new_n237), .A3(G101), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT80), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n238), .B(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n237), .B1(new_n216), .B2(G101), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n217), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n233), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n195), .A2(new_n244), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n236), .B1(new_n243), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT65), .B(KEYINPUT11), .ZN(new_n252));
  INV_X1    g066(.A(G134), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(G137), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT66), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT11), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT65), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT65), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT11), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n261));
  INV_X1    g075(.A(G137), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G134), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n255), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n262), .A2(G134), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n262), .A2(KEYINPUT11), .A3(G134), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT67), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n262), .A2(KEYINPUT67), .A3(KEYINPUT11), .A4(G134), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G131), .ZN(new_n273));
  INV_X1    g087(.A(G131), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n252), .A2(KEYINPUT66), .A3(new_n254), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n261), .B1(new_n260), .B2(new_n263), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n274), .B(new_n271), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  NOR3_X1   g092(.A1(new_n229), .A2(new_n251), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(G110), .B(G140), .ZN(new_n280));
  INV_X1    g094(.A(G953), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n281), .A2(G227), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n280), .B(new_n282), .Z(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n187), .B1(new_n279), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n222), .A2(new_n228), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT10), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n278), .ZN(new_n289));
  OR2_X1    g103(.A1(new_n238), .A2(new_n239), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n238), .A2(new_n239), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n290), .A2(new_n291), .B1(new_n217), .B2(new_n241), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n249), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n288), .A2(new_n289), .A3(new_n293), .A4(new_n236), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(KEYINPUT82), .A3(new_n283), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n199), .A2(new_n204), .B1(new_n233), .B2(new_n232), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n222), .A2(new_n228), .B1(new_n296), .B2(new_n221), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(KEYINPUT12), .A3(new_n278), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT12), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n297), .B2(new_n289), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n285), .A2(new_n295), .A3(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n229), .A2(new_n251), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(new_n289), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n284), .B1(new_n305), .B2(new_n279), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G469), .ZN(new_n308));
  INV_X1    g122(.A(G902), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  OR3_X1    g124(.A1(new_n305), .A2(new_n279), .A3(new_n284), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n279), .B1(new_n299), .B2(new_n301), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n311), .B(G469), .C1(new_n312), .C2(new_n283), .ZN(new_n313));
  NAND2_X1  g127(.A1(G469), .A2(G902), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  XOR2_X1   g129(.A(KEYINPUT9), .B(G234), .Z(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G221), .B1(new_n317), .B2(G902), .ZN(new_n318));
  XOR2_X1   g132(.A(new_n318), .B(KEYINPUT78), .Z(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  XOR2_X1   g135(.A(G110), .B(G122), .Z(new_n322));
  XOR2_X1   g136(.A(G116), .B(G119), .Z(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT2), .B(G113), .ZN(new_n324));
  XOR2_X1   g138(.A(new_n323), .B(new_n324), .Z(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n240), .A2(new_n326), .A3(new_n242), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT5), .ZN(new_n328));
  INV_X1    g142(.A(G119), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(G116), .ZN(new_n330));
  OAI211_X1 g144(.A(G113), .B(new_n330), .C1(new_n323), .C2(new_n328), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n323), .B2(new_n324), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n221), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n322), .B1(new_n327), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n322), .ZN(new_n335));
  INV_X1    g149(.A(new_n333), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n335), .B(new_n336), .C1(new_n243), .C2(new_n325), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(KEYINPUT6), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT74), .B(G125), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n249), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n296), .B2(new_n339), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n281), .A2(G224), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT83), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n341), .B(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT6), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n345), .B(new_n322), .C1(new_n327), .C2(new_n333), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n338), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n342), .A2(KEYINPUT7), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n341), .B(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT84), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n221), .A2(new_n332), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n336), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  XOR2_X1   g166(.A(new_n322), .B(KEYINPUT8), .Z(new_n353));
  NAND3_X1  g167(.A1(new_n221), .A2(KEYINPUT84), .A3(new_n332), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n349), .A2(new_n355), .A3(new_n337), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n347), .A2(new_n309), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(G210), .B1(G237), .B2(G902), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n347), .A2(new_n356), .A3(new_n309), .A4(new_n358), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(KEYINPUT85), .A3(new_n361), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n347), .A2(new_n309), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT85), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n363), .A2(new_n364), .A3(new_n358), .A4(new_n356), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(G214), .B1(G237), .B2(G902), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  XOR2_X1   g183(.A(KEYINPUT89), .B(KEYINPUT13), .Z(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(G128), .A3(new_n202), .ZN(new_n371));
  XOR2_X1   g185(.A(G128), .B(G143), .Z(new_n372));
  OAI211_X1 g186(.A(new_n371), .B(G134), .C1(new_n372), .C2(new_n370), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n372), .A2(G134), .ZN(new_n374));
  XNOR2_X1  g188(.A(G116), .B(G122), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(new_n211), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT14), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G116), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(KEYINPUT14), .A3(G122), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(G107), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(KEYINPUT90), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n372), .A2(G134), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n374), .A2(new_n384), .B1(new_n211), .B2(new_n375), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n383), .A2(KEYINPUT91), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(KEYINPUT91), .B1(new_n383), .B2(new_n385), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n377), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G217), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n317), .A2(new_n389), .A3(G953), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n377), .B(new_n390), .C1(new_n386), .C2(new_n387), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(KEYINPUT92), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT92), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n388), .A2(new_n395), .A3(new_n391), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n394), .A2(KEYINPUT93), .A3(new_n309), .A4(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G478), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(KEYINPUT15), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n397), .A2(new_n399), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n281), .A2(G952), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(G234), .B2(G237), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  XOR2_X1   g219(.A(KEYINPUT21), .B(G898), .Z(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(KEYINPUT94), .ZN(new_n407));
  AOI211_X1 g221(.A(new_n309), .B(new_n281), .C1(G234), .C2(G237), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n405), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(G125), .A2(G140), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(new_n339), .B2(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G146), .ZN(new_n413));
  XNOR2_X1  g227(.A(G125), .B(G140), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n194), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G237), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(new_n281), .A3(G214), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(G143), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(KEYINPUT18), .A2(G131), .ZN(new_n421));
  XOR2_X1   g235(.A(new_n421), .B(KEYINPUT87), .Z(new_n422));
  XOR2_X1   g236(.A(new_n419), .B(KEYINPUT86), .Z(new_n423));
  OAI221_X1 g237(.A(new_n416), .B1(new_n420), .B2(new_n422), .C1(new_n423), .C2(new_n421), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT16), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n339), .A2(new_n425), .ZN(new_n426));
  OAI22_X1  g240(.A1(new_n412), .A2(new_n425), .B1(new_n426), .B2(G140), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n427), .A2(new_n189), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n419), .B(new_n274), .ZN(new_n429));
  MUX2_X1   g243(.A(new_n414), .B(new_n412), .S(KEYINPUT19), .Z(new_n430));
  OAI211_X1 g244(.A(new_n428), .B(new_n429), .C1(new_n201), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n424), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G113), .B(G122), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(new_n213), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n427), .B(new_n189), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n420), .A2(KEYINPUT17), .A3(G131), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n438), .B(new_n439), .C1(KEYINPUT17), .C2(new_n429), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(new_n434), .A3(new_n424), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G475), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n443), .A3(new_n309), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT20), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n442), .A2(new_n446), .A3(new_n443), .A4(new_n309), .ZN(new_n447));
  INV_X1    g261(.A(new_n441), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n434), .B1(new_n424), .B2(new_n440), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n309), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT88), .B(G475), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n445), .A2(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n402), .A2(new_n410), .A3(new_n452), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n321), .A2(new_n369), .A3(new_n453), .ZN(new_n454));
  XOR2_X1   g268(.A(KEYINPUT26), .B(KEYINPUT27), .Z(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(G101), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n417), .A2(new_n281), .A3(G210), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n456), .B(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(G131), .B1(new_n254), .B2(new_n266), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n277), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT69), .B1(new_n462), .B2(new_n296), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT69), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n235), .A2(new_n464), .A3(new_n277), .A4(new_n461), .ZN(new_n465));
  INV_X1    g279(.A(new_n277), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n274), .B1(new_n265), .B2(new_n271), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n249), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n463), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT30), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n277), .A2(new_n461), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n278), .A2(new_n249), .B1(new_n472), .B2(new_n235), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT30), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n326), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n235), .A2(new_n277), .A3(new_n461), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(new_n468), .A3(new_n325), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT70), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT70), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n476), .A2(new_n468), .A3(new_n479), .A4(new_n325), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n460), .B1(new_n475), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT28), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n478), .A2(new_n480), .B1(new_n326), .B2(new_n469), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n484), .B1(new_n485), .B2(new_n483), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n459), .B(KEYINPUT72), .ZN(new_n488));
  AOI211_X1 g302(.A(KEYINPUT29), .B(new_n482), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n473), .A2(new_n325), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(new_n478), .B2(new_n480), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n484), .B1(new_n491), .B2(new_n483), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n460), .A2(KEYINPUT29), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n309), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G472), .B1(new_n489), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(G472), .A2(G902), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n479), .B1(new_n473), .B2(new_n325), .ZN(new_n498));
  INV_X1    g312(.A(new_n480), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n460), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT71), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n481), .A2(KEYINPUT71), .A3(new_n460), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n475), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n488), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n504), .A2(KEYINPUT31), .B1(new_n486), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT31), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n502), .A2(new_n507), .A3(new_n475), .A4(new_n503), .ZN(new_n508));
  AOI211_X1 g322(.A(KEYINPUT32), .B(new_n497), .C1(new_n506), .C2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT32), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n504), .A2(KEYINPUT31), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n486), .A2(new_n505), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n510), .B1(new_n513), .B2(new_n496), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n495), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT73), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT23), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n517), .B1(G119), .B2(new_n197), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n329), .A2(KEYINPUT23), .A3(G128), .ZN(new_n519));
  OAI22_X1  g333(.A1(new_n518), .A2(new_n519), .B1(G119), .B2(new_n197), .ZN(new_n520));
  XNOR2_X1  g334(.A(G119), .B(G128), .ZN(new_n521));
  XOR2_X1   g335(.A(KEYINPUT24), .B(G110), .Z(new_n522));
  AOI22_X1  g336(.A1(new_n520), .A2(G110), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n437), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT75), .B(G110), .ZN(new_n525));
  OAI22_X1  g339(.A1(new_n520), .A2(new_n525), .B1(new_n521), .B2(new_n522), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n428), .A2(new_n415), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n281), .A2(G221), .A3(G234), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(KEYINPUT22), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(G137), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT76), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n524), .A2(KEYINPUT76), .A3(new_n527), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n533), .B1(new_n537), .B2(new_n532), .ZN(new_n538));
  OR2_X1    g352(.A1(new_n538), .A2(KEYINPUT77), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(KEYINPUT77), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n389), .B1(G234), .B2(new_n309), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(G902), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n538), .ZN(new_n546));
  OR3_X1    g360(.A1(new_n546), .A2(KEYINPUT25), .A3(G902), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT25), .B1(new_n546), .B2(G902), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n543), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT73), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n552), .B(new_n495), .C1(new_n509), .C2(new_n514), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n454), .A2(new_n516), .A3(new_n551), .A4(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(G101), .ZN(G3));
  OR2_X1    g369(.A1(new_n360), .A2(KEYINPUT95), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n360), .A2(KEYINPUT95), .A3(new_n361), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n556), .A2(new_n367), .A3(new_n410), .A4(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n394), .A2(new_n396), .ZN(new_n560));
  AOI21_X1  g374(.A(G478), .B1(new_n560), .B2(new_n309), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n392), .A2(KEYINPUT33), .A3(new_n393), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT33), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n394), .A2(new_n563), .A3(new_n396), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n394), .A2(KEYINPUT96), .A3(new_n563), .A4(new_n396), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n562), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n398), .A2(G902), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n561), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(new_n452), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n559), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT97), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n559), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n513), .A2(new_n309), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G472), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT71), .B1(new_n481), .B2(new_n460), .ZN(new_n580));
  AOI211_X1 g394(.A(new_n501), .B(new_n459), .C1(new_n478), .C2(new_n480), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n471), .A2(new_n326), .A3(new_n474), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n512), .B1(new_n583), .B2(new_n507), .ZN(new_n584));
  INV_X1    g398(.A(new_n508), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n496), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n579), .A2(new_n586), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n587), .A2(new_n550), .A3(new_n319), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n315), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n577), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT34), .B(G104), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G6));
  OAI21_X1  g406(.A(new_n452), .B1(new_n400), .B2(new_n401), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n558), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT35), .B(G107), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G9));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n532), .A2(KEYINPUT36), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n537), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n544), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n549), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n599), .B1(new_n587), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n579), .A2(KEYINPUT98), .A3(new_n603), .A4(new_n586), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n454), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT37), .ZN(new_n608));
  XOR2_X1   g422(.A(new_n608), .B(G110), .Z(G12));
  AND3_X1   g423(.A1(new_n556), .A2(new_n367), .A3(new_n557), .ZN(new_n610));
  AND4_X1   g424(.A1(new_n516), .A2(new_n553), .A3(new_n610), .A4(new_n603), .ZN(new_n611));
  INV_X1    g425(.A(G900), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n404), .B1(new_n408), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n593), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n611), .A2(new_n321), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G128), .ZN(G30));
  XOR2_X1   g430(.A(new_n613), .B(KEYINPUT39), .Z(new_n617));
  NAND2_X1  g431(.A1(new_n321), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n618), .B(KEYINPUT40), .Z(new_n619));
  XOR2_X1   g433(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n366), .B(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n402), .A2(new_n452), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n603), .A2(new_n368), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n504), .B(G472), .C1(new_n488), .C2(new_n491), .ZN(new_n625));
  NAND2_X1  g439(.A1(G472), .A2(G902), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT100), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n586), .A2(KEYINPUT32), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n513), .A2(new_n510), .A3(new_n496), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n619), .A2(new_n623), .A3(new_n624), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G143), .ZN(G45));
  INV_X1    g448(.A(new_n613), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n571), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n611), .A2(new_n321), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G146), .ZN(G48));
  NAND2_X1  g453(.A1(new_n307), .A2(new_n309), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(G469), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n641), .A2(KEYINPUT101), .A3(new_n310), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n640), .A2(new_n643), .A3(G469), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n319), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n516), .A2(new_n551), .A3(new_n553), .A4(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n577), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT41), .B(G113), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G15));
  NOR2_X1   g463(.A1(new_n646), .A2(new_n595), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(new_n380), .ZN(G18));
  AOI21_X1  g465(.A(KEYINPUT102), .B1(new_n645), .B2(new_n610), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n645), .A2(KEYINPUT102), .A3(new_n610), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n516), .A2(new_n553), .A3(new_n453), .A4(new_n603), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G119), .ZN(G21));
  NAND2_X1  g473(.A1(new_n492), .A2(new_n505), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n511), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT103), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n511), .A2(new_n663), .A3(new_n660), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n662), .A2(new_n508), .A3(new_n664), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n665), .A2(new_n496), .B1(G472), .B2(new_n578), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n666), .A2(new_n645), .A3(new_n551), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n558), .A2(new_n402), .A3(new_n452), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n666), .A2(new_n645), .A3(new_n669), .A4(new_n551), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT104), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G122), .ZN(G24));
  INV_X1    g488(.A(new_n666), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n675), .A2(new_n636), .A3(new_n604), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n655), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G125), .ZN(G27));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(new_n366), .B2(new_n367), .ZN(new_n680));
  AOI211_X1 g494(.A(KEYINPUT106), .B(new_n368), .C1(new_n362), .C2(new_n365), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n636), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n314), .B(KEYINPUT105), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n313), .A2(new_n685), .ZN(new_n686));
  AOI211_X1 g500(.A(G469), .B(G902), .C1(new_n303), .C2(new_n306), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n320), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n550), .B1(new_n631), .B2(new_n495), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n684), .A2(KEYINPUT42), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n552), .B1(new_n631), .B2(new_n495), .ZN(new_n693));
  INV_X1    g507(.A(new_n553), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n680), .A2(new_n681), .A3(new_n688), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n695), .A2(new_n551), .A3(new_n637), .A4(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT42), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n692), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n516), .A2(new_n696), .A3(new_n551), .A4(new_n553), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n692), .B(new_n698), .C1(new_n700), .C2(new_n636), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n691), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G131), .ZN(G33));
  INV_X1    g518(.A(new_n614), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n253), .ZN(G36));
  INV_X1    g521(.A(new_n570), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n452), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n708), .A2(KEYINPUT43), .A3(new_n452), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n587), .A3(new_n603), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n713), .A2(KEYINPUT44), .A3(new_n587), .A4(new_n603), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n682), .A3(new_n717), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n718), .A2(KEYINPUT109), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n311), .B1(new_n312), .B2(new_n283), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(G469), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n685), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT46), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT108), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n724), .A2(KEYINPUT46), .A3(new_n685), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n725), .A2(new_n730), .A3(new_n726), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n728), .A2(new_n310), .A3(new_n729), .A4(new_n731), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n732), .A2(new_n320), .A3(new_n617), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n718), .A2(KEYINPUT109), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n719), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G137), .ZN(G39));
  INV_X1    g550(.A(KEYINPUT47), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(KEYINPUT110), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n732), .B2(new_n320), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n732), .A2(new_n320), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n737), .A2(KEYINPUT110), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n740), .B1(new_n743), .B2(new_n739), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n516), .A2(new_n553), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n684), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(new_n550), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G140), .ZN(G42));
  OR2_X1    g562(.A1(G952), .A2(G953), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n698), .B1(new_n700), .B2(new_n636), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT107), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n701), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n706), .B1(new_n753), .B2(new_n691), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n402), .A2(new_n452), .A3(new_n635), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n683), .B1(new_n756), .B2(KEYINPUT114), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n757), .A2(new_n321), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n756), .A2(KEYINPUT114), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n745), .A2(new_n604), .A3(new_n759), .ZN(new_n760));
  AOI22_X1  g574(.A1(new_n758), .A2(new_n760), .B1(new_n676), .B2(new_n696), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n611), .B(new_n321), .C1(new_n614), .C2(new_n637), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n610), .A2(new_n622), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n603), .A2(new_n613), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n632), .A2(new_n689), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n762), .A2(new_n677), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT52), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n762), .A2(new_n768), .A3(new_n677), .A4(new_n765), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n754), .A2(new_n761), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n593), .B1(new_n570), .B2(new_n452), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n771), .A2(new_n369), .A3(new_n410), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n588), .A2(new_n772), .A3(new_n315), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n554), .A2(new_n773), .A3(new_n607), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT113), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n650), .B1(new_n670), .B2(new_n672), .ZN(new_n777));
  INV_X1    g591(.A(new_n646), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n655), .A2(new_n657), .B1(new_n778), .B2(new_n576), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n777), .A2(KEYINPUT112), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT112), .B1(new_n777), .B2(new_n779), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n750), .B1(new_n770), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n706), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n703), .A2(new_n784), .A3(new_n761), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n767), .A2(new_n769), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n654), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n652), .ZN(new_n789));
  OAI22_X1  g603(.A1(new_n789), .A2(new_n656), .B1(new_n577), .B2(new_n646), .ZN(new_n790));
  INV_X1    g604(.A(new_n650), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n673), .A2(new_n791), .ZN(new_n792));
  NOR4_X1   g606(.A1(new_n775), .A2(new_n750), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n787), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n783), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(KEYINPUT54), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT115), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n798));
  INV_X1    g612(.A(new_n781), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n777), .A2(new_n779), .A3(KEYINPUT112), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n775), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n787), .A2(new_n801), .A3(KEYINPUT53), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n783), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n798), .B1(new_n803), .B2(KEYINPUT54), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n797), .B1(new_n796), .B2(new_n804), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n403), .B(KEYINPUT118), .Z(new_n806));
  OR2_X1    g620(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n807));
  NAND2_X1  g621(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n713), .A2(KEYINPUT116), .A3(new_n404), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT116), .B1(new_n713), .B2(new_n404), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n368), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n667), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n812), .A2(new_n621), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n807), .B(new_n808), .C1(new_n811), .C2(new_n813), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n809), .A2(new_n810), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n682), .A2(new_n645), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n815), .A2(new_n603), .A3(new_n666), .A4(new_n817), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n816), .A2(new_n632), .A3(new_n550), .A4(new_n405), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n452), .A3(new_n570), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n814), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n815), .A2(new_n551), .A3(new_n666), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n642), .A2(new_n644), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n319), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n822), .B(new_n682), .C1(new_n744), .C2(new_n825), .ZN(new_n826));
  OR3_X1    g640(.A1(new_n811), .A2(new_n813), .A3(new_n807), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n821), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n821), .A2(new_n826), .A3(KEYINPUT51), .A4(new_n827), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n822), .A2(new_n655), .ZN(new_n832));
  AND4_X1   g646(.A1(new_n806), .A2(new_n830), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n815), .A2(new_n690), .A3(new_n817), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT48), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n819), .A2(new_n571), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n749), .B1(new_n805), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n551), .A2(new_n320), .A3(new_n367), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT111), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n632), .A2(new_n621), .A3(new_n709), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n823), .B(KEYINPUT49), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n838), .A2(new_n843), .ZN(G75));
  NAND3_X1  g658(.A1(new_n795), .A2(G210), .A3(G902), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT56), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n338), .A2(new_n346), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(new_n344), .ZN(new_n849));
  XOR2_X1   g663(.A(new_n849), .B(KEYINPUT55), .Z(new_n850));
  NAND2_X1  g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n281), .A2(G952), .ZN(new_n854));
  XNOR2_X1  g668(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n854), .B1(new_n845), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n847), .A2(KEYINPUT119), .A3(new_n850), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n853), .A2(new_n857), .A3(new_n858), .ZN(G51));
  NAND2_X1  g673(.A1(new_n685), .A2(KEYINPUT57), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n783), .B2(new_n794), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n860), .B1(new_n796), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n685), .A2(KEYINPUT57), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n307), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n795), .A2(G902), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n866), .A2(new_n724), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n854), .B1(new_n865), .B2(new_n867), .ZN(G54));
  NAND4_X1  g682(.A1(new_n795), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n869));
  INV_X1    g683(.A(new_n442), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n871), .A2(new_n872), .A3(new_n854), .ZN(G60));
  NAND2_X1  g687(.A1(G478), .A2(G902), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT59), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n568), .B(KEYINPUT121), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n875), .B(new_n877), .C1(new_n796), .C2(new_n862), .ZN(new_n878));
  INV_X1    g692(.A(new_n854), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n805), .A2(new_n875), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n880), .B1(new_n881), .B2(new_n876), .ZN(G63));
  INV_X1    g696(.A(KEYINPUT61), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(KEYINPUT125), .ZN(new_n884));
  XOR2_X1   g698(.A(KEYINPUT122), .B(KEYINPUT60), .Z(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT123), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n389), .A2(new_n309), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n886), .B(new_n887), .Z(new_n888));
  AOI21_X1  g702(.A(KEYINPUT53), .B1(new_n787), .B2(new_n801), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n776), .A2(KEYINPUT53), .A3(new_n779), .A4(new_n777), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(new_n770), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n601), .B(new_n888), .C1(new_n889), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT124), .ZN(new_n893));
  INV_X1    g707(.A(new_n888), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n783), .B2(new_n794), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n896), .A3(new_n601), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n883), .A2(KEYINPUT125), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n879), .B(new_n899), .C1(new_n895), .C2(new_n542), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n884), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n900), .ZN(new_n902));
  INV_X1    g716(.A(new_n884), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n902), .A2(new_n903), .A3(new_n893), .A4(new_n897), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n901), .A2(new_n904), .ZN(G66));
  NAND2_X1  g719(.A1(new_n407), .A2(G224), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(G953), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n907), .B1(new_n801), .B2(G953), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n848), .B1(G898), .B2(new_n281), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n908), .B(new_n909), .ZN(G69));
  AND2_X1   g724(.A1(new_n747), .A2(new_n735), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n762), .A2(new_n677), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n733), .A2(new_n690), .A3(new_n763), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n911), .A2(new_n754), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n281), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n612), .A2(G953), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT127), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n471), .A2(new_n474), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n430), .B(KEYINPUT126), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n921), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n912), .A2(new_n633), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n683), .A2(new_n618), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n695), .A2(new_n927), .A3(new_n551), .A4(new_n771), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n926), .A2(new_n911), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n923), .B1(new_n929), .B2(G953), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n922), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n281), .B1(G227), .B2(G900), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(G72));
  NAND2_X1  g747(.A1(new_n475), .A2(new_n481), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n929), .A2(new_n801), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n626), .B(KEYINPUT63), .Z(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n460), .B(new_n934), .C1(new_n935), .C2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n936), .B1(new_n914), .B2(new_n782), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n939), .A2(new_n475), .A3(new_n481), .A4(new_n459), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n803), .B(new_n936), .C1(new_n583), .C2(new_n482), .ZN(new_n941));
  AND4_X1   g755(.A1(new_n879), .A2(new_n938), .A3(new_n940), .A4(new_n941), .ZN(G57));
endmodule


