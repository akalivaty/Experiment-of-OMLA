//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G122), .ZN(new_n188));
  XNOR2_X1  g002(.A(G116), .B(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT2), .A2(G113), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT67), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT67), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT2), .A3(G113), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  OR2_X1    g008(.A1(KEYINPUT2), .A2(G113), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n189), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n195), .A3(new_n189), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G104), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(new_n200), .B2(G107), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G104), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(G107), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G101), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n201), .A2(new_n204), .A3(new_n208), .A4(new_n205), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(KEYINPUT4), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT4), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n206), .A2(new_n211), .A3(G101), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n199), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n200), .A2(G107), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n203), .A2(G104), .ZN(new_n215));
  OAI21_X1  g029(.A(G101), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n209), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G119), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G116), .ZN(new_n219));
  INV_X1    g033(.A(G116), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G119), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT5), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT5), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n218), .A3(G116), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G113), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT80), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT5), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT80), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n227), .A2(new_n228), .A3(G113), .A4(new_n224), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n217), .A2(new_n226), .A3(new_n198), .A4(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n188), .B1(new_n213), .B2(new_n230), .ZN(new_n231));
  OR2_X1    g045(.A1(new_n231), .A2(KEYINPUT6), .ZN(new_n232));
  INV_X1    g046(.A(new_n198), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n212), .B1(new_n233), .B2(new_n196), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n207), .A2(KEYINPUT4), .A3(new_n209), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n230), .B(new_n188), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT81), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT81), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n213), .A2(new_n238), .A3(new_n188), .A4(new_n230), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n231), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT6), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n232), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G146), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G143), .ZN(new_n244));
  INV_X1    g058(.A(G143), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT1), .B1(new_n245), .B2(G146), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(G128), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G128), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n244), .B(new_n246), .C1(KEYINPUT1), .C2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(G125), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G125), .ZN(new_n254));
  AND2_X1   g068(.A1(KEYINPUT0), .A2(G128), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n244), .A2(new_n246), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(G143), .B(G146), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT0), .B(G128), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  OAI22_X1  g074(.A1(new_n253), .A2(KEYINPUT82), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n253), .A2(KEYINPUT82), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT84), .ZN(new_n264));
  INV_X1    g078(.A(G224), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n264), .B1(new_n265), .B2(G953), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT84), .A3(G224), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XOR2_X1   g083(.A(new_n269), .B(KEYINPUT83), .Z(new_n270));
  XNOR2_X1  g084(.A(new_n263), .B(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n242), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n268), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n273), .B1(new_n261), .B2(new_n262), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n198), .B1(new_n222), .B2(new_n225), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n217), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n188), .B(KEYINPUT8), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n226), .A2(new_n198), .A3(new_n229), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n276), .B(new_n277), .C1(new_n278), .C2(new_n217), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  NOR3_X1   g094(.A1(new_n261), .A2(new_n262), .A3(new_n273), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n237), .A2(new_n239), .ZN(new_n283));
  AOI21_X1  g097(.A(G902), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(G210), .B1(G237), .B2(G902), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(KEYINPUT85), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n272), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n287), .B1(new_n272), .B2(new_n284), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n187), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G469), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  XNOR2_X1  g106(.A(G110), .B(G140), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n267), .A2(G227), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n293), .B(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n255), .ZN(new_n297));
  OR2_X1    g111(.A1(KEYINPUT0), .A2(G128), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n247), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n212), .A2(new_n256), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT79), .B1(new_n235), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT79), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n210), .A2(new_n302), .A3(new_n260), .A4(new_n212), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT68), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n248), .A2(G128), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(new_n257), .ZN(new_n307));
  INV_X1    g121(.A(new_n251), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n249), .A2(KEYINPUT68), .A3(new_n251), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n209), .A2(new_n216), .A3(KEYINPUT10), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT10), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n249), .A2(new_n251), .A3(new_n209), .A4(new_n216), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n311), .A2(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n304), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G134), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT11), .B1(new_n317), .B2(G137), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT11), .ZN(new_n319));
  INV_X1    g133(.A(G137), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(G134), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT65), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n320), .B2(G134), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n317), .A2(KEYINPUT65), .A3(G137), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G131), .ZN(new_n327));
  INV_X1    g141(.A(G131), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n322), .A2(new_n328), .A3(new_n324), .A4(new_n325), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n316), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n329), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n324), .A2(new_n325), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n328), .B1(new_n333), .B2(new_n322), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n304), .A2(new_n335), .A3(new_n315), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n296), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n314), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n249), .A2(new_n251), .B1(new_n209), .B2(new_n216), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n330), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT12), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n330), .B(KEYINPUT12), .C1(new_n338), .C2(new_n339), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n336), .A2(new_n296), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n291), .B(new_n292), .C1(new_n337), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(G469), .A2(G902), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n336), .A2(new_n344), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n295), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n331), .A2(new_n336), .A3(new_n296), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(G469), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n347), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT9), .B(G234), .ZN(new_n354));
  OAI21_X1  g168(.A(G221), .B1(new_n354), .B2(G902), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT77), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(KEYINPUT78), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n254), .A2(KEYINPUT16), .A3(G140), .ZN(new_n360));
  XNOR2_X1  g174(.A(G125), .B(G140), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n360), .B1(new_n361), .B2(KEYINPUT16), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(G146), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT16), .ZN(new_n364));
  INV_X1    g178(.A(G140), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(G125), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(G125), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n254), .A2(G140), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(G146), .B(new_n366), .C1(new_n369), .C2(new_n364), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n363), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G237), .ZN(new_n373));
  AND4_X1   g187(.A1(G143), .A2(new_n373), .A3(new_n267), .A4(G214), .ZN(new_n374));
  NOR2_X1   g188(.A1(G237), .A2(G953), .ZN(new_n375));
  AOI21_X1  g189(.A(G143), .B1(new_n375), .B2(G214), .ZN(new_n376));
  OAI21_X1  g190(.A(G131), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT17), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n373), .A2(new_n267), .A3(G214), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n245), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n375), .A2(G143), .A3(G214), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n328), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n377), .A2(new_n378), .A3(new_n382), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n377), .A2(KEYINPUT89), .A3(new_n378), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT89), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n328), .B1(new_n380), .B2(new_n381), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n385), .B1(new_n386), .B2(KEYINPUT17), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n372), .B(new_n383), .C1(new_n384), .C2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G113), .B(G122), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(new_n200), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n369), .A2(G146), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n367), .A2(new_n368), .A3(new_n243), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(KEYINPUT18), .A2(G131), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n395), .B1(new_n374), .B2(new_n376), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n380), .A2(new_n381), .A3(new_n394), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n393), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT86), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT86), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n393), .A2(new_n396), .A3(new_n400), .A4(new_n397), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n388), .A2(new_n390), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n390), .B1(new_n388), .B2(new_n402), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n292), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n406), .A2(G475), .ZN(new_n407));
  NOR2_X1   g221(.A1(G475), .A2(G902), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n377), .A2(new_n382), .B1(new_n362), .B2(G146), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT19), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n369), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT19), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT87), .B1(new_n413), .B2(new_n243), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT87), .ZN(new_n415));
  AOI211_X1 g229(.A(new_n415), .B(G146), .C1(new_n411), .C2(new_n412), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n409), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n402), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT88), .ZN(new_n419));
  INV_X1    g233(.A(new_n390), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n403), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n419), .B1(new_n418), .B2(new_n420), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n408), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT20), .ZN(new_n425));
  INV_X1    g239(.A(new_n412), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT19), .B1(new_n367), .B2(new_n368), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n243), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n415), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n413), .A2(KEYINPUT87), .A3(new_n243), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n431), .A2(new_n409), .B1(new_n399), .B2(new_n401), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT88), .B1(new_n432), .B2(new_n390), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n403), .A3(new_n421), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(new_n408), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n407), .B1(new_n425), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G217), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n354), .A2(new_n438), .A3(G953), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n220), .A2(G122), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(KEYINPUT14), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n220), .A2(G122), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n441), .B1(new_n443), .B2(KEYINPUT14), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n442), .B1(new_n444), .B2(KEYINPUT90), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT90), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n446), .B(new_n441), .C1(new_n443), .C2(KEYINPUT14), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n203), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n443), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(new_n441), .A3(new_n203), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n245), .A2(G128), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n250), .A2(G143), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n317), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n317), .B1(new_n451), .B2(new_n452), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n450), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n448), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n203), .B1(new_n449), .B2(new_n441), .ZN(new_n458));
  INV_X1    g272(.A(new_n441), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n459), .A2(G107), .A3(new_n443), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n453), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT13), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n451), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n245), .A2(KEYINPUT13), .A3(G128), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n464), .A3(new_n452), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n465), .A2(G134), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n440), .B1(new_n457), .B2(new_n467), .ZN(new_n468));
  OAI221_X1 g282(.A(new_n439), .B1(new_n461), .B2(new_n466), .C1(new_n448), .C2(new_n456), .ZN(new_n469));
  AOI21_X1  g283(.A(G902), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G478), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(KEYINPUT15), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  AOI211_X1 g288(.A(G902), .B(new_n472), .C1(new_n468), .C2(new_n469), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n267), .A2(G952), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(G234), .B2(G237), .ZN(new_n478));
  AOI211_X1 g292(.A(new_n292), .B(new_n267), .C1(G234), .C2(G237), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT21), .B(G898), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n437), .A2(new_n482), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n290), .A2(new_n359), .A3(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(G472), .A2(G902), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n259), .A2(KEYINPUT64), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT64), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n299), .A2(new_n487), .A3(new_n256), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT66), .B1(new_n335), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT66), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n330), .A2(new_n491), .A3(new_n486), .A4(new_n488), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n317), .A2(G137), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n320), .A2(G134), .ZN(new_n494));
  OAI21_X1  g308(.A(G131), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n329), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n249), .A2(new_n251), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n490), .A2(new_n492), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n496), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n311), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n330), .A2(new_n260), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(KEYINPUT30), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT69), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n311), .A2(new_n503), .B1(new_n330), .B2(new_n260), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT69), .A3(KEYINPUT30), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n502), .A2(new_n508), .A3(new_n199), .A4(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n233), .A2(new_n196), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT70), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT70), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n199), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n509), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n375), .A2(G210), .ZN(new_n518));
  XOR2_X1   g332(.A(new_n518), .B(KEYINPUT27), .Z(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT26), .B(G101), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n511), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT31), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT31), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n511), .A2(new_n525), .A3(new_n522), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n521), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n509), .A2(new_n516), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT28), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  XOR2_X1   g346(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n486), .B(new_n488), .C1(new_n332), .C2(new_n334), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n498), .B1(new_n535), .B2(KEYINPUT66), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n512), .B1(new_n536), .B2(new_n492), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n534), .B1(new_n537), .B2(new_n517), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT72), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n532), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(KEYINPUT72), .B(new_n534), .C1(new_n537), .C2(new_n517), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n528), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n485), .B1(new_n527), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT32), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n485), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(new_n544), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n547), .B1(new_n527), .B2(new_n542), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n500), .A2(new_n199), .B1(new_n509), .B2(new_n516), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n539), .B1(new_n549), .B2(new_n533), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n550), .A2(new_n528), .A3(new_n541), .A4(new_n531), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n511), .A2(new_n529), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n521), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT29), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n509), .A2(new_n516), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT28), .B1(new_n517), .B2(new_n556), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n557), .A2(new_n531), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n521), .A2(new_n554), .ZN(new_n559));
  AOI21_X1  g373(.A(G902), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G472), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n545), .A2(new_n548), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n438), .B1(G234), .B2(new_n292), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(KEYINPUT73), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT23), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n218), .B2(G128), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n218), .A2(G128), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n250), .A2(KEYINPUT23), .A3(G119), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G110), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT24), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT24), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(G110), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT74), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n250), .B2(G119), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n218), .A2(KEYINPUT74), .A3(G128), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n250), .A2(G119), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n570), .A2(new_n571), .B1(new_n576), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n370), .A2(new_n392), .ZN(new_n583));
  OR2_X1    g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n575), .A2(new_n578), .A3(new_n579), .A4(new_n580), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(G110), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n585), .B(new_n587), .C1(new_n363), .C2(new_n371), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT75), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n584), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n587), .A2(new_n585), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n366), .B1(new_n369), .B2(new_n364), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n243), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n591), .B1(new_n370), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n582), .A2(new_n583), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT75), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT22), .B(G137), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n590), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n584), .A2(new_n588), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n602), .A2(KEYINPUT75), .A3(new_n599), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT25), .B1(new_n604), .B2(new_n292), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT25), .ZN(new_n606));
  AOI211_X1 g420(.A(new_n606), .B(G902), .C1(new_n601), .C2(new_n603), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n565), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n604), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n564), .A2(G902), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n608), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n563), .A2(KEYINPUT76), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT76), .B1(new_n563), .B2(new_n613), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n484), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(G101), .ZN(G3));
  AND3_X1   g431(.A1(new_n511), .A2(new_n525), .A3(new_n522), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n525), .B1(new_n511), .B2(new_n522), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n550), .A2(new_n541), .A3(new_n531), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n521), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n546), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(G472), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n620), .A2(new_n622), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n624), .B1(new_n625), .B2(new_n292), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT91), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(G902), .B1(new_n620), .B2(new_n622), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT91), .B1(new_n629), .B2(new_n624), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n285), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n272), .B2(new_n284), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n481), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n272), .A2(new_n284), .A3(new_n633), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n635), .A2(new_n187), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n471), .A2(G902), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT33), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n468), .A2(new_n469), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n640), .B1(new_n468), .B2(new_n469), .ZN(new_n643));
  OAI211_X1 g457(.A(KEYINPUT92), .B(new_n639), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n639), .ZN(new_n645));
  INV_X1    g459(.A(new_n643), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n645), .B1(new_n646), .B2(new_n641), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT92), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(new_n470), .B2(G478), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n644), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n425), .A2(new_n436), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n406), .A2(G475), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n638), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n359), .A2(new_n612), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n632), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT34), .B(G104), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G6));
  NAND3_X1  g473(.A1(new_n425), .A2(KEYINPUT93), .A3(new_n436), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n436), .A2(KEYINPUT93), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n660), .A2(new_n652), .A3(new_n476), .A4(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n638), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n632), .A2(new_n656), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT94), .Z(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT35), .B(G107), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  NOR2_X1   g481(.A1(new_n600), .A2(KEYINPUT36), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n602), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n610), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n608), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n437), .A2(new_n671), .A3(new_n482), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n290), .A2(new_n672), .A3(new_n359), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n292), .B1(new_n527), .B2(new_n542), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n627), .A3(G472), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n673), .A2(new_n543), .A3(new_n675), .A4(new_n630), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT37), .B(G110), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G12));
  NAND3_X1  g492(.A1(new_n635), .A2(new_n187), .A3(new_n637), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n353), .A2(new_n671), .A3(new_n358), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n563), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(G900), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n479), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n478), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n662), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n250), .ZN(G30));
  AND3_X1   g504(.A1(new_n434), .A2(new_n435), .A3(new_n408), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n435), .B1(new_n434), .B2(new_n408), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n652), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n476), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n552), .A2(new_n528), .ZN(new_n696));
  OR3_X1    g510(.A1(new_n517), .A2(new_n556), .A3(new_n528), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n292), .A3(new_n697), .ZN(new_n698));
  AOI22_X1  g512(.A1(new_n625), .A2(new_n547), .B1(G472), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n545), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n272), .A2(new_n284), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n286), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n272), .A2(new_n284), .A3(new_n287), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n187), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n671), .A2(new_n707), .ZN(new_n708));
  AND4_X1   g522(.A1(new_n695), .A2(new_n700), .A3(new_n706), .A4(new_n708), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n709), .A2(KEYINPUT96), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(KEYINPUT96), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n686), .B(KEYINPUT39), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n359), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT40), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n710), .A2(new_n711), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G143), .ZN(G45));
  INV_X1    g531(.A(new_n650), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n693), .A2(new_n718), .A3(new_n686), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n682), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n243), .ZN(G48));
  OAI21_X1  g536(.A(new_n292), .B1(new_n337), .B2(new_n346), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(G469), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT97), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n725), .A3(new_n347), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n723), .A2(KEYINPUT97), .A3(G469), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n356), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n563), .A2(new_n613), .A3(new_n655), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT41), .B(G113), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  NAND4_X1  g545(.A1(new_n563), .A2(new_n613), .A3(new_n663), .A4(new_n728), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G116), .ZN(G18));
  NAND2_X1  g547(.A1(new_n726), .A2(new_n727), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n272), .A2(new_n284), .A3(new_n633), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n735), .A2(new_n634), .A3(new_n707), .ZN(new_n736));
  INV_X1    g550(.A(new_n356), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n672), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n563), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  AOI21_X1  g555(.A(new_n528), .B1(new_n557), .B2(new_n531), .ZN(new_n742));
  OR3_X1    g556(.A1(new_n619), .A2(new_n742), .A3(KEYINPUT98), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT98), .B1(new_n619), .B2(new_n742), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n526), .A3(new_n744), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n745), .A2(new_n485), .B1(new_n674), .B2(G472), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n638), .A2(new_n694), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n746), .A2(new_n747), .A3(new_n613), .A4(new_n728), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  NAND4_X1  g563(.A1(new_n738), .A2(new_n671), .A3(new_n746), .A4(new_n720), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  INV_X1    g565(.A(KEYINPUT42), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n352), .A2(new_n348), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n304), .A2(new_n335), .A3(new_n315), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n335), .B1(new_n304), .B2(new_n315), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n295), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI211_X1 g570(.A(G469), .B(G902), .C1(new_n756), .C2(new_n345), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT99), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT99), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n347), .A2(new_n759), .A3(new_n348), .A4(new_n352), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n758), .A2(new_n737), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n702), .A2(new_n187), .A3(new_n703), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n563), .A2(new_n763), .A3(new_n613), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n752), .B1(new_n764), .B2(new_n719), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT100), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n766), .B1(new_n625), .B2(new_n547), .ZN(new_n767));
  INV_X1    g581(.A(new_n547), .ZN(new_n768));
  AOI211_X1 g582(.A(KEYINPUT100), .B(new_n768), .C1(new_n620), .C2(new_n622), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n544), .A2(new_n543), .B1(new_n561), .B2(G472), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n612), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n288), .A2(new_n289), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n773), .A2(new_n653), .A3(new_n187), .A4(new_n686), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n758), .A2(KEYINPUT42), .A3(new_n737), .A4(new_n760), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT101), .B1(new_n772), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n548), .A2(KEYINPUT100), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n625), .A2(new_n766), .A3(new_n547), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n545), .A2(new_n778), .A3(new_n562), .A4(new_n779), .ZN(new_n780));
  AND4_X1   g594(.A1(KEYINPUT101), .A2(new_n776), .A3(new_n780), .A4(new_n613), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n765), .B1(new_n777), .B2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT102), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g598(.A(KEYINPUT102), .B(new_n765), .C1(new_n777), .C2(new_n781), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XOR2_X1   g600(.A(KEYINPUT103), .B(G131), .Z(new_n787));
  XNOR2_X1  g601(.A(new_n786), .B(new_n787), .ZN(G33));
  NAND4_X1  g602(.A1(new_n563), .A2(new_n763), .A3(new_n613), .A4(new_n688), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G134), .ZN(G36));
  NAND2_X1  g604(.A1(new_n631), .A2(new_n671), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT105), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT105), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n631), .A2(new_n793), .A3(new_n671), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n437), .A2(new_n718), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n796), .B(KEYINPUT43), .Z(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT44), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n795), .A2(KEYINPUT44), .A3(new_n797), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n350), .A2(new_n351), .ZN(new_n802));
  OAI21_X1  g616(.A(G469), .B1(new_n802), .B2(KEYINPUT45), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n803), .A2(KEYINPUT104), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(KEYINPUT45), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(KEYINPUT104), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT46), .B1(new_n807), .B2(new_n348), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n757), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(KEYINPUT46), .A3(new_n348), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n737), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n812), .A2(new_n713), .A3(new_n762), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n800), .A2(new_n801), .A3(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G137), .ZN(G39));
  INV_X1    g629(.A(KEYINPUT47), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n811), .A2(KEYINPUT47), .A3(new_n737), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n563), .A2(new_n613), .A3(new_n774), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G140), .ZN(G42));
  OAI211_X1 g636(.A(new_n187), .B(new_n636), .C1(new_n288), .C2(new_n289), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n652), .B(new_n476), .C1(new_n691), .C2(new_n692), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n823), .B1(new_n654), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n628), .A2(new_n825), .A3(new_n630), .A4(new_n656), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n826), .A2(new_n729), .A3(new_n732), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n474), .A2(new_n475), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n828), .A2(new_n652), .A3(new_n686), .ZN(new_n829));
  AND4_X1   g643(.A1(KEYINPUT107), .A2(new_n660), .A3(new_n661), .A4(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n830), .A2(new_n680), .A3(new_n762), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n660), .A2(new_n829), .A3(new_n661), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT107), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n831), .A2(new_n563), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n761), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n762), .A2(new_n719), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n746), .A2(new_n671), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n789), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n740), .A2(new_n676), .A3(new_n748), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n616), .A2(new_n827), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n563), .B(new_n681), .C1(new_n688), .C2(new_n720), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n679), .A2(new_n671), .A3(new_n687), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n700), .A2(new_n843), .A3(new_n695), .A4(new_n836), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n750), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n842), .A2(new_n750), .A3(new_n844), .A4(KEYINPUT52), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n841), .A2(new_n784), .A3(new_n785), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n850), .A2(KEYINPUT108), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT108), .B1(new_n850), .B2(new_n851), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n850), .A2(new_n851), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT109), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n841), .A2(KEYINPUT53), .A3(new_n782), .A4(new_n849), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n850), .A2(new_n851), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n859), .A2(KEYINPUT110), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(KEYINPUT110), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n856), .B(new_n858), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT108), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n854), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n850), .A2(KEYINPUT108), .A3(new_n851), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT109), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n868), .A3(KEYINPUT54), .ZN(new_n869));
  INV_X1    g683(.A(new_n700), .ZN(new_n870));
  INV_X1    g684(.A(new_n762), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n728), .A2(new_n871), .ZN(new_n872));
  AND4_X1   g686(.A1(new_n613), .A2(new_n870), .A3(new_n478), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n437), .A2(new_n650), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n797), .A2(new_n478), .A3(new_n872), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n746), .A2(new_n671), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n873), .A2(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n797), .A2(new_n478), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n773), .B(new_n705), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n707), .A3(new_n728), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n746), .A2(new_n613), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n883), .A2(KEYINPUT50), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(KEYINPUT50), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n878), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n734), .A2(new_n357), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n817), .A2(new_n818), .A3(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n879), .A2(new_n882), .A3(new_n762), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT111), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n888), .A2(KEYINPUT111), .A3(new_n889), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT51), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT112), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n886), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(KEYINPUT112), .B(new_n878), .C1(new_n884), .C2(new_n885), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n896), .A2(new_n890), .A3(KEYINPUT51), .A4(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n876), .A2(new_n772), .ZN(new_n899));
  AND2_X1   g713(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n900));
  NOR2_X1   g714(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n899), .A2(new_n900), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n477), .B(KEYINPUT113), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n873), .B2(new_n653), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n879), .A2(new_n882), .ZN(new_n907));
  AOI211_X1 g721(.A(new_n902), .B(new_n906), .C1(new_n738), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n898), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n894), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n857), .A2(new_n862), .A3(new_n869), .A4(new_n910), .ZN(new_n911));
  OR2_X1    g725(.A1(G952), .A2(G953), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n734), .B(KEYINPUT49), .ZN(new_n914));
  NOR4_X1   g728(.A1(new_n796), .A2(new_n612), .A3(new_n707), .A4(new_n357), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n914), .A2(new_n870), .A3(new_n880), .A4(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT106), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT115), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT115), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n913), .A2(new_n920), .A3(new_n917), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(G75));
  NOR2_X1   g736(.A1(new_n267), .A2(G952), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT116), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(G210), .A3(G902), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT56), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n242), .B(new_n271), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT55), .Z(new_n931));
  OR2_X1    g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n929), .A2(new_n931), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n925), .B1(new_n932), .B2(new_n933), .ZN(G51));
  INV_X1    g748(.A(new_n807), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n926), .A2(G902), .A3(new_n935), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT117), .Z(new_n937));
  XNOR2_X1  g751(.A(new_n926), .B(new_n856), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n348), .B(KEYINPUT57), .ZN(new_n939));
  OAI22_X1  g753(.A1(new_n938), .A2(new_n939), .B1(new_n337), .B2(new_n346), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n923), .B1(new_n937), .B2(new_n940), .ZN(G54));
  NAND4_X1  g755(.A1(new_n926), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n942));
  INV_X1    g756(.A(new_n434), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(new_n945), .A3(new_n923), .ZN(G60));
  NAND2_X1  g760(.A1(G478), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT59), .Z(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n642), .B2(new_n643), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n924), .B1(new_n938), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n642), .A2(new_n643), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n857), .A2(new_n862), .A3(new_n869), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n949), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n951), .B1(new_n952), .B2(new_n954), .ZN(G63));
  XNOR2_X1  g769(.A(KEYINPUT118), .B(KEYINPUT60), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n438), .A2(new_n292), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n926), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n609), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n669), .B(KEYINPUT119), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n926), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n960), .A2(new_n924), .A3(new_n962), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g778(.A(G953), .B1(new_n480), .B2(new_n265), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n827), .A2(new_n616), .A3(new_n840), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n966), .B2(G953), .ZN(new_n967));
  INV_X1    g781(.A(new_n242), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(G898), .B2(new_n267), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT120), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n967), .B(new_n970), .ZN(G69));
  NAND3_X1  g785(.A1(new_n502), .A2(new_n508), .A3(new_n510), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(new_n413), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n842), .A2(new_n750), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n716), .A2(new_n974), .A3(KEYINPUT62), .ZN(new_n975));
  AOI21_X1  g789(.A(KEYINPUT62), .B1(new_n716), .B2(new_n974), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n821), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n714), .A2(new_n871), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n654), .B2(new_n824), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(new_n614), .B2(new_n615), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n814), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT121), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n814), .A2(KEYINPUT121), .A3(new_n980), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n977), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n973), .B1(new_n985), .B2(G953), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(KEYINPUT122), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT122), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n988), .B(new_n973), .C1(new_n985), .C2(G953), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT123), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n772), .A2(new_n736), .A3(new_n695), .ZN(new_n992));
  OR3_X1    g806(.A1(new_n812), .A2(new_n713), .A3(new_n992), .ZN(new_n993));
  AND4_X1   g807(.A1(new_n786), .A2(new_n821), .A3(new_n789), .A4(new_n993), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n814), .A2(KEYINPUT124), .A3(new_n974), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT124), .B1(new_n814), .B2(new_n974), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(KEYINPUT125), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT125), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n994), .B(new_n999), .C1(new_n995), .C2(new_n996), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n998), .A2(new_n267), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n973), .B1(G900), .B2(G953), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n990), .A2(new_n991), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n267), .B1(G227), .B2(G900), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1005), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n990), .A2(new_n991), .A3(new_n1007), .A4(new_n1003), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1006), .A2(new_n1008), .ZN(G72));
  XNOR2_X1  g823(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n624), .A2(new_n292), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1010), .B(new_n1011), .Z(new_n1012));
  INV_X1    g826(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1013), .B1(new_n553), .B2(new_n523), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n923), .B1(new_n867), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n985), .A2(new_n966), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n696), .B1(new_n1016), .B2(new_n1012), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI211_X1 g833(.A(KEYINPUT127), .B(new_n696), .C1(new_n1016), .C2(new_n1012), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1015), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n998), .A2(new_n966), .A3(new_n1000), .ZN(new_n1022));
  AOI211_X1 g836(.A(new_n528), .B(new_n552), .C1(new_n1022), .C2(new_n1012), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1021), .A2(new_n1023), .ZN(G57));
endmodule


