//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1255,
    new_n1256, new_n1257, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n212), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n210), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n201), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n215), .B1(KEYINPUT1), .B2(new_n225), .C1(new_n228), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n225), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT64), .Z(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G68), .Z(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G1), .A3(G13), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  AOI21_X1  g0055(.A(G1698), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n256), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(new_n255), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G257), .A3(G1698), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n251), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT5), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n209), .B(G45), .C1(new_n261), .C2(KEYINPUT5), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n262), .B1(new_n263), .B2(KEYINPUT83), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT83), .ZN(new_n265));
  INV_X1    g0065(.A(G45), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G1), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT5), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G41), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n265), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  OAI211_X1 g0070(.A(G264), .B(new_n251), .C1(new_n264), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT89), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n263), .A2(KEYINPUT83), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n267), .A2(new_n265), .A3(new_n269), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(new_n274), .A3(new_n262), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT89), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n275), .A2(new_n276), .A3(G264), .A4(new_n251), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n260), .B1(new_n272), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n281), .A2(new_n274), .A3(new_n273), .A4(new_n262), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n278), .A2(G190), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n226), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT23), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(new_n210), .B2(G107), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G116), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n289), .B1(G20), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n258), .A2(new_n210), .A3(G87), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT22), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT22), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n258), .A2(new_n294), .A3(new_n210), .A4(G87), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n291), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  XOR2_X1   g0096(.A(KEYINPUT88), .B(KEYINPUT24), .Z(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  AOI211_X1 g0099(.A(new_n297), .B(new_n291), .C1(new_n293), .C2(new_n295), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n285), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(new_n226), .A3(new_n284), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n209), .B2(G33), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT25), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(new_n302), .B2(G107), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n302), .A2(new_n305), .A3(G107), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n304), .A2(G107), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n283), .A2(new_n301), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G200), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n278), .B2(new_n282), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n272), .A2(new_n277), .ZN(new_n314));
  INV_X1    g0114(.A(new_n260), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(new_n315), .A3(new_n282), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G169), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT90), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT90), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(new_n319), .A3(G169), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n278), .A2(G179), .A3(new_n282), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n301), .A2(new_n309), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n313), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n210), .A2(G33), .ZN(new_n325));
  INV_X1    g0125(.A(G77), .ZN(new_n326));
  OAI22_X1  g0126(.A1(new_n325), .A2(new_n326), .B1(new_n210), .B2(G68), .ZN(new_n327));
  NOR2_X1   g0127(.A1(G20), .A2(G33), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n327), .A2(KEYINPUT74), .B1(new_n202), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n327), .A2(KEYINPUT74), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n285), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  XOR2_X1   g0132(.A(new_n332), .B(KEYINPUT11), .Z(new_n333));
  INV_X1    g0133(.A(new_n302), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n217), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT12), .B1(new_n335), .B2(KEYINPUT75), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(KEYINPUT75), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n303), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT71), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT71), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n303), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n209), .A2(G20), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n340), .A2(G68), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n333), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n258), .A2(G232), .A3(G1698), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G97), .ZN(new_n349));
  INV_X1    g0149(.A(G1698), .ZN(new_n350));
  AND2_X1   g0150(.A1(KEYINPUT3), .A2(G33), .ZN(new_n351));
  NOR2_X1   g0151(.A1(KEYINPUT3), .A2(G33), .ZN(new_n352));
  OAI211_X1 g0152(.A(G226), .B(new_n350), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n348), .A2(new_n349), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n279), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(new_n280), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT66), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n209), .B(KEYINPUT66), .C1(G41), .C2(G45), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(new_n251), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT67), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n361), .A2(KEYINPUT67), .A3(new_n251), .A4(new_n362), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n218), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT13), .B1(new_n359), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n366), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G238), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT13), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(new_n358), .A4(new_n355), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n368), .A2(new_n372), .A3(G179), .ZN(new_n373));
  INV_X1    g0173(.A(G169), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n368), .B2(new_n372), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT14), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI211_X1 g0177(.A(KEYINPUT14), .B(new_n374), .C1(new_n368), .C2(new_n372), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n347), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n368), .A2(new_n372), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G190), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n381), .B(new_n346), .C1(new_n311), .C2(new_n380), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G20), .A2(G77), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT15), .B(G87), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT8), .B(G58), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n383), .B1(new_n384), .B2(new_n325), .C1(new_n329), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n285), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n340), .A2(G77), .A3(new_n342), .A4(new_n343), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n334), .A2(new_n326), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G244), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(new_n365), .B2(new_n366), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n258), .A2(G232), .A3(new_n350), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n351), .A2(new_n352), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G107), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n258), .A2(G1698), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n394), .B(new_n396), .C1(new_n397), .C2(new_n218), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n357), .B1(new_n398), .B2(new_n279), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n390), .B1(new_n400), .B2(new_n374), .ZN(new_n401));
  INV_X1    g0201(.A(G179), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n393), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n398), .A2(new_n279), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n358), .ZN(new_n406));
  OAI21_X1  g0206(.A(G200), .B1(new_n406), .B2(new_n392), .ZN(new_n407));
  INV_X1    g0207(.A(G190), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n407), .B(new_n390), .C1(new_n408), .C2(new_n400), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n379), .A2(new_n382), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT68), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n256), .A2(new_n412), .A3(G222), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n412), .B1(new_n256), .B2(G222), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(G223), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n397), .A2(new_n416), .B1(new_n326), .B2(new_n258), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n279), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n369), .A2(G226), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n418), .A2(new_n419), .A3(G190), .A4(new_n358), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n343), .A2(G50), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n303), .A2(new_n421), .B1(G50), .B2(new_n302), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT69), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI221_X1 g0224(.A(KEYINPUT69), .B1(G50), .B2(new_n302), .C1(new_n303), .C2(new_n421), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n328), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n325), .B2(new_n385), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n424), .A2(new_n425), .B1(new_n427), .B2(new_n285), .ZN(new_n428));
  NAND2_X1  g0228(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n428), .B2(new_n430), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n420), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n418), .A2(new_n419), .A3(new_n358), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G200), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT73), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n435), .B(new_n437), .C1(new_n438), .C2(KEYINPUT10), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n428), .B1(new_n436), .B2(new_n374), .ZN(new_n440));
  INV_X1    g0240(.A(new_n436), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT70), .B1(new_n441), .B2(new_n402), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT70), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n436), .A2(new_n443), .A3(G179), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n440), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT10), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n420), .A2(new_n431), .A3(new_n438), .A4(new_n433), .ZN(new_n447));
  INV_X1    g0247(.A(new_n437), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n446), .B(new_n447), .C1(new_n448), .C2(new_n434), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n439), .A2(new_n445), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n411), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT78), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n361), .A2(G232), .A3(new_n251), .A4(new_n362), .ZN(new_n453));
  NOR2_X1   g0253(.A1(G223), .A2(G1698), .ZN(new_n454));
  INV_X1    g0254(.A(G226), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(G1698), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n456), .A2(new_n258), .B1(G33), .B2(G87), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n358), .B(new_n453), .C1(new_n457), .C2(new_n251), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(G190), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n455), .A2(G1698), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(G223), .B2(G1698), .ZN(new_n461));
  OAI22_X1  g0261(.A1(new_n461), .A2(new_n395), .B1(new_n253), .B2(new_n219), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n357), .B1(new_n462), .B2(new_n279), .ZN(new_n463));
  AOI21_X1  g0263(.A(G200), .B1(new_n463), .B2(new_n453), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n452), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n458), .A2(new_n311), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n466), .B(KEYINPUT78), .C1(G190), .C2(new_n458), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n385), .B1(new_n209), .B2(G20), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n469), .A2(new_n339), .B1(new_n334), .B2(new_n385), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n254), .A2(new_n210), .A3(new_n255), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT7), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT7), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n254), .A2(new_n473), .A3(new_n210), .A4(new_n255), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(G68), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT76), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n472), .A2(KEYINPUT76), .A3(G68), .A4(new_n474), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g0279(.A(G58), .B(G68), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n480), .A2(G20), .B1(G159), .B2(new_n328), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(KEYINPUT16), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n475), .A2(new_n481), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT16), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT77), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n483), .A2(KEYINPUT77), .A3(new_n484), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n482), .A2(new_n487), .A3(new_n285), .A4(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n468), .A2(new_n470), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT17), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n470), .ZN(new_n493));
  INV_X1    g0293(.A(new_n481), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n477), .B2(new_n478), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n495), .A2(KEYINPUT16), .B1(new_n226), .B2(new_n284), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT77), .B1(new_n483), .B2(new_n484), .ZN(new_n497));
  AOI211_X1 g0297(.A(new_n486), .B(KEYINPUT16), .C1(new_n475), .C2(new_n481), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n493), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n458), .A2(new_n402), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n501), .B1(G169), .B2(new_n458), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT18), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n489), .A2(new_n470), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT18), .ZN(new_n505));
  INV_X1    g0305(.A(new_n502), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n500), .A2(KEYINPUT17), .A3(new_n468), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n492), .A2(new_n503), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT79), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n492), .A2(new_n508), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n503), .A2(new_n507), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT79), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n451), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n264), .A2(new_n270), .ZN(new_n516));
  OAI211_X1 g0316(.A(G264), .B(G1698), .C1(new_n351), .C2(new_n352), .ZN(new_n517));
  OAI211_X1 g0317(.A(G257), .B(new_n350), .C1(new_n351), .C2(new_n352), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n254), .A2(G303), .A3(new_n255), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n516), .A2(new_n281), .B1(new_n520), .B2(new_n279), .ZN(new_n521));
  OAI211_X1 g0321(.A(G270), .B(new_n251), .C1(new_n264), .C2(new_n270), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT86), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT86), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n275), .A2(new_n524), .A3(G270), .A4(new_n251), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n521), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(G13), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n527), .A2(G1), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(G116), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G20), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G283), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n533), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(new_n285), .A3(new_n531), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT20), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n534), .A2(KEYINPUT20), .A3(new_n285), .A4(new_n531), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n532), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n530), .B1(new_n209), .B2(G33), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n340), .A2(new_n342), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n374), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT87), .B1(new_n526), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT21), .ZN(new_n544));
  OR2_X1    g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n521), .A2(new_n523), .A3(G179), .A4(new_n525), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n539), .A2(new_n541), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n543), .A2(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n548), .B1(new_n526), .B2(G200), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(new_n408), .B2(new_n526), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n545), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n258), .A2(G244), .A3(new_n350), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT4), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n554), .A2(KEYINPUT82), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n533), .B1(new_n554), .B2(KEYINPUT82), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n350), .A2(KEYINPUT4), .A3(G244), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n220), .B2(new_n350), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n557), .B1(new_n559), .B2(new_n258), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n279), .ZN(new_n562));
  OAI211_X1 g0362(.A(G257), .B(new_n251), .C1(new_n264), .C2(new_n270), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n562), .A2(new_n402), .A3(new_n282), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n282), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n251), .B1(new_n556), .B2(new_n560), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n374), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G97), .A2(G107), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n207), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT6), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT80), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n205), .A2(KEYINPUT6), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n207), .A2(new_n573), .A3(new_n576), .A4(new_n570), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n210), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n329), .A2(new_n326), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT81), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n472), .A2(G107), .A3(new_n474), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n578), .A2(KEYINPUT81), .A3(new_n579), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n285), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n302), .A2(G97), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n585), .B1(new_n304), .B2(G97), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n569), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n586), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n575), .A2(new_n577), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n579), .B1(new_n590), .B2(G20), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT81), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n580), .A3(new_n581), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n589), .B1(new_n594), .B2(new_n285), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n311), .B1(new_n565), .B2(new_n566), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n562), .A2(new_n282), .A3(new_n563), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n596), .B1(new_n597), .B2(G190), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT85), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n220), .B1(new_n209), .B2(G45), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n251), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n267), .A2(G274), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT84), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT84), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n602), .A2(new_n606), .A3(new_n603), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n258), .A2(G238), .A3(new_n350), .ZN(new_n609));
  OAI211_X1 g0409(.A(G244), .B(G1698), .C1(new_n351), .C2(new_n352), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n290), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n279), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n608), .A2(new_n612), .A3(G179), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n374), .B1(new_n608), .B2(new_n612), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n600), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n608), .A2(new_n612), .A3(G179), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n605), .A2(new_n607), .B1(new_n611), .B2(new_n279), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n616), .B(KEYINPUT85), .C1(new_n374), .C2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n258), .A2(new_n210), .A3(G68), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT19), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n210), .B1(new_n349), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(G87), .B2(new_n207), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n620), .B1(new_n325), .B2(new_n205), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n619), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n285), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n384), .A2(new_n334), .ZN(new_n626));
  INV_X1    g0426(.A(new_n304), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n384), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n615), .A2(new_n618), .A3(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n625), .B(new_n626), .C1(new_n219), .C2(new_n627), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n608), .A2(new_n612), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n630), .B1(G200), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n617), .A2(G190), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n588), .A2(new_n599), .A3(new_n629), .A4(new_n634), .ZN(new_n635));
  AND4_X1   g0435(.A1(new_n324), .A2(new_n515), .A3(new_n552), .A4(new_n635), .ZN(G372));
  INV_X1    g0436(.A(new_n312), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n637), .A2(new_n301), .A3(new_n309), .A4(new_n283), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n616), .B1(new_n617), .B2(new_n374), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n632), .A2(new_n633), .B1(new_n639), .B2(new_n628), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n638), .A2(new_n588), .A3(new_n599), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n526), .A2(new_n542), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT87), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(new_n643), .A3(new_n544), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n547), .A2(new_n548), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n543), .A2(new_n544), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT91), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT91), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n545), .A2(new_n549), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n320), .A2(new_n321), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n319), .B1(new_n316), .B2(G169), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n323), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n641), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n595), .A2(new_n568), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(new_n634), .A3(new_n629), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(KEYINPUT26), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n639), .A2(new_n628), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT92), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n569), .A2(new_n587), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT92), .B1(new_n595), .B2(new_n568), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n661), .A2(new_n662), .A3(new_n640), .A4(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n658), .A2(new_n659), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n515), .B1(new_n655), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n445), .ZN(new_n667));
  INV_X1    g0467(.A(new_n379), .ZN(new_n668));
  INV_X1    g0468(.A(new_n404), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n512), .A2(new_n382), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n513), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n439), .A2(new_n449), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n667), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n666), .A2(new_n674), .ZN(G369));
  OR3_X1    g0475(.A1(new_n529), .A2(KEYINPUT27), .A3(G20), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT27), .B1(new_n529), .B2(G20), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n654), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n680), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n654), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT93), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n323), .A2(new_n680), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n685), .B1(new_n324), .B2(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n654), .A2(new_n685), .A3(new_n638), .A4(new_n686), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n684), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT94), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n654), .A2(new_n638), .A3(new_n686), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT93), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n688), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(KEYINPUT94), .A3(new_n684), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n682), .B1(new_n646), .B2(new_n647), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT95), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n681), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G330), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n548), .A2(new_n680), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n651), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n552), .A2(new_n702), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n701), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n697), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n700), .A2(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n213), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G1), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT96), .ZN(new_n713));
  OAI22_X1  g0513(.A1(new_n712), .A2(new_n713), .B1(new_n230), .B2(new_n710), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n713), .B2(new_n712), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n715), .B(KEYINPUT28), .Z(new_n716));
  NAND4_X1  g0516(.A1(new_n656), .A2(new_n629), .A3(new_n663), .A4(new_n634), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n661), .A2(new_n662), .A3(new_n640), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n659), .B(new_n717), .C1(new_n718), .C2(new_n663), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n646), .A2(new_n647), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n641), .B1(new_n654), .B2(new_n720), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT29), .B(new_n682), .C1(new_n719), .C2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n682), .B1(new_n655), .B2(new_n665), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n724), .B2(KEYINPUT29), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n324), .A2(new_n635), .A3(new_n552), .A4(new_n682), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n597), .A2(new_n631), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n727), .A2(new_n547), .A3(KEYINPUT30), .A4(new_n278), .ZN(new_n728));
  XNOR2_X1  g0528(.A(KEYINPUT97), .B(KEYINPUT30), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n565), .A2(new_n566), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n278), .A2(new_n731), .A3(new_n617), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n730), .B1(new_n732), .B2(new_n546), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n526), .A2(new_n402), .A3(new_n631), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n731), .B1(new_n278), .B2(new_n282), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT98), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n316), .A2(new_n736), .A3(new_n597), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n728), .B(new_n733), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n680), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT31), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n726), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n680), .A2(KEYINPUT31), .ZN(new_n744));
  INV_X1    g0544(.A(new_n728), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n733), .B1(new_n737), .B2(new_n738), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n745), .B1(new_n746), .B2(KEYINPUT99), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT99), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n748), .B(new_n733), .C1(new_n737), .C2(new_n738), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n744), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(G330), .B1(new_n743), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n725), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n716), .B1(new_n753), .B2(G1), .ZN(G364));
  INV_X1    g0554(.A(new_n705), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n703), .A2(new_n701), .A3(new_n704), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n527), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n209), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n709), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n755), .A2(new_n756), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G13), .A2(G33), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n703), .A2(new_n704), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n708), .A2(new_n395), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n767), .A2(G355), .B1(new_n530), .B2(new_n708), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n708), .A2(new_n258), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(G45), .B2(new_n230), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n248), .A2(new_n266), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n768), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n226), .B1(G20), .B2(new_n374), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n765), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n761), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT100), .Z(new_n776));
  NOR2_X1   g0576(.A1(new_n210), .A2(G190), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G179), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G159), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT32), .Z(new_n782));
  NAND2_X1  g0582(.A1(new_n778), .A2(G190), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G20), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G97), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n210), .A2(new_n408), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n402), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n395), .B1(new_n789), .B2(G58), .ZN(new_n790));
  AND3_X1   g0590(.A1(new_n782), .A2(new_n785), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n311), .A2(G179), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT101), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n786), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G87), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n402), .A2(new_n311), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n786), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n797), .A2(new_n777), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G50), .A2(new_n799), .B1(new_n801), .B2(G68), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n777), .A2(new_n787), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n326), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n793), .A2(new_n777), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n804), .B1(G107), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n791), .A2(new_n796), .A3(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G283), .A2(new_n806), .B1(new_n795), .B2(G303), .ZN(new_n809));
  INV_X1    g0609(.A(G326), .ZN(new_n810));
  INV_X1    g0610(.A(G322), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n798), .A2(new_n810), .B1(new_n788), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G329), .B2(new_n780), .ZN(new_n813));
  INV_X1    g0613(.A(G311), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n395), .B1(new_n803), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(G294), .B2(new_n784), .ZN(new_n816));
  XNOR2_X1  g0616(.A(KEYINPUT33), .B(G317), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n800), .B1(new_n818), .B2(KEYINPUT102), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(KEYINPUT102), .B2(new_n818), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n809), .A2(new_n813), .A3(new_n816), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n808), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n776), .B1(new_n773), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n766), .A2(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n762), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  INV_X1    g0626(.A(KEYINPUT105), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n401), .A2(new_n403), .A3(new_n682), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n390), .A2(new_n682), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n409), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n827), .B(new_n828), .C1(new_n830), .C2(new_n669), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n409), .A2(new_n829), .B1(new_n401), .B2(new_n403), .ZN(new_n832));
  INV_X1    g0632(.A(new_n828), .ZN(new_n833));
  OAI21_X1  g0633(.A(KEYINPUT105), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n723), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n682), .B(new_n835), .C1(new_n655), .C2(new_n665), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n839), .A2(new_n751), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n760), .B1(new_n839), .B2(new_n751), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n836), .A2(new_n763), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n773), .A2(new_n763), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n760), .B1(G77), .B2(new_n845), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT103), .Z(new_n847));
  INV_X1    g0647(.A(new_n803), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G143), .A2(new_n789), .B1(new_n848), .B2(G159), .ZN(new_n849));
  INV_X1    g0649(.A(G137), .ZN(new_n850));
  INV_X1    g0650(.A(G150), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n849), .B1(new_n850), .B2(new_n798), .C1(new_n851), .C2(new_n800), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT34), .Z(new_n853));
  NAND2_X1  g0653(.A1(new_n795), .A2(G50), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n806), .A2(G68), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n784), .A2(G58), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n395), .B1(new_n780), .B2(G132), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G294), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n395), .B1(new_n779), .B2(new_n814), .C1(new_n859), .C2(new_n788), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(G97), .B2(new_n784), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n861), .B1(new_n219), .B2(new_n805), .C1(new_n206), .C2(new_n794), .ZN(new_n862));
  INV_X1    g0662(.A(G283), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n800), .A2(new_n863), .B1(new_n803), .B2(new_n530), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(G303), .B2(new_n799), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT104), .Z(new_n866));
  OAI22_X1  g0666(.A1(new_n853), .A2(new_n858), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n847), .B1(new_n867), .B2(new_n773), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n843), .A2(new_n868), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n842), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(G384));
  XOR2_X1   g0671(.A(new_n590), .B(KEYINPUT106), .Z(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n530), .B(new_n228), .C1(new_n873), .C2(KEYINPUT35), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(KEYINPUT35), .B2(new_n873), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n875), .B(KEYINPUT36), .Z(new_n876));
  AOI211_X1 g0676(.A(new_n326), .B(new_n230), .C1(G58), .C2(G68), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n877), .A2(KEYINPUT107), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n877), .A2(KEYINPUT107), .B1(new_n202), .B2(G68), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n209), .B(G13), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n496), .B1(KEYINPUT16), .B2(new_n495), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n678), .B1(new_n882), .B2(new_n470), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n509), .A2(new_n883), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n882), .A2(new_n470), .B1(new_n502), .B2(new_n678), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n468), .A2(new_n470), .A3(new_n489), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT37), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n504), .A2(new_n506), .ZN(new_n888));
  INV_X1    g0688(.A(new_n678), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n504), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT37), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n888), .A2(new_n890), .A3(new_n891), .A4(new_n490), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n884), .A2(KEYINPUT38), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n884), .B2(new_n893), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT39), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n884), .A2(new_n893), .A3(KEYINPUT38), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n888), .A2(new_n890), .A3(new_n490), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT37), .ZN(new_n900));
  INV_X1    g0700(.A(new_n890), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n900), .A2(new_n892), .B1(new_n509), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n898), .B1(new_n902), .B2(KEYINPUT38), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n897), .B1(KEYINPUT39), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n668), .A2(new_n682), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n347), .A2(new_n680), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n379), .A2(new_n382), .A3(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n347), .B(new_n680), .C1(new_n377), .C2(new_n378), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n838), .B2(new_n828), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n894), .B2(new_n895), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n513), .A2(new_n889), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n907), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n515), .B(new_n722), .C1(new_n724), .C2(KEYINPUT29), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n674), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n915), .B(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT108), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n726), .A2(new_n742), .A3(new_n920), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n909), .A2(new_n910), .B1(new_n831), .B2(new_n834), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT40), .B1(new_n904), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n884), .A2(new_n893), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT38), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT40), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(new_n928), .A3(new_n898), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n919), .A2(new_n928), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n929), .A2(new_n921), .A3(new_n922), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n924), .A2(new_n932), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n933), .A2(new_n515), .A3(new_n921), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n933), .B1(new_n515), .B2(new_n921), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n934), .A2(new_n935), .A3(new_n701), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n918), .A2(new_n936), .B1(new_n209), .B2(new_n757), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n918), .A2(new_n936), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n881), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT109), .ZN(G367));
  INV_X1    g0740(.A(new_n659), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n630), .A2(new_n680), .ZN(new_n942));
  MUX2_X1   g0742(.A(new_n941), .B(new_n640), .S(new_n942), .Z(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n588), .B(new_n599), .C1(new_n595), .C2(new_n682), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n656), .A2(new_n680), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n697), .A2(new_n705), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT110), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT94), .B1(new_n695), .B2(new_n684), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n691), .B(new_n683), .C1(new_n694), .C2(new_n688), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n699), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n948), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT42), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT42), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n697), .A2(new_n958), .A3(new_n699), .A4(new_n948), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n588), .B1(new_n946), .B2(new_n654), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n682), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n957), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n951), .B1(new_n952), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n952), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n949), .B(KEYINPUT110), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n945), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n964), .A2(new_n965), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n951), .A2(new_n952), .A3(new_n962), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(new_n969), .A3(new_n944), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n709), .B(KEYINPUT41), .Z(new_n972));
  INV_X1    g0772(.A(new_n681), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n955), .A2(KEYINPUT45), .A3(new_n973), .A4(new_n948), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT45), .B1(new_n700), .B2(new_n948), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n955), .A2(new_n973), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT44), .B1(new_n977), .B2(new_n956), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT44), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n979), .B(new_n948), .C1(new_n955), .C2(new_n973), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n975), .A2(new_n976), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n706), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n979), .B1(new_n700), .B2(new_n948), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n977), .A2(KEYINPUT44), .A3(new_n956), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n955), .A2(new_n973), .A3(new_n948), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT45), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n974), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n706), .A3(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n697), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n755), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n993), .A2(new_n706), .A3(new_n699), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n699), .B1(new_n993), .B2(new_n706), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n995), .A2(new_n996), .A3(new_n752), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n983), .A2(new_n991), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n972), .B1(new_n998), .B2(new_n753), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n971), .B1(new_n999), .B2(new_n759), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n774), .B1(new_n213), .B2(new_n384), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n769), .B2(new_n241), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n784), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(new_n217), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n395), .B(new_n1004), .C1(G143), .C2(new_n799), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G58), .A2(new_n795), .B1(new_n806), .B2(G77), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(G50), .A2(new_n848), .B1(new_n780), .B2(G137), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G150), .A2(new_n789), .B1(new_n801), .B2(G159), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n794), .A2(new_n530), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT46), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n806), .A2(G97), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n799), .A2(G311), .B1(new_n780), .B2(G317), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G303), .A2(new_n789), .B1(new_n848), .B2(G283), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n395), .B1(new_n800), .B2(new_n859), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G107), .B2(new_n784), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1009), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT47), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n761), .B(new_n1002), .C1(new_n1019), .C2(new_n773), .ZN(new_n1020));
  OR3_X1    g0820(.A1(new_n943), .A2(G20), .A3(new_n764), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1000), .A2(new_n1022), .ZN(G387));
  NOR2_X1   g0823(.A1(new_n995), .A2(new_n996), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n992), .A2(new_n765), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n238), .A2(G45), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT111), .Z(new_n1027));
  XOR2_X1   g0827(.A(KEYINPUT8), .B(G58), .Z(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n202), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT50), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n711), .B(new_n266), .C1(new_n217), .C2(new_n326), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1027), .B(new_n769), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n711), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n767), .A2(new_n1033), .B1(new_n206), .B2(new_n708), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n765), .B(new_n773), .C1(new_n1032), .C2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1003), .A2(new_n384), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G50), .B2(new_n789), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT112), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n258), .B1(new_n779), .B2(new_n851), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n800), .A2(new_n385), .B1(new_n803), .B2(new_n217), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(G159), .C2(new_n799), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n795), .A2(G77), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1038), .A2(new_n1012), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n795), .A2(G294), .B1(G283), .B2(new_n784), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G317), .A2(new_n789), .B1(new_n848), .B2(G303), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n814), .B2(new_n800), .C1(new_n811), .C2(new_n798), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT48), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n1047), .B2(new_n1046), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(KEYINPUT49), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n258), .B1(new_n780), .B2(G326), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(new_n530), .C2(new_n805), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1049), .A2(KEYINPUT49), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1043), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n761), .B(new_n1035), .C1(new_n1054), .C2(new_n773), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n1024), .A2(new_n759), .B1(new_n1025), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n996), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1057), .A2(new_n753), .A3(new_n994), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n709), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1024), .A2(new_n753), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1056), .B1(new_n1059), .B2(new_n1060), .ZN(G393));
  AND3_X1   g0861(.A1(new_n986), .A2(new_n706), .A3(new_n990), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n706), .B1(new_n986), .B2(new_n990), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n956), .A2(new_n765), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n769), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n774), .B1(new_n205), .B2(new_n213), .C1(new_n1066), .C2(new_n245), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n760), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT52), .ZN(new_n1069));
  INV_X1    g0869(.A(G317), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n798), .A2(new_n1070), .B1(new_n788), .B2(new_n814), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n795), .A2(G283), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n1069), .B2(new_n1071), .C1(new_n206), .C2(new_n805), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G294), .A2(new_n848), .B1(new_n780), .B2(G322), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n258), .B1(new_n801), .B2(G303), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(new_n530), .C2(new_n1003), .ZN(new_n1076));
  INV_X1    g0876(.A(G159), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n798), .A2(new_n851), .B1(new_n788), .B2(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1078), .B(new_n1079), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1080), .B1(new_n217), .B2(new_n794), .C1(new_n219), .C2(new_n805), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G50), .A2(new_n801), .B1(new_n848), .B2(new_n1028), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n395), .B1(new_n780), .B2(G143), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1082), .B(new_n1083), .C1(new_n326), .C2(new_n1003), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n1073), .A2(new_n1076), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1068), .B1(new_n1085), .B2(new_n773), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1064), .A2(new_n759), .B1(new_n1065), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1058), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1088), .A2(new_n998), .A3(new_n709), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(G390));
  NAND2_X1  g0890(.A1(new_n905), .A2(new_n763), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n760), .B1(new_n1028), .B2(new_n845), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n395), .B1(new_n800), .B2(new_n206), .C1(new_n1003), .C2(new_n326), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n788), .A2(new_n530), .B1(new_n803), .B2(new_n205), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n798), .A2(new_n863), .B1(new_n779), .B2(new_n859), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1096), .A2(new_n796), .A3(new_n855), .ZN(new_n1097));
  INV_X1    g0897(.A(G132), .ZN(new_n1098));
  INV_X1    g0898(.A(G125), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n788), .A2(new_n1098), .B1(new_n779), .B2(new_n1099), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n395), .B(new_n1100), .C1(G128), .C2(new_n799), .ZN(new_n1101));
  OR3_X1    g0901(.A1(new_n794), .A2(KEYINPUT53), .A3(new_n851), .ZN(new_n1102));
  OAI21_X1  g0902(.A(KEYINPUT53), .B1(new_n794), .B2(new_n851), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n784), .A2(G159), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT54), .B(G143), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n800), .A2(new_n850), .B1(new_n803), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n806), .A2(G50), .B1(new_n1108), .B2(KEYINPUT114), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(KEYINPUT114), .B2(new_n1108), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1097), .B1(new_n1105), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1092), .B1(new_n1111), .B2(new_n773), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1091), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n900), .A2(new_n892), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n509), .A2(new_n901), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n926), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT39), .B1(new_n1117), .B2(new_n898), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT39), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n894), .A2(new_n895), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n906), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n1118), .A2(new_n1120), .B1(new_n912), .B2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n682), .B(new_n835), .C1(new_n719), .C2(new_n721), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1123), .A2(new_n828), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n906), .B(new_n903), .C1(new_n1124), .C2(new_n911), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n922), .B(G330), .C1(new_n743), .C2(new_n750), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1122), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n921), .A2(G330), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n922), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1113), .B1(new_n1131), .B2(new_n758), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(KEYINPUT115), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1128), .A2(new_n515), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n916), .A2(new_n674), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n921), .A2(G330), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n911), .B1(new_n1136), .B2(new_n836), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1137), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n838), .A2(new_n828), .ZN(new_n1140));
  OAI211_X1 g0940(.A(G330), .B(new_n835), .C1(new_n743), .C2(new_n750), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n911), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1140), .B1(new_n1129), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1135), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1131), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1144), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1145), .A2(new_n1148), .A3(new_n709), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT115), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1150), .B(new_n1113), .C1(new_n1131), .C2(new_n758), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1133), .A2(new_n1149), .A3(new_n1151), .ZN(G378));
  NAND2_X1  g0952(.A1(new_n921), .A2(new_n922), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(KEYINPUT108), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n928), .B1(new_n1154), .B2(new_n903), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n921), .A2(new_n922), .A3(new_n931), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n896), .B2(new_n928), .ZN(new_n1157));
  OAI21_X1  g0957(.A(G330), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(KEYINPUT119), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT119), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1160), .B(G330), .C1(new_n1155), .C2(new_n1157), .ZN(new_n1161));
  XOR2_X1   g0961(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1162));
  XNOR2_X1  g0962(.A(new_n450), .B(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n428), .A2(new_n678), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT118), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1163), .B(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1159), .A2(new_n1161), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1161), .A2(new_n1167), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1160), .B1(new_n933), .B2(G330), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n907), .A2(new_n913), .A3(new_n914), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1168), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1172), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n759), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(G50), .B1(new_n255), .B2(new_n261), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1004), .B1(G116), .B2(new_n799), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT116), .Z(new_n1178));
  OAI211_X1 g0978(.A(new_n261), .B(new_n395), .C1(new_n779), .C2(new_n863), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n788), .A2(new_n206), .B1(new_n803), .B2(new_n384), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(G97), .C2(new_n801), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n806), .A2(G58), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1178), .A2(new_n1042), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT58), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1176), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n800), .A2(new_n1098), .B1(new_n803), .B2(new_n850), .ZN(new_n1186));
  INV_X1    g0986(.A(G128), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n798), .A2(new_n1099), .B1(new_n788), .B2(new_n1187), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1186), .B(new_n1188), .C1(G150), .C2(new_n784), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n794), .B2(new_n1106), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1190), .B(new_n1191), .ZN(new_n1192));
  AOI211_X1 g0992(.A(G33), .B(G41), .C1(new_n780), .C2(G124), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n1077), .B2(new_n805), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1185), .B1(new_n1184), .B2(new_n1183), .C1(new_n1192), .C2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n773), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n761), .B1(new_n202), .B2(new_n844), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(new_n1166), .C2(new_n764), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1175), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1148), .A2(new_n1135), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT57), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n710), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1158), .A2(KEYINPUT119), .A3(new_n1166), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n915), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT120), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1168), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n915), .B(KEYINPUT120), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n916), .A2(new_n674), .A3(new_n1134), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1212), .A2(new_n1202), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1209), .A2(new_n1210), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1199), .B1(new_n1203), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(G375));
  OAI21_X1  g1016(.A(new_n759), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n911), .A2(new_n763), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT122), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n258), .B(new_n1036), .C1(G303), .C2(new_n780), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G77), .A2(new_n806), .B1(new_n795), .B2(G97), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G116), .A2(new_n801), .B1(new_n848), .B2(G107), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G294), .A2(new_n799), .B1(new_n789), .B2(G283), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n788), .A2(new_n850), .B1(new_n779), .B2(new_n1187), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n799), .A2(G132), .B1(new_n848), .B2(G150), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n800), .B2(new_n1106), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1225), .B(new_n1227), .C1(G50), .C2(new_n784), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1182), .A2(new_n258), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT123), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(new_n1077), .C2(new_n794), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1229), .A2(KEYINPUT123), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1224), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n773), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n761), .B1(new_n217), .B2(new_n844), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1219), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1217), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1129), .A2(new_n1142), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1211), .B(new_n1138), .C1(new_n1239), .C2(new_n1140), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT121), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1143), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT121), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1242), .A2(new_n1243), .A3(new_n1211), .A4(new_n1138), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n972), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1144), .A2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1238), .B1(new_n1245), .B2(new_n1247), .ZN(G381));
  INV_X1    g1048(.A(G378), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1215), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(G390), .ZN(new_n1251));
  NOR4_X1   g1051(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  OR3_X1    g1053(.A1(new_n1250), .A2(G387), .A3(new_n1253), .ZN(G407));
  NAND2_X1  g1054(.A1(new_n679), .A2(G213), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(KEYINPUT124), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G407), .B(G213), .C1(new_n1250), .C2(new_n1257), .ZN(G409));
  XNOR2_X1  g1058(.A(G393), .B(new_n825), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1000), .A2(new_n1022), .A3(G390), .ZN(new_n1261));
  AOI21_X1  g1061(.A(G390), .B1(new_n1000), .B2(new_n1022), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1260), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n967), .A2(new_n970), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1062), .A2(new_n1063), .A3(new_n1058), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1246), .B1(new_n1265), .B2(new_n752), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1264), .B1(new_n1266), .B2(new_n758), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1022), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1251), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1000), .A2(new_n1022), .A3(G390), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(new_n1259), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1263), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1144), .A2(KEYINPUT60), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(new_n1241), .A3(new_n1244), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1240), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n710), .B1(new_n1275), .B2(KEYINPUT60), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G384), .B1(new_n1277), .B2(new_n1238), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n870), .B(new_n1237), .C1(new_n1274), .C2(new_n1276), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT61), .B1(new_n1281), .B2(KEYINPUT62), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1198), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1212), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1283), .B1(new_n1284), .B2(new_n1246), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1209), .A2(new_n759), .A3(new_n1210), .ZN(new_n1286));
  AOI21_X1  g1086(.A(G378), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1215), .B2(G378), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1288), .A2(new_n1256), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1278), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1279), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1255), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(G2897), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1290), .A2(new_n1291), .A3(new_n1293), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1256), .A2(G2897), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1295), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT125), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1294), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(KEYINPUT125), .B(new_n1295), .C1(new_n1278), .C2(new_n1279), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1300), .A2(KEYINPUT62), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1282), .B1(new_n1289), .B2(new_n1301), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1175), .A2(new_n1198), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1214), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n709), .B1(new_n1284), .B2(KEYINPUT57), .ZN(new_n1305));
  OAI211_X1 g1105(.A(G378), .B(new_n1303), .C1(new_n1304), .C2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1198), .B1(new_n1201), .B2(new_n972), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1209), .A2(new_n759), .A3(new_n1210), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1249), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1292), .B1(new_n1306), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1280), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1311), .A2(KEYINPUT62), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1272), .B1(new_n1302), .B2(new_n1312), .ZN(new_n1313));
  AOI211_X1 g1113(.A(new_n1292), .B(new_n1281), .C1(new_n1306), .C2(new_n1309), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1300), .B1(new_n1288), .B2(new_n1292), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1314), .B1(new_n1315), .B2(KEYINPUT63), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1306), .A2(new_n1309), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1280), .A2(KEYINPUT63), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1317), .A2(new_n1257), .A3(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT61), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1320), .A2(new_n1321), .A3(new_n1271), .A4(new_n1263), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1316), .A2(new_n1322), .A3(KEYINPUT126), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT126), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1263), .A2(new_n1271), .A3(new_n1321), .ZN(new_n1325));
  AOI211_X1 g1125(.A(new_n1256), .B(new_n1318), .C1(new_n1306), .C2(new_n1309), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1299), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT125), .B1(new_n1280), .B2(new_n1293), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1328), .B1(new_n1329), .B2(new_n1296), .ZN(new_n1330));
  OAI21_X1  g1130(.A(KEYINPUT63), .B1(new_n1310), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1311), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1324), .B1(new_n1327), .B2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1313), .B1(new_n1323), .B2(new_n1333), .ZN(G405));
  NAND2_X1  g1134(.A1(new_n1281), .A2(KEYINPUT127), .ZN(new_n1335));
  AND3_X1   g1135(.A1(new_n1263), .A2(new_n1271), .A3(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1335), .B1(new_n1263), .B2(new_n1271), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(G375), .A2(new_n1249), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1339), .B(new_n1306), .C1(KEYINPUT127), .C2(new_n1281), .ZN(new_n1340));
  XNOR2_X1  g1140(.A(new_n1338), .B(new_n1340), .ZN(G402));
endmodule


