//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT69), .B(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G210), .A3(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(G101), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G113), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT2), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G113), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G116), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G119), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G116), .ZN(new_n202));
  INV_X1    g016(.A(G119), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n198), .B(new_n201), .C1(new_n202), .C2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT67), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(KEYINPUT66), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G116), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G119), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n210), .A2(new_n211), .A3(new_n201), .A4(new_n198), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n201), .B1(new_n202), .B2(new_n203), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT2), .B(G113), .ZN(new_n214));
  AOI22_X1  g028(.A1(new_n205), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G134), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT11), .B1(new_n216), .B2(G137), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT11), .ZN(new_n218));
  INV_X1    g032(.A(G137), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(G134), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n216), .A2(G137), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n226), .B1(new_n216), .B2(G137), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n223), .A2(new_n225), .ZN(new_n228));
  OAI21_X1  g042(.A(G131), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G143), .ZN(new_n231));
  INV_X1    g045(.A(G143), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G146), .ZN(new_n233));
  INV_X1    g047(.A(G128), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT65), .B(KEYINPUT1), .Z(new_n237));
  XNOR2_X1  g051(.A(G143), .B(G146), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n236), .B1(new_n239), .B2(G128), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n237), .A2(new_n233), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n224), .B(new_n229), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n232), .A2(G146), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n230), .A2(G143), .ZN(new_n245));
  OAI21_X1  g059(.A(G128), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(KEYINPUT0), .A3(new_n235), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n231), .A2(new_n233), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT0), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(G128), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n218), .B1(G134), .B2(new_n219), .ZN(new_n252));
  NOR3_X1   g066(.A1(new_n216), .A2(KEYINPUT11), .A3(G137), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n223), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G131), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n224), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n243), .B1(new_n251), .B2(new_n256), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n222), .B1(new_n221), .B2(new_n223), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n247), .A2(new_n250), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT68), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n215), .B(new_n242), .C1(new_n257), .C2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n256), .A2(new_n250), .A3(new_n247), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT30), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n242), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n242), .B1(new_n257), .B2(new_n262), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(KEYINPUT30), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n193), .B(new_n263), .C1(new_n268), .C2(new_n215), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n272));
  OAI21_X1  g086(.A(G128), .B1(new_n248), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n235), .ZN(new_n274));
  INV_X1    g088(.A(new_n241), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n258), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n276), .A2(new_n229), .B1(new_n251), .B2(new_n256), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n265), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT68), .B1(new_n260), .B2(new_n261), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n251), .A2(new_n243), .A3(new_n256), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n279), .A2(new_n280), .B1(new_n229), .B2(new_n276), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n278), .B1(new_n281), .B2(new_n265), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n213), .A2(new_n214), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n200), .B1(new_n209), .B2(G119), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n211), .B1(new_n284), .B2(new_n198), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n203), .B1(new_n206), .B2(new_n208), .ZN(new_n286));
  NOR4_X1   g100(.A1(new_n286), .A2(new_n214), .A3(KEYINPUT67), .A4(new_n200), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n283), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n289), .A2(KEYINPUT70), .A3(new_n193), .A4(new_n263), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n271), .A2(KEYINPUT31), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT31), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n269), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT28), .B1(new_n277), .B2(new_n215), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT71), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n297), .B1(new_n277), .B2(new_n215), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n242), .A2(new_n264), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(KEYINPUT71), .A3(new_n288), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n263), .A3(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n301), .A2(KEYINPUT72), .A3(KEYINPUT28), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT72), .B1(new_n301), .B2(KEYINPUT28), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n296), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n193), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n294), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(G472), .A2(G902), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n187), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n291), .A2(new_n293), .B1(new_n304), .B2(new_n305), .ZN(new_n310));
  INV_X1    g124(.A(new_n308), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n310), .A2(KEYINPUT32), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n193), .B(new_n296), .C1(new_n302), .C2(new_n303), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n315));
  INV_X1    g129(.A(new_n263), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n316), .B1(new_n282), .B2(new_n288), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n315), .B1(new_n317), .B2(new_n193), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n279), .A2(new_n280), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n215), .B1(new_n321), .B2(new_n242), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT28), .B1(new_n316), .B2(new_n322), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n323), .A2(KEYINPUT29), .A3(new_n193), .A4(new_n296), .ZN(new_n324));
  INV_X1    g138(.A(G902), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n320), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n313), .B1(new_n328), .B2(G472), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n326), .B1(new_n314), .B2(new_n319), .ZN(new_n330));
  INV_X1    g144(.A(G472), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n330), .A2(KEYINPUT73), .A3(new_n331), .ZN(new_n332));
  OAI22_X1  g146(.A1(new_n309), .A2(new_n312), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(G214), .B1(G237), .B2(G902), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n241), .B1(new_n235), .B2(new_n273), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT86), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n336), .A2(KEYINPUT86), .A3(new_n337), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G224), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(G953), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n261), .A2(G125), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n342), .A2(KEYINPUT7), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G107), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(G104), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(G104), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n349), .B1(KEYINPUT3), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT3), .ZN(new_n352));
  AND2_X1   g166(.A1(KEYINPUT82), .A2(G107), .ZN(new_n353));
  NOR2_X1   g167(.A1(KEYINPUT82), .A2(G107), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n352), .B(G104), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT4), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(G101), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(G101), .ZN(new_n359));
  INV_X1    g173(.A(G101), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n351), .A2(new_n360), .A3(new_n355), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(KEYINPUT4), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n288), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT83), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n348), .ZN(new_n366));
  INV_X1    g180(.A(G104), .ZN(new_n367));
  NAND2_X1  g181(.A1(KEYINPUT82), .A2(G107), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n350), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n364), .B1(new_n370), .B2(G101), .ZN(new_n371));
  AOI211_X1 g185(.A(KEYINPUT83), .B(new_n360), .C1(new_n369), .C2(new_n350), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n205), .A2(new_n212), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT5), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n200), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(G113), .B(new_n376), .C1(new_n213), .C2(new_n375), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n373), .A2(new_n374), .A3(new_n361), .A4(new_n377), .ZN(new_n378));
  XOR2_X1   g192(.A(G110), .B(G122), .Z(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n363), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n340), .A2(new_n346), .A3(new_n341), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT7), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n382), .B1(new_n383), .B2(new_n344), .ZN(new_n384));
  INV_X1    g198(.A(new_n350), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n353), .A2(new_n354), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n385), .B1(new_n386), .B2(new_n367), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT83), .B1(new_n387), .B2(new_n360), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n370), .A2(new_n364), .A3(G101), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n388), .A2(new_n389), .A3(new_n361), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n374), .A2(new_n377), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT87), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n388), .A2(new_n389), .A3(new_n361), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT87), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n374), .B(new_n377), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  XOR2_X1   g209(.A(new_n379), .B(KEYINPUT8), .Z(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n347), .A2(new_n381), .A3(new_n384), .A4(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n362), .A2(new_n358), .ZN(new_n399));
  OAI22_X1  g213(.A1(new_n399), .A2(new_n215), .B1(new_n391), .B2(new_n393), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT85), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n400), .A2(new_n379), .B1(new_n401), .B2(KEYINPUT6), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(KEYINPUT6), .ZN(new_n403));
  AOI211_X1 g217(.A(new_n380), .B(new_n403), .C1(new_n363), .C2(new_n378), .ZN(new_n404));
  INV_X1    g218(.A(new_n381), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n382), .B(new_n345), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n325), .B(new_n398), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G210), .B1(G237), .B2(G902), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n407), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n400), .A2(new_n379), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n403), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT6), .A4(new_n379), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n381), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n417), .A2(new_n325), .A3(new_n409), .A4(new_n398), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n335), .B1(new_n411), .B2(new_n418), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n189), .A2(G952), .ZN(new_n420));
  NAND2_X1  g234(.A1(G234), .A2(G237), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  XOR2_X1   g237(.A(KEYINPUT21), .B(G898), .Z(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n421), .A2(G902), .A3(G953), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n423), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n419), .A2(new_n429), .ZN(new_n430));
  AND2_X1   g244(.A1(KEYINPUT69), .A2(G237), .ZN(new_n431));
  NOR2_X1   g245(.A1(KEYINPUT69), .A2(G237), .ZN(new_n432));
  OAI211_X1 g246(.A(G214), .B(new_n189), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n232), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n188), .A2(G143), .A3(G214), .A4(new_n189), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G131), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT17), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n434), .A2(new_n435), .A3(new_n222), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  XOR2_X1   g254(.A(G125), .B(G140), .Z(new_n441));
  INV_X1    g255(.A(KEYINPUT16), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(G125), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(G140), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n230), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(G125), .B(G140), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n445), .B1(new_n447), .B2(KEYINPUT16), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G146), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n222), .B1(new_n434), .B2(new_n435), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT17), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n440), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n436), .A2(KEYINPUT18), .A3(G131), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT88), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n447), .B(G146), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n434), .A2(new_n435), .ZN(new_n458));
  NAND2_X1  g272(.A1(KEYINPUT18), .A2(G131), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n451), .A2(KEYINPUT88), .A3(KEYINPUT18), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n456), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n453), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G113), .B(G122), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(new_n367), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n453), .A2(new_n462), .A3(new_n465), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n325), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G475), .ZN(new_n471));
  NOR2_X1   g285(.A1(G475), .A2(G902), .ZN(new_n472));
  XOR2_X1   g286(.A(new_n472), .B(KEYINPUT89), .Z(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n453), .A2(new_n462), .A3(new_n465), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n437), .A2(new_n439), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n441), .A2(KEYINPUT19), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n441), .A2(KEYINPUT19), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n230), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n476), .A2(new_n449), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n465), .B1(new_n462), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n474), .B1(new_n475), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT90), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT20), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT20), .B1(new_n482), .B2(new_n483), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n462), .A2(new_n480), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n466), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n473), .B1(new_n488), .B2(new_n468), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(KEYINPUT90), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n471), .B(new_n485), .C1(new_n486), .C2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(G128), .B(G143), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT13), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n232), .A2(G128), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n493), .B(G134), .C1(KEYINPUT13), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n216), .ZN(new_n496));
  INV_X1    g310(.A(new_n386), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n209), .A2(G122), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n199), .A2(G122), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n497), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G122), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n502), .B1(new_n206), .B2(new_n208), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n503), .A2(new_n386), .A3(new_n499), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n495), .B(new_n496), .C1(new_n501), .C2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT14), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n506), .B(new_n500), .C1(new_n202), .C2(new_n502), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n209), .A2(KEYINPUT14), .A3(G122), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(G107), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n498), .A2(new_n497), .A3(new_n500), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n492), .B(new_n216), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT9), .B(G234), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT81), .ZN(new_n515));
  INV_X1    g329(.A(G217), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n515), .A2(new_n516), .A3(G953), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n505), .A2(new_n512), .A3(new_n517), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(KEYINPUT91), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT91), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n505), .A2(new_n512), .A3(new_n517), .A4(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n325), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G478), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(KEYINPUT15), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n524), .B(new_n526), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n491), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G469), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n245), .A2(KEYINPUT1), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n274), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n531), .A2(new_n361), .A3(new_n388), .A4(new_n389), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT10), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n336), .A2(new_n533), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n390), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n362), .A2(new_n251), .A3(new_n358), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n534), .A2(new_n260), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(G110), .B(G140), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n189), .A2(G227), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n393), .A2(new_n336), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n532), .A3(KEYINPUT84), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT84), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n393), .A2(new_n545), .A3(new_n336), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n544), .A2(new_n256), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT12), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n544), .A2(KEYINPUT12), .A3(new_n256), .A4(new_n546), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n542), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n534), .A2(new_n537), .A3(new_n536), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n256), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n541), .B1(new_n553), .B2(new_n538), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n529), .B(new_n325), .C1(new_n551), .C2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n538), .A3(new_n541), .ZN(new_n556));
  INV_X1    g370(.A(new_n538), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(new_n549), .B2(new_n550), .ZN(new_n558));
  OAI211_X1 g372(.A(G469), .B(new_n556), .C1(new_n558), .C2(new_n541), .ZN(new_n559));
  NAND2_X1  g373(.A1(G469), .A2(G902), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n555), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G221), .ZN(new_n562));
  INV_X1    g376(.A(new_n515), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n562), .B1(new_n563), .B2(new_n325), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n430), .A2(new_n528), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n441), .A2(G146), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n448), .B2(G146), .ZN(new_n569));
  OR3_X1    g383(.A1(new_n203), .A2(KEYINPUT78), .A3(G128), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n234), .A2(G119), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT78), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT77), .B(KEYINPUT23), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n234), .A2(G119), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n570), .B(new_n572), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n234), .A2(KEYINPUT23), .A3(G119), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT76), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XOR2_X1   g392(.A(KEYINPUT79), .B(G110), .Z(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT80), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n575), .A2(new_n578), .A3(KEYINPUT80), .A4(new_n579), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT24), .B(G110), .Z(new_n585));
  NAND2_X1  g399(.A1(new_n203), .A2(G128), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n571), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT74), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT74), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n571), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n585), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n569), .B1(new_n584), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n588), .A2(new_n590), .A3(new_n585), .ZN(new_n593));
  XOR2_X1   g407(.A(new_n593), .B(KEYINPUT75), .Z(new_n594));
  NAND2_X1  g408(.A1(new_n575), .A2(new_n578), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n446), .A2(new_n449), .B1(new_n595), .B2(G110), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT22), .B(G137), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n599), .B(new_n600), .Z(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n592), .A2(new_n597), .A3(new_n601), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(new_n325), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT25), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n516), .B1(G234), .B2(new_n325), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT25), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n603), .A2(new_n608), .A3(new_n325), .A4(new_n604), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  OR2_X1    g424(.A1(new_n605), .A2(new_n607), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n333), .A2(new_n567), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G101), .ZN(G3));
  AND3_X1   g428(.A1(new_n612), .A2(new_n561), .A3(new_n565), .ZN(new_n615));
  OAI21_X1  g429(.A(G472), .B1(new_n310), .B2(G902), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n307), .A2(new_n308), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT92), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n430), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n615), .A2(new_n616), .A3(new_n617), .A4(KEYINPUT92), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(G475), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n469), .B2(new_n325), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n484), .B1(new_n489), .B2(KEYINPUT90), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n482), .A2(new_n483), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n521), .A2(new_n629), .A3(new_n523), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n525), .A2(G902), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n519), .A2(KEYINPUT33), .A3(new_n520), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT93), .B(G478), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n524), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT94), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT94), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n633), .A2(new_n638), .A3(new_n635), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n628), .A2(new_n485), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n623), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT95), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n642), .B(new_n644), .ZN(G6));
  INV_X1    g459(.A(new_n491), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n527), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n623), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT35), .B(G107), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NOR2_X1   g464(.A1(new_n607), .A2(G902), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n598), .A2(KEYINPUT96), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n602), .A2(KEYINPUT36), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n598), .A2(KEYINPUT96), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n653), .B1(new_n652), .B2(new_n654), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n610), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n567), .A2(new_n617), .A3(new_n616), .A4(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT97), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n659), .B(new_n661), .ZN(G12));
  INV_X1    g476(.A(new_n419), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n658), .A2(new_n561), .A3(new_n565), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n422), .B(KEYINPUT98), .Z(new_n666));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n666), .B1(new_n667), .B2(new_n427), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n647), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n333), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  INV_X1    g485(.A(new_n418), .ZN(new_n672));
  AOI21_X1  g486(.A(G902), .B1(new_n412), .B2(new_n416), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n409), .B1(new_n673), .B2(new_n398), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT38), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n307), .A2(new_n187), .A3(new_n308), .ZN(new_n678));
  OAI21_X1  g492(.A(KEYINPUT32), .B1(new_n310), .B2(new_n311), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n271), .A2(new_n290), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n316), .A2(new_n322), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n681), .B1(new_n305), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(G472), .B1(new_n683), .B2(G902), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n491), .A2(new_n527), .A3(new_n334), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n686), .A2(new_n658), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n687), .A2(KEYINPUT99), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(KEYINPUT99), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n677), .A2(new_n685), .A3(new_n688), .A4(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT100), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n668), .B(KEYINPUT39), .Z(new_n694));
  AND3_X1   g508(.A1(new_n561), .A2(new_n565), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT40), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n692), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G143), .ZN(G45));
  INV_X1    g512(.A(new_n668), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n419), .A2(new_n640), .A3(KEYINPUT101), .A4(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n664), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n637), .A2(new_n639), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n703), .A2(new_n491), .A3(new_n699), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT101), .B1(new_n704), .B2(new_n419), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n333), .A2(new_n702), .A3(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n301), .A2(KEYINPUT28), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT72), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n301), .A2(KEYINPUT72), .A3(KEYINPUT28), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n295), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n318), .B1(new_n714), .B2(new_n193), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n313), .B(G472), .C1(new_n715), .C2(new_n326), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT73), .B1(new_n330), .B2(new_n331), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n705), .B1(new_n680), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(KEYINPUT102), .A3(new_n702), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n709), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G146), .ZN(G48));
  OAI21_X1  g536(.A(new_n325), .B1(new_n551), .B2(new_n554), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(G469), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT103), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n725), .A3(new_n555), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n723), .A2(KEYINPUT103), .A3(G469), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n565), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n430), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n333), .A2(new_n730), .A3(new_n612), .A4(new_n640), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT41), .B(G113), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G15));
  INV_X1    g547(.A(new_n647), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n333), .A2(new_n730), .A3(new_n612), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G116), .ZN(G18));
  NOR2_X1   g550(.A1(new_n729), .A2(new_n663), .ZN(new_n737));
  INV_X1    g551(.A(new_n658), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n528), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n333), .A2(new_n737), .A3(new_n429), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  OR2_X1    g555(.A1(new_n675), .A2(new_n686), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n428), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n331), .B1(new_n307), .B2(new_n325), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n323), .A2(new_n296), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n305), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n311), .B1(new_n294), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n729), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n743), .A2(new_n748), .A3(new_n612), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(KEYINPUT104), .B(G122), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(G24));
  NOR3_X1   g566(.A1(new_n744), .A2(new_n738), .A3(new_n747), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n737), .A3(new_n704), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  XNOR2_X1  g569(.A(new_n560), .B(KEYINPUT105), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n555), .A2(new_n559), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n555), .A2(new_n559), .A3(KEYINPUT106), .A4(new_n756), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n565), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n411), .A2(new_n334), .A3(new_n418), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n333), .A2(new_n612), .A3(new_n704), .A4(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT42), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n640), .A2(new_n699), .ZN(new_n768));
  NOR4_X1   g582(.A1(new_n761), .A2(new_n768), .A3(new_n765), .A4(new_n762), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n678), .A2(new_n679), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n718), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n770), .B1(new_n678), .B2(new_n679), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n612), .B(new_n769), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n766), .A2(new_n767), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n767), .B1(new_n766), .B2(new_n774), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n222), .ZN(G33));
  NAND4_X1  g592(.A1(new_n333), .A2(new_n612), .A3(new_n669), .A4(new_n763), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G134), .ZN(G36));
  OAI21_X1  g594(.A(new_n556), .B1(new_n558), .B2(new_n541), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT45), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(G469), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT109), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(KEYINPUT109), .A3(G469), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(KEYINPUT46), .A3(new_n756), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n555), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT110), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT46), .ZN(new_n791));
  INV_X1    g605(.A(new_n787), .ZN(new_n792));
  INV_X1    g606(.A(new_n756), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n788), .A2(new_n795), .A3(new_n555), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n790), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n565), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n703), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n491), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT43), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n616), .A2(new_n617), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n803), .A3(new_n658), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT44), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n762), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n804), .A2(new_n805), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n799), .A2(new_n694), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G137), .ZN(G39));
  INV_X1    g624(.A(KEYINPUT47), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n798), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n797), .A2(KEYINPUT47), .A3(new_n565), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n678), .A2(new_n679), .B1(new_n716), .B2(new_n717), .ZN(new_n815));
  INV_X1    g629(.A(new_n612), .ZN(new_n816));
  INV_X1    g630(.A(new_n762), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n815), .A2(new_n816), .A3(new_n704), .A4(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT111), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(KEYINPUT112), .B(G140), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n820), .B(new_n821), .ZN(G42));
  XNOR2_X1  g636(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT102), .B1(new_n719), .B2(new_n702), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n700), .A2(new_n701), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n815), .A2(new_n825), .A3(new_n708), .A4(new_n705), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n670), .B(new_n754), .C1(new_n824), .C2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n742), .B1(new_n680), .B2(new_n684), .ZN(new_n828));
  INV_X1    g642(.A(new_n761), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n828), .A2(new_n738), .A3(new_n829), .A4(new_n699), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n823), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n670), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(new_n709), .B2(new_n720), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(KEYINPUT52), .A3(new_n754), .A4(new_n830), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n734), .A2(KEYINPUT113), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n647), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(new_n641), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n620), .A2(new_n841), .A3(new_n621), .A4(new_n622), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n613), .A3(new_n659), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n766), .B2(new_n774), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n731), .A2(new_n735), .A3(new_n750), .A4(new_n740), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n528), .A2(new_n668), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n333), .A2(new_n701), .A3(new_n817), .A4(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n753), .A2(new_n704), .A3(new_n763), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n779), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n844), .A2(new_n846), .A3(new_n847), .A4(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n836), .A2(new_n837), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n837), .B1(new_n836), .B2(new_n853), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n844), .A2(new_n847), .A3(new_n852), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT114), .B1(new_n777), .B2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n731), .A2(new_n735), .A3(new_n750), .A4(new_n740), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n860), .A2(new_n843), .A3(new_n851), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT114), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n861), .B(new_n862), .C1(new_n776), .C2(new_n775), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT52), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(new_n827), .B2(new_n831), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n835), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n859), .A2(new_n863), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n845), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n856), .A2(new_n857), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n867), .A2(KEYINPUT53), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n859), .A2(new_n863), .A3(new_n845), .A4(new_n836), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(KEYINPUT54), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  AND4_X1   g688(.A1(new_n612), .A2(new_n802), .A3(new_n666), .A4(new_n748), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n737), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n335), .A3(new_n676), .A4(new_n749), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT50), .Z(new_n878));
  NOR2_X1   g692(.A1(new_n729), .A2(new_n762), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n802), .A2(new_n879), .A3(new_n666), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT117), .Z(new_n881));
  NAND2_X1  g695(.A1(new_n612), .A2(new_n423), .ZN(new_n882));
  NOR4_X1   g696(.A1(new_n685), .A2(new_n729), .A3(new_n762), .A4(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n703), .A2(new_n491), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n881), .A2(new_n753), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n878), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n728), .A2(new_n564), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n812), .A2(new_n813), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT118), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n875), .A2(new_n817), .ZN(new_n890));
  OAI211_X1 g704(.A(KEYINPUT51), .B(new_n886), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n888), .A2(new_n817), .A3(new_n875), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT51), .B1(new_n892), .B2(new_n886), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n612), .B1(new_n772), .B2(new_n773), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n881), .A2(new_n895), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n896), .A2(KEYINPUT48), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(KEYINPUT48), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n883), .A2(new_n640), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n897), .A2(new_n420), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n893), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n874), .A2(new_n876), .A3(new_n891), .A4(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n902), .B1(G952), .B2(G953), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n677), .A2(new_n685), .A3(new_n816), .ZN(new_n904));
  NOR4_X1   g718(.A1(new_n800), .A2(new_n491), .A3(new_n564), .A4(new_n335), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n728), .B(KEYINPUT49), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n903), .A2(new_n907), .ZN(G75));
  XNOR2_X1  g722(.A(new_n416), .B(new_n407), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT55), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT56), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n911), .B1(KEYINPUT119), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(G210), .ZN(new_n915));
  AOI211_X1 g729(.A(new_n915), .B(new_n325), .C1(new_n856), .C2(new_n868), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n914), .B1(new_n916), .B2(KEYINPUT56), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n189), .A2(G952), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n856), .A2(new_n868), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n920), .A2(G210), .A3(G902), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(new_n912), .A3(new_n913), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n917), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n917), .A2(KEYINPUT120), .A3(new_n922), .A4(new_n919), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(G51));
  INV_X1    g741(.A(KEYINPUT121), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n869), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n920), .A2(KEYINPUT54), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n856), .A2(new_n868), .A3(KEYINPUT121), .A4(new_n857), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n756), .B(KEYINPUT57), .Z(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n551), .A2(new_n554), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n920), .A2(G902), .A3(new_n792), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n918), .B1(new_n936), .B2(new_n937), .ZN(G54));
  INV_X1    g752(.A(KEYINPUT58), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT122), .B1(new_n939), .B2(new_n624), .ZN(new_n940));
  OR3_X1    g754(.A1(new_n939), .A2(new_n624), .A3(KEYINPUT122), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n920), .A2(G902), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n475), .A2(new_n481), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n942), .A2(KEYINPUT123), .A3(new_n943), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT123), .B1(new_n942), .B2(new_n943), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n919), .B(new_n944), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(G60));
  XNOR2_X1  g762(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n525), .A2(new_n325), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n932), .A2(new_n630), .A3(new_n632), .A4(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n873), .A2(new_n951), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n630), .A2(new_n632), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n918), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n952), .A2(new_n955), .ZN(G63));
  NAND2_X1  g770(.A1(G217), .A2(G902), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT125), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT60), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n920), .B(new_n959), .C1(new_n655), .C2(new_n656), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n920), .A2(new_n959), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n603), .A2(new_n604), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n960), .B(new_n919), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n964));
  AOI21_X1  g778(.A(KEYINPUT61), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n963), .B(new_n965), .ZN(G66));
  NAND2_X1  g780(.A1(new_n844), .A2(new_n847), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n189), .ZN(new_n968));
  OAI21_X1  g782(.A(G953), .B1(new_n425), .B2(new_n343), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n406), .B1(G898), .B2(new_n189), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(G69));
  NAND2_X1  g786(.A1(new_n477), .A2(new_n478), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n268), .B(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n827), .ZN(new_n975));
  NAND2_X1  g789(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n697), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n697), .A2(new_n975), .ZN(new_n978));
  AND2_X1   g792(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n979));
  NOR2_X1   g793(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n820), .A2(new_n809), .A3(new_n977), .A4(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n815), .A2(new_n816), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n983), .A2(new_n695), .A3(new_n817), .A4(new_n841), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n974), .B1(new_n986), .B2(new_n189), .ZN(new_n987));
  INV_X1    g801(.A(new_n742), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n799), .A2(new_n694), .A3(new_n988), .A4(new_n895), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n820), .A2(new_n809), .A3(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n777), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n991), .A2(new_n779), .A3(new_n975), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n990), .A2(G953), .A3(new_n992), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n282), .B(new_n973), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n667), .A2(new_n189), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n997));
  OR3_X1    g811(.A1(new_n987), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n997), .B1(new_n987), .B2(new_n996), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(G72));
  NAND2_X1  g814(.A1(G472), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT63), .Z(new_n1002));
  INV_X1    g816(.A(new_n681), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1003), .B1(new_n193), .B2(new_n317), .ZN(new_n1004));
  AND4_X1   g818(.A1(new_n870), .A2(new_n871), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n982), .A2(new_n967), .A3(new_n985), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1002), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n193), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NOR3_X1   g822(.A1(new_n990), .A2(new_n967), .A3(new_n992), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n317), .B1(new_n1009), .B2(new_n1007), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  AOI211_X1 g825(.A(new_n918), .B(new_n1005), .C1(new_n1011), .C2(new_n269), .ZN(G57));
endmodule


