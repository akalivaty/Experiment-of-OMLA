//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n813, new_n814,
    new_n815, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  NAND2_X1  g001(.A1(G225gat), .A2(G233gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n203), .B(KEYINPUT82), .Z(new_n204));
  XNOR2_X1  g003(.A(G155gat), .B(G162gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT79), .ZN(new_n206));
  XNOR2_X1  g005(.A(G141gat), .B(G148gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(KEYINPUT80), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(KEYINPUT80), .ZN(new_n209));
  INV_X1    g008(.A(G155gat), .ZN(new_n210));
  INV_X1    g009(.A(G162gat), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT2), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n206), .B1(new_n208), .B2(new_n213), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n207), .A2(KEYINPUT81), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n207), .A2(KEYINPUT81), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n215), .A2(new_n216), .A3(new_n205), .A4(new_n212), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G113gat), .ZN(new_n220));
  INV_X1    g019(.A(G120gat), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT1), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(new_n220), .B2(new_n221), .ZN(new_n223));
  XOR2_X1   g022(.A(G127gat), .B(G134gat), .Z(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(KEYINPUT69), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT68), .B(G134gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G127gat), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n228), .B(new_n223), .C1(G127gat), .C2(G134gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n219), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT83), .B(KEYINPUT4), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n204), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n226), .A2(new_n229), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(new_n218), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT4), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n218), .A2(KEYINPUT3), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n218), .A2(KEYINPUT3), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n237), .A3(new_n233), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n232), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n233), .A2(new_n218), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n230), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n204), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n239), .A2(KEYINPUT5), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G1gat), .B(G29gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT0), .ZN(new_n245));
  XNOR2_X1  g044(.A(G57gat), .B(G85gat), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n245), .B(new_n246), .Z(new_n247));
  OR2_X1    g046(.A1(new_n234), .A2(KEYINPUT4), .ZN(new_n248));
  OR2_X1    g047(.A1(new_n230), .A2(new_n231), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n204), .A2(KEYINPUT5), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n238), .A4(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n243), .A2(new_n247), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT84), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n243), .A2(new_n251), .ZN(new_n254));
  INV_X1    g053(.A(new_n247), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT6), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT84), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n243), .A2(new_n258), .A3(new_n247), .A4(new_n251), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n253), .A2(new_n256), .A3(new_n257), .A4(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n254), .A2(KEYINPUT6), .A3(new_n255), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G197gat), .B(G204gat), .ZN(new_n263));
  INV_X1    g062(.A(G211gat), .ZN(new_n264));
  INV_X1    g063(.A(G218gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n263), .B1(KEYINPUT22), .B2(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(G211gat), .B(G218gat), .Z(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G226gat), .A2(G233gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT24), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n274), .B1(G183gat), .B2(G190gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT66), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT23), .ZN(new_n279));
  INV_X1    g078(.A(G169gat), .ZN(new_n280));
  INV_X1    g079(.A(G176gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT23), .ZN(new_n283));
  INV_X1    g082(.A(new_n276), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AND4_X1   g084(.A1(KEYINPUT25), .A2(new_n275), .A3(new_n279), .A4(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n276), .A2(KEYINPUT23), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT65), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n290), .B1(G183gat), .B2(G190gat), .ZN(new_n291));
  OR3_X1    g090(.A1(new_n290), .A2(G183gat), .A3(G190gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n287), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  OR2_X1    g093(.A1(new_n286), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT27), .B(G183gat), .ZN(new_n296));
  INV_X1    g095(.A(G190gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT67), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(KEYINPUT28), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT26), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n278), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n282), .B1(KEYINPUT26), .B2(new_n284), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n302), .A2(new_n303), .B1(G183gat), .B2(G190gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n295), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT29), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n272), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n271), .B1(new_n295), .B2(new_n305), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n270), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n306), .A2(new_n272), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT29), .B1(new_n295), .B2(new_n305), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n311), .B(new_n269), .C1(new_n272), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G8gat), .B(G36gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(G64gat), .B(G92gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(KEYINPUT30), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n310), .A2(new_n313), .A3(KEYINPUT30), .A4(new_n317), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n314), .A2(new_n318), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n324), .A2(new_n322), .A3(new_n321), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n320), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n262), .A2(new_n326), .A3(KEYINPUT87), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n226), .A2(new_n229), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n300), .A2(new_n304), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n286), .A2(new_n294), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n295), .A2(new_n233), .A3(new_n305), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n331), .A2(new_n332), .A3(G227gat), .A4(G233gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT33), .ZN(new_n334));
  XNOR2_X1  g133(.A(G15gat), .B(G43gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT71), .ZN(new_n336));
  XNOR2_X1  g135(.A(G71gat), .B(G99gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n333), .B(KEYINPUT32), .C1(new_n334), .C2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n338), .B1(new_n333), .B2(KEYINPUT32), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n333), .A2(KEYINPUT70), .A3(new_n334), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT70), .B1(new_n333), .B2(new_n334), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n339), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n331), .A2(new_n332), .B1(G227gat), .B2(G233gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT73), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT34), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n347), .B(KEYINPUT74), .Z(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n346), .A2(KEYINPUT34), .ZN(new_n350));
  OR3_X1    g149(.A1(new_n345), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n349), .B1(new_n345), .B2(new_n350), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n344), .A2(new_n353), .A3(KEYINPUT76), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT76), .B1(new_n344), .B2(new_n353), .ZN(new_n355));
  OR2_X1    g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT3), .B1(new_n269), .B2(new_n307), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n219), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n236), .A2(new_n307), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(new_n270), .ZN(new_n360));
  XNOR2_X1  g159(.A(G78gat), .B(G106gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  NAND2_X1  g161(.A1(G228gat), .A2(G233gat), .ZN(new_n363));
  INV_X1    g162(.A(G22gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT31), .B(G50gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n362), .B(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT75), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(new_n344), .B2(new_n353), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n351), .A2(new_n352), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n333), .A2(new_n334), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT70), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(new_n341), .A3(new_n340), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n371), .A2(new_n375), .A3(KEYINPUT75), .A4(new_n339), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n370), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n327), .A2(new_n356), .A3(new_n368), .A4(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT87), .B1(new_n262), .B2(new_n326), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n202), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT86), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT37), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n310), .A2(new_n382), .A3(new_n313), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n382), .B1(new_n310), .B2(new_n313), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n383), .A2(new_n384), .A3(new_n317), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT38), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n381), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n319), .B1(new_n385), .B2(new_n386), .ZN(new_n388));
  OR2_X1    g187(.A1(new_n384), .A2(new_n317), .ZN(new_n389));
  OAI211_X1 g188(.A(KEYINPUT86), .B(KEYINPUT38), .C1(new_n389), .C2(new_n383), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n248), .A2(new_n249), .A3(new_n238), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT39), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n393), .A3(new_n204), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n247), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT40), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT39), .B1(new_n241), .B2(new_n204), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n397), .B1(new_n392), .B2(new_n204), .ZN(new_n398));
  OR3_X1    g197(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n396), .B1(new_n395), .B2(new_n398), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n256), .A3(new_n400), .ZN(new_n401));
  OAI22_X1  g200(.A1(new_n391), .A2(new_n262), .B1(new_n326), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT36), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n356), .A2(new_n403), .A3(new_n377), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n351), .A2(KEYINPUT72), .A3(new_n352), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n405), .A2(new_n344), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n344), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT36), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n402), .A2(new_n404), .A3(new_n368), .A4(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n368), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n370), .B(new_n376), .C1(new_n354), .C2(new_n355), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n410), .B(new_n408), .C1(new_n411), .C2(KEYINPUT36), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n410), .A2(new_n406), .A3(new_n407), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT35), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n256), .B(KEYINPUT85), .Z(new_n416));
  NAND3_X1  g215(.A1(new_n253), .A2(new_n257), .A3(new_n259), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n261), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n325), .A2(new_n323), .ZN(new_n419));
  OR2_X1    g218(.A1(new_n419), .A2(KEYINPUT78), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n320), .B1(new_n419), .B2(KEYINPUT78), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n380), .B(new_n409), .C1(new_n415), .C2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT17), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT90), .ZN(new_n425));
  INV_X1    g224(.A(G43gat), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n425), .B1(new_n426), .B2(G50gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(G50gat), .ZN(new_n428));
  INV_X1    g227(.A(G50gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n429), .A2(KEYINPUT90), .A3(G43gat), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n427), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT15), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AND3_X1   g232(.A1(KEYINPUT89), .A2(G29gat), .A3(G36gat), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT89), .B1(G29gat), .B2(G36gat), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT14), .ZN(new_n437));
  INV_X1    g236(.A(G29gat), .ZN(new_n438));
  INV_X1    g237(.A(G36gat), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n429), .A2(G43gat), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(new_n428), .A3(KEYINPUT15), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n436), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n433), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT88), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n440), .A2(new_n447), .ZN(new_n448));
  NOR3_X1   g247(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT88), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n450), .A3(new_n441), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n444), .B1(new_n451), .B2(new_n436), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n424), .B1(new_n446), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT91), .ZN(new_n454));
  XNOR2_X1  g253(.A(G15gat), .B(G22gat), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n454), .B1(new_n455), .B2(G1gat), .ZN(new_n456));
  INV_X1    g255(.A(G1gat), .ZN(new_n457));
  INV_X1    g256(.A(G15gat), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n458), .A2(G22gat), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n364), .A2(G15gat), .ZN(new_n460));
  OAI211_X1 g259(.A(KEYINPUT91), .B(new_n457), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n457), .A2(KEYINPUT16), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n455), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n456), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n465));
  INV_X1    g264(.A(G8gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n364), .A2(G15gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n458), .A2(G22gat), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT92), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n467), .A2(new_n468), .A3(new_n462), .A4(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n465), .A2(new_n466), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n463), .A2(KEYINPUT92), .ZN(new_n472));
  AOI22_X1  g271(.A1(G8gat), .A2(new_n464), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n441), .B1(new_n449), .B2(KEYINPUT88), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n440), .A2(new_n447), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n436), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n444), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n431), .A2(new_n432), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n479), .A2(new_n444), .A3(new_n436), .A4(new_n442), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n480), .A3(KEYINPUT17), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n453), .A2(new_n473), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n464), .A2(G8gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n471), .A2(new_n472), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n478), .A2(new_n480), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G229gat), .A2(G233gat), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n482), .A2(KEYINPUT18), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n488), .B(KEYINPUT13), .Z(new_n490));
  NOR2_X1   g289(.A1(new_n485), .A2(new_n486), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n483), .A2(new_n484), .B1(new_n478), .B2(new_n480), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G113gat), .B(G141gat), .ZN(new_n495));
  INV_X1    g294(.A(G197gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT11), .B(G169gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  XOR2_X1   g298(.A(new_n499), .B(KEYINPUT12), .Z(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n482), .A2(new_n487), .A3(new_n488), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT18), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n494), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT93), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n502), .A2(KEYINPUT93), .A3(new_n503), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n494), .A3(new_n508), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n509), .A2(KEYINPUT94), .A3(new_n500), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT94), .B1(new_n509), .B2(new_n500), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G71gat), .A2(G78gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(KEYINPUT95), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT96), .B1(G71gat), .B2(G78gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(G71gat), .A2(G78gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT96), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n514), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT97), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n514), .A2(KEYINPUT97), .A3(new_n515), .A4(new_n518), .ZN(new_n522));
  INV_X1    g321(.A(G57gat), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n523), .A2(G64gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(G64gat), .ZN(new_n525));
  INV_X1    g324(.A(new_n513), .ZN(new_n526));
  OAI22_X1  g325(.A1(new_n524), .A2(new_n525), .B1(new_n526), .B2(KEYINPUT9), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n521), .A2(new_n522), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n523), .A2(KEYINPUT98), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT98), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(G57gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(new_n531), .A3(G64gat), .ZN(new_n532));
  INV_X1    g331(.A(new_n525), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n532), .A2(KEYINPUT99), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT99), .B1(new_n532), .B2(new_n533), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT100), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n526), .B1(KEYINPUT9), .B2(new_n516), .ZN(new_n537));
  NOR4_X1   g336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n532), .A2(new_n533), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT99), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT98), .B(G57gat), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n525), .B1(new_n542), .B2(G64gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT99), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT100), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n528), .B1(new_n538), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT21), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G231gat), .A2(G233gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(G127gat), .ZN(new_n551));
  XOR2_X1   g350(.A(G183gat), .B(G211gat), .Z(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n473), .B1(new_n546), .B2(new_n547), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(KEYINPUT101), .Z(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(new_n210), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n555), .B(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n552), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n551), .B(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n558), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G85gat), .A2(G92gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT7), .ZN(new_n566));
  INV_X1    g365(.A(G85gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT103), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT103), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(G85gat), .ZN(new_n570));
  INV_X1    g369(.A(G92gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G99gat), .A2(G106gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT8), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n572), .A2(KEYINPUT104), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT104), .B1(new_n572), .B2(new_n574), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n566), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G99gat), .B(G106gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n578), .B(new_n566), .C1(new_n575), .C2(new_n576), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(new_n481), .A3(new_n453), .ZN(new_n583));
  NAND3_X1  g382(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n486), .A3(new_n581), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT105), .ZN(new_n587));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n583), .A2(new_n590), .A3(new_n584), .A4(new_n585), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n592), .B(KEYINPUT102), .Z(new_n593));
  XNOR2_X1  g392(.A(G134gat), .B(G162gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  NAND3_X1  g394(.A1(new_n589), .A2(new_n591), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n587), .B1(new_n586), .B2(new_n588), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT106), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n597), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT106), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n591), .A2(new_n595), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n599), .A2(new_n600), .A3(new_n589), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n604), .A2(new_n591), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n605), .A2(new_n595), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G120gat), .B(G148gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(G176gat), .B(G204gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  NAND2_X1  g409(.A1(new_n546), .A2(new_n582), .ZN(new_n611));
  INV_X1    g410(.A(new_n537), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n612), .B1(new_n543), .B2(KEYINPUT99), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n536), .B1(new_n613), .B2(new_n534), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n541), .A2(KEYINPUT100), .A3(new_n544), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n616), .A2(new_n581), .A3(new_n580), .A4(new_n528), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G230gat), .A2(G233gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT108), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT10), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n611), .A2(new_n617), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n582), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n626), .A2(KEYINPUT10), .A3(new_n616), .A4(new_n528), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n619), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n610), .B1(new_n623), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT107), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n620), .B1(new_n625), .B2(new_n627), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT107), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n623), .A2(new_n633), .A3(new_n610), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n564), .A2(new_n607), .A3(new_n637), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n423), .A2(new_n512), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n418), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G1gat), .ZN(G1324gat));
  INV_X1    g441(.A(new_n326), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT16), .B(G8gat), .Z(new_n644));
  NAND3_X1  g443(.A1(new_n639), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n639), .A2(new_n643), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n645), .B1(new_n647), .B2(new_n466), .ZN(new_n648));
  MUX2_X1   g447(.A(new_n645), .B(new_n648), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g448(.A(new_n411), .ZN(new_n650));
  AOI21_X1  g449(.A(G15gat), .B1(new_n639), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT109), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n404), .A2(new_n408), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n458), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n652), .B1(new_n639), .B2(new_n655), .ZN(G1326gat));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n410), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT43), .B(G22gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1327gat));
  NAND2_X1  g458(.A1(new_n380), .A2(new_n409), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n422), .B1(new_n412), .B2(new_n414), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n607), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n564), .ZN(new_n664));
  INV_X1    g463(.A(new_n512), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n664), .A2(new_n665), .A3(new_n637), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n663), .A2(new_n438), .A3(new_n640), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT45), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n662), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n423), .A2(KEYINPUT44), .A3(new_n607), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND3_X1   g471(.A1(new_n672), .A2(new_n640), .A3(new_n666), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n668), .B1(new_n438), .B2(new_n673), .ZN(G1328gat));
  NAND4_X1  g473(.A1(new_n663), .A2(new_n439), .A3(new_n643), .A4(new_n666), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT46), .Z(new_n676));
  NAND4_X1  g475(.A1(new_n670), .A2(new_n671), .A3(new_n643), .A4(new_n666), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT110), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(G36gat), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n676), .B1(new_n679), .B2(new_n681), .ZN(G1329gat));
  NAND4_X1  g481(.A1(new_n670), .A2(new_n671), .A3(new_n653), .A4(new_n666), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(G43gat), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n663), .A2(new_n426), .A3(new_n650), .A4(new_n666), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT47), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1330gat));
  NAND4_X1  g487(.A1(new_n670), .A2(new_n671), .A3(new_n410), .A4(new_n666), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(G50gat), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n663), .A2(new_n429), .A3(new_n410), .A4(new_n666), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT111), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT48), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT48), .ZN(new_n695));
  AOI211_X1 g494(.A(KEYINPUT111), .B(new_n695), .C1(new_n690), .C2(new_n691), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n694), .A2(new_n696), .ZN(G1331gat));
  NOR2_X1   g496(.A1(new_n564), .A2(new_n607), .ZN(new_n698));
  AND4_X1   g497(.A1(new_n423), .A2(new_n665), .A3(new_n698), .A4(new_n637), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n640), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n700), .B(new_n542), .Z(G1332gat));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n643), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT49), .B(G64gat), .Z(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n702), .B2(new_n704), .ZN(G1333gat));
  INV_X1    g504(.A(G71gat), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n699), .A2(new_n706), .A3(new_n650), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n699), .A2(new_n653), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(new_n709), .B2(new_n706), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT50), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1334gat));
  NAND2_X1  g511(.A1(new_n699), .A2(new_n410), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g513(.A1(new_n664), .A2(new_n512), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n607), .B(new_n715), .C1(new_n660), .C2(new_n661), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT51), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT113), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n423), .A2(KEYINPUT51), .A3(new_n607), .A4(new_n715), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n716), .A2(KEYINPUT113), .A3(new_n717), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n568), .A2(new_n570), .ZN(new_n723));
  INV_X1    g522(.A(new_n637), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n418), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n721), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n664), .A2(new_n512), .A3(new_n724), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n670), .A2(new_n671), .A3(new_n640), .A4(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n723), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n728), .A2(new_n729), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n726), .B1(new_n731), .B2(new_n732), .ZN(G1336gat));
  NAND4_X1  g532(.A1(new_n670), .A2(new_n671), .A3(new_n643), .A4(new_n727), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G92gat), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n724), .A2(new_n326), .A3(G92gat), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n721), .A2(new_n722), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n718), .A2(new_n720), .ZN(new_n740));
  AOI22_X1  g539(.A1(G92gat), .A2(new_n734), .B1(new_n740), .B2(new_n738), .ZN(new_n741));
  OAI22_X1  g540(.A1(new_n737), .A2(new_n739), .B1(new_n741), .B2(new_n736), .ZN(G1337gat));
  NAND3_X1  g541(.A1(new_n672), .A2(new_n653), .A3(new_n727), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G99gat), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n411), .A2(G99gat), .A3(new_n724), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT114), .Z(new_n746));
  NAND3_X1  g545(.A1(new_n721), .A2(new_n722), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n747), .ZN(G1338gat));
  NAND4_X1  g547(.A1(new_n670), .A2(new_n671), .A3(new_n410), .A4(new_n727), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT53), .B1(new_n749), .B2(G106gat), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n724), .A2(G106gat), .A3(new_n368), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n721), .A2(new_n722), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n749), .A2(G106gat), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n755), .B1(new_n740), .B2(new_n751), .ZN(new_n756));
  INV_X1    g555(.A(new_n751), .ZN(new_n757));
  AOI211_X1 g556(.A(KEYINPUT115), .B(new_n757), .C1(new_n718), .C2(new_n720), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n754), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n753), .B1(new_n759), .B2(new_n760), .ZN(G1339gat));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n634), .A2(KEYINPUT107), .ZN(new_n763));
  AOI211_X1 g562(.A(new_n632), .B(new_n620), .C1(new_n625), .C2(new_n627), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n625), .A2(new_n627), .A3(new_n620), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT54), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT54), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n610), .B1(new_n634), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n762), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n765), .A2(KEYINPUT54), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n633), .A2(new_n772), .A3(new_n635), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n773), .A2(new_n769), .A3(KEYINPUT55), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n771), .A2(new_n512), .A3(new_n636), .A4(new_n774), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n491), .A2(new_n492), .A3(new_n490), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n488), .B1(new_n482), .B2(new_n487), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n499), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AND4_X1   g577(.A1(new_n623), .A2(new_n610), .A3(new_n633), .A4(new_n635), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n505), .B(new_n778), .C1(new_n779), .C2(new_n630), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n607), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n505), .A2(new_n778), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n784), .B1(new_n603), .B2(new_n606), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n785), .A2(new_n636), .A3(new_n771), .A4(new_n774), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n783), .A2(KEYINPUT116), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n607), .B1(new_n775), .B2(new_n780), .ZN(new_n789));
  INV_X1    g588(.A(new_n786), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n787), .A2(new_n564), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n638), .A2(new_n665), .ZN(new_n793));
  AOI211_X1 g592(.A(new_n410), .B(new_n411), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n418), .A2(new_n643), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT117), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n794), .A2(KEYINPUT117), .A3(new_n795), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n798), .A2(G113gat), .A3(new_n512), .A4(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n418), .B1(new_n792), .B2(new_n793), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(new_n413), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n326), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n220), .B1(new_n803), .B2(new_n665), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n805), .B(new_n806), .ZN(G1340gat));
  INV_X1    g606(.A(new_n803), .ZN(new_n808));
  AOI21_X1  g607(.A(G120gat), .B1(new_n808), .B2(new_n637), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n798), .A2(new_n799), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n724), .A2(new_n221), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(G1341gat));
  INV_X1    g611(.A(G127gat), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n808), .A2(new_n813), .A3(new_n664), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n810), .A2(new_n664), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(new_n813), .ZN(G1342gat));
  NAND2_X1  g615(.A1(new_n810), .A2(new_n607), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(G134gat), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n643), .A2(new_n227), .A3(new_n782), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g619(.A(new_n820), .B(KEYINPUT56), .Z(new_n821));
  NAND2_X1  g620(.A1(new_n818), .A2(new_n821), .ZN(G1343gat));
  INV_X1    g621(.A(G141gat), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n654), .A2(new_n795), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n783), .A2(new_n786), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n564), .A2(new_n825), .B1(new_n638), .B2(new_n665), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n826), .A2(new_n827), .A3(new_n368), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n791), .A2(new_n564), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n789), .A2(new_n790), .A3(new_n788), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n793), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT57), .B1(new_n831), .B2(new_n410), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n828), .B1(new_n832), .B2(KEYINPUT119), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n368), .B1(new_n792), .B2(new_n793), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n834), .B1(new_n835), .B2(KEYINPUT57), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n824), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n823), .B1(new_n837), .B2(new_n512), .ZN(new_n838));
  AOI211_X1 g637(.A(new_n418), .B(new_n412), .C1(new_n792), .C2(new_n793), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n839), .A2(new_n326), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n512), .A2(new_n823), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT120), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT58), .B1(new_n838), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n832), .A2(KEYINPUT119), .ZN(new_n846));
  INV_X1    g645(.A(new_n828), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n836), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n824), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n512), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(G141gat), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n852), .A3(new_n843), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n845), .A2(new_n853), .ZN(G1344gat));
  INV_X1    g653(.A(G148gat), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n855), .A3(new_n637), .ZN(new_n856));
  AOI211_X1 g655(.A(KEYINPUT59), .B(new_n855), .C1(new_n837), .C2(new_n637), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n835), .A2(KEYINPUT57), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n827), .B1(new_n826), .B2(new_n368), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n724), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n849), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n858), .B1(new_n862), .B2(G148gat), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n856), .B1(new_n857), .B2(new_n863), .ZN(G1345gat));
  AOI21_X1  g663(.A(G155gat), .B1(new_n840), .B2(new_n664), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n564), .A2(new_n210), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT121), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n865), .B1(new_n837), .B2(new_n867), .ZN(G1346gat));
  NAND4_X1  g667(.A1(new_n839), .A2(new_n211), .A3(new_n326), .A4(new_n607), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n837), .A2(new_n607), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(new_n211), .ZN(G1347gat));
  AOI21_X1  g670(.A(new_n640), .B1(new_n792), .B2(new_n793), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n872), .A2(new_n413), .A3(new_n643), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n280), .A3(new_n512), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n640), .A2(new_n326), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n794), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(G169gat), .B1(new_n876), .B2(new_n665), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n877), .A2(KEYINPUT122), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(KEYINPUT122), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n874), .B1(new_n878), .B2(new_n879), .ZN(G1348gat));
  OAI21_X1  g679(.A(G176gat), .B1(new_n876), .B2(new_n724), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n873), .A2(new_n281), .A3(new_n637), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1349gat));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(KEYINPUT60), .ZN(new_n885));
  OAI21_X1  g684(.A(G183gat), .B1(new_n876), .B2(new_n564), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n873), .A2(new_n296), .A3(new_n664), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n884), .A2(KEYINPUT60), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n888), .B(new_n889), .ZN(G1350gat));
  NAND3_X1  g689(.A1(new_n794), .A2(new_n607), .A3(new_n875), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n297), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n873), .A2(new_n297), .A3(new_n607), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G1351gat));
  NOR2_X1   g697(.A1(new_n412), .A2(new_n326), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT125), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n900), .A2(new_n872), .ZN(new_n901));
  AOI21_X1  g700(.A(G197gat), .B1(new_n901), .B2(new_n512), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n654), .A2(new_n875), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n903), .B1(new_n859), .B2(new_n860), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n665), .A2(new_n496), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(G1352gat));
  INV_X1    g705(.A(G204gat), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n901), .A2(new_n907), .A3(new_n637), .ZN(new_n908));
  XOR2_X1   g707(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n909));
  XNOR2_X1  g708(.A(new_n908), .B(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n903), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n861), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n910), .B1(new_n907), .B2(new_n912), .ZN(G1353gat));
  NAND3_X1  g712(.A1(new_n901), .A2(new_n264), .A3(new_n664), .ZN(new_n914));
  AOI211_X1 g713(.A(new_n827), .B(new_n368), .C1(new_n792), .C2(new_n793), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n825), .A2(new_n564), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n793), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT57), .B1(new_n917), .B2(new_n410), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n664), .B(new_n911), .C1(new_n915), .C2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT127), .ZN(new_n920));
  OAI21_X1  g719(.A(G211gat), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT127), .B1(new_n904), .B2(new_n664), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT63), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT63), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n921), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n914), .B1(new_n925), .B2(new_n927), .ZN(G1354gat));
  NAND3_X1  g727(.A1(new_n901), .A2(new_n265), .A3(new_n607), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n904), .A2(new_n607), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n930), .B2(new_n265), .ZN(G1355gat));
endmodule


