//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT66), .ZN(new_n213));
  XOR2_X1   g0013(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n208), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n215), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n213), .A2(new_n214), .ZN(new_n222));
  XOR2_X1   g0022(.A(KEYINPUT67), .B(G244), .Z(new_n223));
  AND2_X1   g0023(.A1(new_n223), .A2(G77), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G87), .A2(G250), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n210), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n221), .A2(new_n222), .A3(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G226), .B(G232), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(KEYINPUT69), .B(KEYINPUT70), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G68), .Z(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G169), .ZN(new_n251));
  INV_X1    g0051(.A(G238), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT74), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n252), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(new_n257), .B2(new_n256), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G232), .A3(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(G226), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G97), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n268), .B(new_n270), .C1(new_n265), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n253), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n259), .A2(new_n262), .A3(new_n273), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n274), .A2(KEYINPUT13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(KEYINPUT13), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n251), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT14), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n275), .A2(G179), .A3(new_n276), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(new_n277), .B2(new_n278), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT76), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  OR2_X1    g0083(.A1(new_n277), .A2(new_n278), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT76), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n284), .A2(new_n285), .A3(new_n279), .A4(new_n281), .ZN(new_n286));
  INV_X1    g0086(.A(G13), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n287), .A2(new_n208), .A3(G1), .ZN(new_n288));
  INV_X1    g0088(.A(G68), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT12), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n216), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(G1), .B2(new_n208), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n265), .A2(G20), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G77), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n297), .A2(new_n298), .B1(new_n208), .B2(G68), .ZN(new_n299));
  NOR2_X1   g0099(.A1(G20), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(new_n202), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n293), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT11), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n291), .B1(new_n289), .B2(new_n295), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n304), .B2(new_n303), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT75), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT77), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n283), .A2(new_n286), .A3(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n256), .A2(G226), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n267), .A2(G222), .A3(new_n269), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n267), .A2(G1698), .ZN(new_n312));
  INV_X1    g0112(.A(G223), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n311), .B1(new_n298), .B2(new_n267), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  AOI211_X1 g0114(.A(new_n261), .B(new_n310), .C1(new_n314), .C2(new_n253), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G190), .ZN(new_n316));
  NOR2_X1   g0116(.A1(KEYINPUT8), .A2(G58), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT71), .B(G58), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(KEYINPUT8), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n296), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n300), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n293), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n288), .A2(new_n202), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n323), .B(new_n324), .C1(new_n202), .C2(new_n295), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT9), .ZN(new_n326));
  OR2_X1    g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n326), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n316), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT73), .ZN(new_n330));
  AOI21_X1  g0130(.A(KEYINPUT10), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G200), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n329), .B1(new_n332), .B2(new_n315), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  OAI221_X1 g0134(.A(new_n329), .B1(new_n330), .B2(KEYINPUT10), .C1(new_n332), .C2(new_n315), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n315), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n325), .B1(new_n315), .B2(G169), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n275), .A2(new_n276), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G200), .ZN(new_n343));
  INV_X1    g0143(.A(G190), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n343), .B(new_n307), .C1(new_n344), .C2(new_n342), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n288), .A2(new_n298), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n295), .B2(new_n298), .ZN(new_n347));
  XOR2_X1   g0147(.A(KEYINPUT8), .B(G58), .Z(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(new_n300), .B1(G20), .B2(G77), .ZN(new_n349));
  XOR2_X1   g0149(.A(KEYINPUT15), .B(G87), .Z(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT72), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n349), .B1(new_n351), .B2(new_n297), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n347), .B1(new_n352), .B2(new_n293), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n267), .A2(G232), .A3(new_n269), .ZN(new_n354));
  INV_X1    g0154(.A(G107), .ZN(new_n355));
  OAI221_X1 g0155(.A(new_n354), .B1(new_n355), .B2(new_n267), .C1(new_n312), .C2(new_n252), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n253), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n261), .B1(new_n256), .B2(new_n223), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n353), .B1(new_n251), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(new_n337), .A3(new_n358), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n359), .A2(G200), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(new_n353), .C1(new_n344), .C2(new_n359), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  AND4_X1   g0165(.A1(new_n309), .A2(new_n341), .A3(new_n345), .A4(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G58), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT71), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT71), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G58), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n370), .A3(G68), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n208), .B1(new_n371), .B2(new_n219), .ZN(new_n372));
  INV_X1    g0172(.A(G159), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n301), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT80), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT80), .ZN(new_n376));
  INV_X1    g0176(.A(new_n374), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n201), .B1(new_n318), .B2(G68), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n376), .B(new_n377), .C1(new_n378), .C2(new_n208), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n264), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n265), .A2(KEYINPUT78), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT78), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G33), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n382), .B1(new_n386), .B2(KEYINPUT3), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT7), .B1(new_n387), .B2(G20), .ZN(new_n388));
  XNOR2_X1  g0188(.A(KEYINPUT78), .B(G33), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n264), .B1(new_n389), .B2(new_n263), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n391), .A3(new_n208), .ZN(new_n392));
  AND4_X1   g0192(.A1(KEYINPUT79), .A2(new_n388), .A3(G68), .A4(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n263), .B1(new_n383), .B2(new_n385), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n208), .B1(new_n394), .B2(new_n382), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n289), .B1(new_n395), .B2(KEYINPUT7), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT79), .B1(new_n396), .B2(new_n392), .ZN(new_n397));
  OAI211_X1 g0197(.A(KEYINPUT16), .B(new_n381), .C1(new_n393), .C2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  OR3_X1    g0199(.A1(new_n263), .A2(KEYINPUT81), .A3(G33), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n266), .A2(KEYINPUT81), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n400), .B(new_n401), .C1(new_n386), .C2(KEYINPUT3), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n391), .A2(G20), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n391), .B1(new_n267), .B2(G20), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n289), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n399), .B1(new_n380), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT82), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI211_X1 g0209(.A(KEYINPUT82), .B(new_n399), .C1(new_n380), .C2(new_n406), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n398), .A2(new_n409), .A3(new_n293), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT83), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n410), .A2(new_n293), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT83), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(new_n398), .A4(new_n409), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n319), .A2(new_n288), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n319), .B2(new_n295), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n261), .B1(new_n256), .B2(G232), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G87), .ZN(new_n422));
  XOR2_X1   g0222(.A(new_n422), .B(KEYINPUT84), .Z(new_n423));
  MUX2_X1   g0223(.A(G223), .B(G226), .S(G1698), .Z(new_n424));
  AOI21_X1  g0224(.A(new_n423), .B1(new_n387), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n421), .B1(new_n254), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(new_n337), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(G169), .B2(new_n426), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT18), .B1(new_n420), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n418), .B1(new_n412), .B2(new_n415), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT18), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n431), .A2(new_n432), .A3(new_n428), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT17), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n426), .A2(G200), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n344), .B2(new_n426), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  AND4_X1   g0237(.A1(new_n434), .A2(new_n416), .A3(new_n419), .A4(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n434), .B1(new_n431), .B2(new_n437), .ZN(new_n439));
  OAI22_X1  g0239(.A1(new_n430), .A2(new_n433), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n366), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n267), .A2(KEYINPUT4), .A3(G244), .A4(new_n269), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n267), .A2(G250), .A3(G1698), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G283), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n387), .A2(G244), .A3(new_n269), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n443), .B(new_n446), .C1(new_n447), .C2(KEYINPUT4), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n253), .ZN(new_n449));
  INV_X1    g0249(.A(G45), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n450), .A2(G1), .ZN(new_n451));
  INV_X1    g0251(.A(G41), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(KEYINPUT5), .B2(new_n452), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n452), .A2(KEYINPUT5), .ZN(new_n454));
  OR3_X1    g0254(.A1(new_n453), .A2(new_n260), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n254), .B1(new_n453), .B2(new_n454), .ZN(new_n456));
  INV_X1    g0256(.A(G257), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n449), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT86), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n332), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n460), .B2(new_n459), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n355), .B1(new_n404), .B2(new_n405), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT6), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n271), .A2(new_n355), .ZN(new_n465));
  NOR2_X1   g0265(.A1(G97), .A2(G107), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n355), .A2(KEYINPUT6), .A3(G97), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI22_X1  g0269(.A1(new_n469), .A2(new_n208), .B1(new_n298), .B2(new_n301), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n293), .B1(new_n463), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n288), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT85), .B1(new_n265), .B2(G1), .ZN(new_n473));
  OR3_X1    g0273(.A1(new_n265), .A2(KEYINPUT85), .A3(G1), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(new_n293), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G97), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n471), .B(new_n477), .C1(G97), .C2(new_n472), .ZN(new_n478));
  INV_X1    g0278(.A(new_n459), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(G190), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n462), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT87), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n462), .A2(KEYINPUT87), .A3(new_n480), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n479), .A2(new_n337), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n459), .A2(new_n251), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(new_n478), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n267), .A2(new_n208), .A3(G87), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT22), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT23), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n208), .B2(G107), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n355), .A2(KEYINPUT23), .A3(G20), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n489), .A2(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G87), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n387), .A2(new_n496), .B1(G116), .B2(new_n389), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n494), .B1(new_n497), .B2(G20), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT24), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n294), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n499), .B2(new_n498), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT25), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n472), .B2(G107), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n288), .A2(KEYINPUT25), .A3(new_n355), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n476), .A2(G107), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(G250), .A2(G1698), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n508), .B1(new_n457), .B2(G1698), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n387), .A2(new_n509), .B1(G294), .B2(new_n389), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(new_n254), .ZN(new_n511));
  INV_X1    g0311(.A(G264), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n455), .B1(new_n456), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G200), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n507), .B(new_n516), .C1(new_n344), .C2(new_n515), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n351), .A2(new_n288), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n387), .A2(new_n208), .A3(G68), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n297), .A2(new_n271), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(KEYINPUT19), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n208), .A2(new_n522), .B1(new_n466), .B2(new_n495), .ZN(new_n523));
  XOR2_X1   g0323(.A(new_n523), .B(KEYINPUT88), .Z(new_n524));
  OAI21_X1  g0324(.A(new_n293), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  XOR2_X1   g0325(.A(new_n351), .B(KEYINPUT89), .Z(new_n526));
  INV_X1    g0326(.A(new_n476), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n518), .B(new_n525), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n387), .A2(G244), .A3(G1698), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n387), .A2(G238), .A3(new_n269), .ZN(new_n530));
  INV_X1    g0330(.A(G116), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n529), .B(new_n530), .C1(new_n531), .C2(new_n386), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n253), .ZN(new_n533));
  INV_X1    g0333(.A(G250), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n253), .A2(new_n534), .A3(new_n451), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(G274), .B2(new_n451), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n251), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n533), .A2(new_n337), .A3(new_n536), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n528), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n525), .A2(new_n518), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(G87), .B2(new_n476), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n537), .A2(G200), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n542), .B(new_n543), .C1(new_n344), .C2(new_n537), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n517), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n485), .A2(new_n488), .A3(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n445), .B(new_n208), .C1(G33), .C2(new_n271), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT90), .ZN(new_n548));
  XNOR2_X1  g0348(.A(new_n547), .B(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n549), .B(new_n293), .C1(new_n208), .C2(G116), .ZN(new_n550));
  XNOR2_X1  g0350(.A(new_n550), .B(KEYINPUT20), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n288), .A2(new_n531), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n527), .B2(new_n531), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(G270), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n455), .B1(new_n456), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(G257), .A2(G1698), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n512), .B2(G1698), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n387), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(G303), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(new_n560), .B2(new_n267), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n556), .B1(new_n253), .B2(new_n561), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n554), .A2(new_n251), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT21), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT91), .ZN(new_n565));
  OR2_X1    g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n562), .A2(G179), .ZN(new_n567));
  OR2_X1    g0367(.A1(new_n554), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n563), .A2(new_n565), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n562), .A2(G190), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n554), .B(new_n570), .C1(new_n332), .C2(new_n562), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n566), .A2(new_n568), .A3(new_n569), .A4(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n514), .A2(G169), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n337), .B2(new_n514), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n506), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NOR4_X1   g0376(.A1(new_n442), .A2(new_n546), .A3(new_n572), .A4(new_n576), .ZN(G372));
  INV_X1    g0377(.A(new_n442), .ZN(new_n578));
  INV_X1    g0378(.A(new_n540), .ZN(new_n579));
  INV_X1    g0379(.A(new_n488), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n580), .A2(KEYINPUT26), .A3(new_n540), .A4(new_n544), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT26), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n544), .A2(new_n540), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n582), .B1(new_n583), .B2(new_n488), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n579), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n586), .A2(new_n576), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n585), .B1(new_n546), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n578), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n430), .A2(new_n433), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n345), .A2(new_n361), .A3(new_n360), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n309), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n438), .A2(new_n439), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n591), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n336), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n340), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n589), .A2(new_n597), .ZN(G369));
  NOR2_X1   g0398(.A1(new_n287), .A2(G20), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n207), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n600), .A2(KEYINPUT27), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(KEYINPUT27), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(G213), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(G343), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n575), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n605), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n517), .B1(new_n507), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n606), .B1(new_n608), .B2(new_n575), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(new_n586), .A3(new_n607), .ZN(new_n610));
  INV_X1    g0410(.A(new_n606), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n554), .A2(new_n607), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n586), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n572), .B2(new_n614), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n616), .A2(G330), .A3(new_n609), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(new_n617), .ZN(G399));
  INV_X1    g0418(.A(new_n211), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(G41), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G1), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n466), .A2(new_n495), .A3(new_n531), .ZN(new_n623));
  OAI22_X1  g0423(.A1(new_n622), .A2(new_n623), .B1(new_n220), .B2(new_n621), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n624), .B(KEYINPUT28), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT92), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n626), .A2(KEYINPUT29), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n588), .B2(new_n607), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n588), .A2(new_n607), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n626), .A2(KEYINPUT29), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n629), .B1(new_n632), .B2(new_n628), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(G330), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n567), .A2(new_n537), .A3(new_n515), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n636), .A2(new_n458), .A3(new_n449), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT30), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n562), .A2(new_n514), .A3(G179), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(new_n459), .A3(new_n537), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n637), .A2(new_n638), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n605), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(KEYINPUT31), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n572), .A2(new_n576), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n580), .B1(new_n483), .B2(new_n484), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n646), .A2(new_n647), .A3(new_n545), .A4(new_n607), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n644), .A2(KEYINPUT31), .ZN(new_n649));
  AOI211_X1 g0449(.A(new_n635), .B(new_n645), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n634), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n625), .B1(new_n653), .B2(G1), .ZN(G364));
  AOI21_X1  g0454(.A(new_n207), .B1(new_n599), .B2(G45), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n620), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n616), .B2(G330), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(G330), .B2(new_n616), .ZN(new_n659));
  OAI211_X1 g0459(.A(G1), .B(G13), .C1(new_n208), .C2(G169), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT93), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT93), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n208), .A2(G190), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(new_n337), .A3(new_n332), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n667), .A2(KEYINPUT94), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(KEYINPUT94), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G329), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n344), .A2(G179), .A3(G200), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(new_n208), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G294), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n208), .A2(new_n337), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(new_n344), .A3(new_n332), .ZN(new_n678));
  INV_X1    g0478(.A(G311), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n208), .A2(new_n344), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n332), .A2(G179), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI22_X1  g0482(.A1(new_n678), .A2(new_n679), .B1(new_n682), .B2(new_n560), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n665), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  AOI211_X1 g0485(.A(new_n267), .B(new_n683), .C1(G283), .C2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n677), .A2(G190), .A3(new_n332), .ZN(new_n687));
  INV_X1    g0487(.A(G322), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n337), .A2(new_n332), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n665), .ZN(new_n691));
  INV_X1    g0491(.A(G317), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n692), .A2(KEYINPUT33), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(KEYINPUT33), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n680), .A2(new_n690), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AOI211_X1 g0497(.A(new_n689), .B(new_n695), .C1(G326), .C2(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n672), .A2(new_n676), .A3(new_n686), .A4(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n267), .ZN(new_n700));
  INV_X1    g0500(.A(new_n318), .ZN(new_n701));
  OAI22_X1  g0501(.A1(new_n701), .A2(new_n687), .B1(new_n691), .B2(new_n289), .ZN(new_n702));
  AOI211_X1 g0502(.A(new_n700), .B(new_n702), .C1(G50), .C2(new_n697), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n667), .A2(G159), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n704), .A2(KEYINPUT32), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n704), .A2(KEYINPUT32), .B1(G97), .B2(new_n675), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n684), .A2(new_n355), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n682), .A2(new_n495), .ZN(new_n708));
  INV_X1    g0508(.A(new_n678), .ZN(new_n709));
  AOI211_X1 g0509(.A(new_n707), .B(new_n708), .C1(G77), .C2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n703), .A2(new_n705), .A3(new_n706), .A4(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n664), .B1(new_n699), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(G13), .A2(G33), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G20), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n663), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n619), .A2(new_n387), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n219), .A2(new_n450), .A3(G50), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n718), .B(new_n719), .C1(new_n249), .C2(new_n450), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n619), .A2(new_n700), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n721), .A2(G355), .B1(new_n531), .B2(new_n619), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n717), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n657), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n712), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n715), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n616), .B2(new_n726), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n659), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(G396));
  OAI21_X1  g0529(.A(new_n364), .B1(new_n353), .B2(new_n607), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n362), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n362), .A2(new_n605), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n630), .B(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n657), .B1(new_n735), .B2(new_n651), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n651), .B2(new_n735), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n663), .A2(new_n713), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n657), .B1(new_n739), .B2(G77), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n671), .A2(G311), .ZN(new_n741));
  INV_X1    g0541(.A(G283), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n678), .A2(new_n531), .B1(new_n691), .B2(new_n742), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n267), .B(new_n743), .C1(G87), .C2(new_n685), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n675), .A2(G97), .ZN(new_n745));
  INV_X1    g0545(.A(G294), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n687), .A2(new_n746), .B1(new_n682), .B2(new_n355), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(G303), .B2(new_n697), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n741), .A2(new_n744), .A3(new_n745), .A4(new_n748), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n709), .A2(G159), .B1(new_n697), .B2(G137), .ZN(new_n750));
  INV_X1    g0550(.A(G150), .ZN(new_n751));
  XOR2_X1   g0551(.A(KEYINPUT95), .B(G143), .Z(new_n752));
  OAI221_X1 g0552(.A(new_n750), .B1(new_n751), .B2(new_n691), .C1(new_n687), .C2(new_n752), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT34), .Z(new_n754));
  OAI22_X1  g0554(.A1(new_n682), .A2(new_n202), .B1(new_n684), .B2(new_n289), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n390), .B(new_n755), .C1(new_n318), .C2(new_n675), .ZN(new_n756));
  INV_X1    g0556(.A(G132), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n756), .B1(new_n757), .B2(new_n670), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n749), .B1(new_n754), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n740), .B1(new_n759), .B2(new_n663), .ZN(new_n760));
  INV_X1    g0560(.A(new_n734), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n760), .B1(new_n761), .B2(new_n714), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT96), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n737), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(G384));
  AOI211_X1 g0565(.A(new_n298), .B(new_n220), .C1(new_n318), .C2(G68), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n289), .A2(G50), .ZN(new_n767));
  OAI211_X1 g0567(.A(G1), .B(new_n287), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n469), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n769), .A2(KEYINPUT35), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(G116), .A3(new_n217), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(KEYINPUT35), .B2(new_n769), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n768), .B1(new_n772), .B2(KEYINPUT36), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(KEYINPUT36), .B2(new_n772), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT38), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT37), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n418), .B(new_n436), .C1(new_n412), .C2(new_n415), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n420), .A2(new_n429), .ZN(new_n779));
  INV_X1    g0579(.A(new_n603), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n420), .A2(new_n780), .ZN(new_n781));
  AND4_X1   g0581(.A1(new_n776), .A2(new_n778), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT99), .ZN(new_n783));
  INV_X1    g0583(.A(new_n398), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n381), .B1(new_n393), .B2(new_n397), .ZN(new_n785));
  AOI21_X1  g0585(.A(KEYINPUT16), .B1(new_n785), .B2(KEYINPUT97), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n388), .A2(G68), .A3(new_n392), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT79), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n396), .A2(KEYINPUT79), .A3(new_n392), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n380), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT97), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n294), .B1(new_n786), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT98), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n784), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n399), .B1(new_n791), .B2(new_n792), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n785), .A2(KEYINPUT97), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n293), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(KEYINPUT98), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n418), .B1(new_n796), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n783), .B1(new_n801), .B2(new_n603), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n795), .B(new_n293), .C1(new_n797), .C2(new_n798), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n398), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n786), .A2(new_n793), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n795), .B1(new_n805), .B2(new_n293), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n419), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n807), .A2(KEYINPUT99), .A3(new_n780), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n777), .B1(new_n807), .B2(new_n429), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n802), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n782), .B1(new_n810), .B2(KEYINPUT37), .ZN(new_n811));
  INV_X1    g0611(.A(new_n594), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n591), .A2(new_n812), .B1(new_n802), .B2(new_n808), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n775), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n808), .ZN(new_n815));
  AOI21_X1  g0615(.A(KEYINPUT99), .B1(new_n807), .B2(new_n780), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n440), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(KEYINPUT38), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n814), .B1(new_n811), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n309), .A2(new_n345), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n820), .A2(new_n308), .A3(new_n605), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n308), .A2(new_n605), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n309), .A2(new_n345), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n645), .B1(new_n648), .B2(new_n649), .ZN(new_n825));
  AND3_X1   g0625(.A1(new_n824), .A2(new_n825), .A3(new_n761), .ZN(new_n826));
  AOI21_X1  g0626(.A(KEYINPUT40), .B1(new_n819), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n778), .A2(new_n779), .A3(new_n781), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT37), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n440), .A2(new_n420), .A3(new_n780), .ZN(new_n830));
  AOI21_X1  g0630(.A(KEYINPUT38), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NOR3_X1   g0632(.A1(new_n818), .A2(new_n811), .A3(KEYINPUT100), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT100), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n810), .A2(KEYINPUT37), .ZN(new_n835));
  INV_X1    g0635(.A(new_n782), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n802), .A2(new_n808), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n775), .B1(new_n838), .B2(new_n440), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n834), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n832), .B1(new_n833), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n824), .A2(KEYINPUT40), .A3(new_n825), .A4(new_n761), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n841), .A2(KEYINPUT102), .A3(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT102), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n837), .A2(new_n834), .A3(new_n839), .ZN(new_n846));
  OAI21_X1  g0646(.A(KEYINPUT100), .B1(new_n818), .B2(new_n811), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n831), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n845), .B1(new_n848), .B2(new_n842), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n827), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n578), .A2(new_n825), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT103), .Z(new_n853));
  OR2_X1    g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n851), .A2(new_n853), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n854), .A2(G330), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n733), .B1(new_n630), .B2(new_n734), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n819), .A2(new_n824), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n591), .B2(new_n780), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n309), .A2(new_n605), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT39), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n861), .B(new_n832), .C1(new_n833), .C2(new_n840), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n859), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n597), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n633), .A2(new_n578), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT101), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n870));
  NOR4_X1   g0670(.A1(new_n870), .A2(new_n442), .A3(new_n868), .A4(new_n629), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n866), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n865), .B(new_n873), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n856), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n856), .A2(new_n874), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT104), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n875), .B1(new_n207), .B2(new_n599), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n774), .B1(new_n878), .B2(new_n880), .ZN(G367));
  INV_X1    g0681(.A(KEYINPUT42), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n478), .A2(new_n605), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n647), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT105), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n647), .A2(KEYINPUT105), .A3(new_n883), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n580), .A2(new_n605), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT106), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n610), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n882), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n890), .B1(new_n886), .B2(new_n887), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n895), .A2(KEYINPUT42), .A3(new_n610), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n488), .B1(new_n895), .B2(new_n575), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n607), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n542), .A2(new_n607), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n583), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n579), .A2(new_n901), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT43), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n904), .A2(KEYINPUT43), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n900), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n897), .A2(new_n906), .A3(new_n905), .A4(new_n899), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n895), .A2(new_n617), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n911), .B(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n620), .B(KEYINPUT41), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n895), .A2(new_n612), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT45), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n895), .A2(new_n612), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT44), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n918), .B(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n617), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT108), .ZN(new_n923));
  INV_X1    g0723(.A(new_n617), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT107), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT107), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n617), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n609), .B1(new_n586), .B2(new_n607), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n893), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n616), .A2(G330), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n925), .A2(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n634), .A2(new_n923), .A3(new_n651), .A4(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n931), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT108), .B1(new_n652), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n917), .A2(new_n617), .A3(new_n920), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n922), .A2(new_n932), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n915), .B1(new_n936), .B2(new_n653), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n913), .B1(new_n937), .B2(new_n656), .ZN(new_n938));
  INV_X1    g0738(.A(new_n718), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(new_n240), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n716), .B1(new_n211), .B2(new_n351), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n657), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n687), .A2(new_n751), .B1(new_n678), .B2(new_n202), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n684), .A2(new_n298), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(G137), .B2(new_n667), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n945), .B(new_n267), .C1(new_n701), .C2(new_n682), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n696), .A2(new_n752), .B1(new_n691), .B2(new_n373), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n674), .A2(new_n289), .ZN(new_n948));
  OR4_X1    g0748(.A1(new_n943), .A2(new_n946), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n682), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(G116), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT46), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n675), .A2(G107), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n709), .A2(G283), .B1(new_n697), .B2(G311), .ZN(new_n954));
  INV_X1    g0754(.A(new_n687), .ZN(new_n955));
  INV_X1    g0755(.A(new_n691), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n955), .A2(G303), .B1(new_n956), .B2(G294), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n952), .A2(new_n953), .A3(new_n954), .A4(new_n957), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n390), .B1(new_n271), .B2(new_n684), .C1(new_n692), .C2(new_n666), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT109), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n949), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT47), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n664), .B1(new_n961), .B2(new_n962), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n942), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n904), .B2(new_n726), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT110), .Z(new_n967));
  NAND2_X1  g0767(.A1(new_n938), .A2(new_n967), .ZN(G387));
  NOR2_X1   g0768(.A1(new_n609), .A2(new_n726), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n678), .A2(new_n289), .B1(new_n696), .B2(new_n373), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n751), .A2(new_n666), .B1(new_n682), .B2(new_n298), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n687), .A2(new_n202), .B1(new_n684), .B2(new_n271), .ZN(new_n972));
  OR4_X1    g0772(.A1(new_n390), .A2(new_n970), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n526), .A2(new_n674), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(new_n319), .C2(new_n956), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n955), .A2(G317), .B1(new_n956), .B2(G311), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n976), .B1(new_n560), .B2(new_n678), .C1(new_n688), .C2(new_n696), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT48), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n742), .B2(new_n674), .C1(new_n746), .C2(new_n682), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT49), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(G326), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n390), .B1(new_n531), .B2(new_n684), .C1(new_n982), .C2(new_n666), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(new_n979), .B2(new_n980), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n975), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n985), .A2(new_n664), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n348), .A2(new_n202), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT112), .Z(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(KEYINPUT50), .ZN(new_n989));
  AOI211_X1 g0789(.A(G45), .B(new_n623), .C1(G68), .C2(G77), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT111), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n988), .A2(KEYINPUT50), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n718), .B1(new_n450), .B2(new_n237), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n721), .A2(new_n623), .B1(new_n355), .B2(new_n619), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n717), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NOR4_X1   g0796(.A1(new_n969), .A2(new_n986), .A3(new_n724), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n931), .B2(new_n656), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n621), .B1(new_n934), .B2(new_n932), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n999), .A2(KEYINPUT113), .B1(new_n653), .B2(new_n931), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n999), .A2(KEYINPUT113), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(G393));
  INV_X1    g0802(.A(new_n935), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n1003), .A2(new_n921), .A3(new_n655), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n246), .A2(new_n939), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n717), .B1(G97), .B2(new_n619), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n724), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n687), .A2(new_n373), .B1(new_n696), .B2(new_n751), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT51), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n387), .B1(new_n289), .B2(new_n682), .C1(new_n495), .C2(new_n684), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n709), .A2(new_n348), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n202), .B2(new_n691), .C1(new_n666), .C2(new_n752), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1011), .B(new_n1013), .C1(G77), .C2(new_n675), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G283), .A2(new_n950), .B1(new_n956), .B2(G303), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n746), .B2(new_n678), .C1(new_n688), .C2(new_n666), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n674), .A2(new_n531), .ZN(new_n1017));
  NOR4_X1   g0817(.A1(new_n1016), .A2(new_n267), .A3(new_n707), .A4(new_n1017), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n687), .A2(new_n679), .B1(new_n696), .B2(new_n692), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT52), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1010), .A2(new_n1014), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1008), .B1(new_n664), .B2(new_n1021), .C1(new_n892), .C2(new_n726), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1004), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n936), .A2(new_n620), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n922), .A2(new_n935), .B1(new_n934), .B2(new_n932), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(G390));
  AOI21_X1  g0827(.A(new_n860), .B1(new_n857), .B2(new_n824), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n862), .A2(new_n863), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n841), .A2(new_n1028), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AND3_X1   g0832(.A1(new_n650), .A2(new_n761), .A3(new_n824), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n650), .A2(new_n761), .A3(new_n824), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1030), .A2(new_n1035), .A3(new_n1031), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n578), .A2(G330), .A3(new_n825), .ZN(new_n1037));
  AOI21_X1  g0837(.A(KEYINPUT101), .B1(new_n633), .B2(new_n578), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n597), .B(new_n1037), .C1(new_n1038), .C2(new_n871), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n824), .B1(new_n650), .B2(new_n761), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1041), .A2(new_n857), .A3(new_n1035), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n857), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n1033), .B2(new_n1040), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1039), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1034), .A2(new_n1036), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n620), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1039), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1045), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1048), .A2(KEYINPUT114), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT114), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1047), .A2(new_n1054), .A3(new_n620), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1034), .A2(new_n656), .A3(new_n1036), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n657), .B1(new_n739), .B2(new_n319), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n955), .A2(G132), .B1(new_n685), .B2(G50), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n682), .A2(new_n751), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1060), .A2(KEYINPUT53), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(KEYINPUT53), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n671), .A2(G125), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G128), .A2(new_n697), .B1(new_n956), .B2(G137), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(KEYINPUT54), .B(G143), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n267), .B1(new_n678), .B2(new_n1065), .C1(new_n674), .C2(new_n373), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  AND4_X1   g0867(.A1(new_n1059), .A2(new_n1063), .A3(new_n1064), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1069), .A2(KEYINPUT115), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n671), .A2(G294), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n675), .A2(G77), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n691), .A2(new_n355), .B1(new_n684), .B2(new_n289), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1073), .A2(new_n267), .A3(new_n708), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n678), .A2(new_n271), .B1(new_n696), .B2(new_n742), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G116), .B2(new_n955), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1069), .A2(KEYINPUT115), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1070), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1058), .B1(new_n1079), .B2(new_n663), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n864), .B2(new_n714), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1056), .A2(new_n1057), .A3(new_n1081), .ZN(G378));
  INV_X1    g0882(.A(G128), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n687), .A2(new_n1083), .B1(new_n691), .B2(new_n757), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n709), .A2(G137), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n697), .A2(G125), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(new_n682), .C2(new_n1065), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1084), .B(new_n1087), .C1(G150), .C2(new_n675), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT59), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n685), .A2(G159), .ZN(new_n1092));
  AOI211_X1 g0892(.A(G33), .B(G41), .C1(new_n667), .C2(G124), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(G50), .B1(new_n265), .B2(new_n452), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n387), .B2(G41), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT58), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n955), .A2(G107), .B1(new_n697), .B2(G116), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n685), .A2(new_n318), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(new_n271), .C2(new_n691), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n948), .B(new_n1100), .C1(G283), .C2(new_n671), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n390), .B(new_n452), .C1(new_n298), .C2(new_n682), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT116), .Z(new_n1103));
  OAI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(new_n526), .C2(new_n678), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1094), .B(new_n1096), .C1(new_n1097), .C2(new_n1104), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1104), .A2(new_n1097), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n663), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1107), .B(new_n657), .C1(G50), .C2(new_n739), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n341), .B(KEYINPUT55), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n325), .A2(new_n780), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1109), .B(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1111), .B(new_n1112), .Z(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1108), .B1(new_n1114), .B2(new_n713), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT118), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n827), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT102), .B1(new_n841), .B2(new_n843), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n848), .A2(new_n845), .A3(new_n842), .ZN(new_n1119));
  OAI211_X1 g0919(.A(G330), .B(new_n1117), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1120), .A2(new_n1114), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1113), .B1(new_n850), .B2(G330), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1116), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n865), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1120), .A2(new_n1114), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n850), .A2(G330), .A3(new_n1113), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n865), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1127), .A2(new_n1116), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1115), .B1(new_n1130), .B2(new_n656), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT57), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1125), .A2(new_n865), .A3(new_n1126), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n865), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT119), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1133), .B(KEYINPUT119), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(new_n620), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1141));
  AOI21_X1  g0941(.A(KEYINPUT57), .B1(new_n1130), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1131), .B1(new_n1140), .B2(new_n1142), .ZN(G375));
  AOI21_X1  g0943(.A(new_n724), .B1(new_n738), .B2(new_n289), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n955), .A2(G283), .B1(new_n956), .B2(G116), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1145), .B1(new_n355), .B2(new_n678), .C1(new_n746), .C2(new_n696), .ZN(new_n1146));
  NOR4_X1   g0946(.A1(new_n974), .A2(new_n267), .A3(new_n944), .A4(new_n1146), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n670), .A2(new_n560), .B1(new_n271), .B2(new_n682), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT121), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n670), .A2(new_n1083), .B1(new_n373), .B2(new_n682), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT122), .Z(new_n1151));
  OAI211_X1 g0951(.A(new_n1099), .B(new_n387), .C1(new_n751), .C2(new_n678), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n955), .A2(G137), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1153), .B1(new_n757), .B2(new_n696), .C1(new_n691), .C2(new_n1065), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1152), .B(new_n1154), .C1(G50), .C2(new_n675), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1147), .A2(new_n1149), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1144), .B1(new_n664), .B2(new_n1156), .C1(new_n824), .C2(new_n714), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n1045), .B2(new_n655), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n914), .B(KEYINPUT120), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1052), .A2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1159), .B1(new_n1161), .B2(new_n1162), .ZN(G381));
  OR2_X1    g0963(.A1(G375), .A2(G378), .ZN(new_n1164));
  OR3_X1    g0964(.A1(G390), .A2(G381), .A3(G384), .ZN(new_n1165));
  OR4_X1    g0965(.A1(G396), .A2(new_n1165), .A3(G387), .A4(G393), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n1164), .A2(new_n1166), .ZN(G407));
  OAI211_X1 g0967(.A(G407), .B(G213), .C1(G343), .C2(new_n1164), .ZN(G409));
  INV_X1    g0968(.A(KEYINPUT61), .ZN(new_n1169));
  INV_X1    g0969(.A(G213), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1170), .A2(G343), .ZN(new_n1171));
  OAI211_X1 g0971(.A(G378), .B(new_n1131), .C1(new_n1140), .C2(new_n1142), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1130), .A2(new_n1141), .A3(new_n1160), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1135), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1125), .A2(new_n865), .A3(new_n1126), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1115), .B1(new_n1176), .B2(new_n656), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1173), .A2(new_n1177), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1056), .A2(new_n1057), .A3(new_n1081), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1171), .B1(new_n1172), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1171), .A2(G2897), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1052), .A2(new_n620), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT60), .B1(new_n1039), .B2(new_n1045), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1162), .A2(KEYINPUT60), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(G384), .B1(new_n1187), .B2(new_n1159), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n764), .B(new_n1158), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1188), .A2(new_n1189), .A3(KEYINPUT123), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT123), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n1162), .A2(KEYINPUT60), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1192), .A2(new_n1184), .A3(new_n1183), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n764), .B1(new_n1193), .B2(new_n1158), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1187), .A2(G384), .A3(new_n1159), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1191), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1182), .B1(new_n1190), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1198));
  OAI211_X1 g0998(.A(G2897), .B(new_n1171), .C1(new_n1198), .C2(KEYINPUT123), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1169), .B1(new_n1181), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1181), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT63), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(G393), .B(new_n728), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n938), .A2(new_n967), .A3(G390), .ZN(new_n1208));
  AOI21_X1  g1008(.A(G390), .B1(new_n938), .B2(new_n967), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1208), .B1(new_n1209), .B2(KEYINPUT124), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT124), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1211), .B(G390), .C1(new_n938), .C2(new_n967), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1207), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT125), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(KEYINPUT125), .B(new_n1207), .C1(new_n1210), .C2(new_n1212), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1209), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1217), .A2(KEYINPUT126), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1208), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1207), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1217), .A2(KEYINPUT126), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1218), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1215), .A2(new_n1216), .A3(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1181), .A2(KEYINPUT63), .A3(new_n1203), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1202), .A2(new_n1206), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT62), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1181), .A2(new_n1226), .A3(new_n1203), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1226), .B1(new_n1181), .B2(new_n1203), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1227), .A2(new_n1201), .A3(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1225), .B1(new_n1229), .B2(new_n1223), .ZN(G405));
  INV_X1    g1030(.A(KEYINPUT127), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1203), .A2(new_n1231), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1223), .B(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1172), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n1231), .B2(new_n1203), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(G375), .A2(new_n1179), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1233), .A2(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1223), .A2(new_n1232), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1223), .A2(new_n1232), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1239), .A2(new_n1236), .A3(new_n1235), .A4(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1238), .A2(new_n1241), .ZN(G402));
endmodule


