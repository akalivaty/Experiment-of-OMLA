//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n562, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n622, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT66), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  NOR2_X1   g051(.A1(new_n466), .A2(G2105), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  NOR2_X1   g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n479), .B(new_n480), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT69), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n463), .A2(new_n465), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n484), .A2(new_n485), .A3(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT67), .B1(new_n466), .B2(new_n473), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI211_X1 g063(.A(new_n478), .B(new_n483), .C1(G124), .C2(new_n488), .ZN(G162));
  NAND2_X1  g064(.A1(G114), .A2(G2104), .ZN(new_n490));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n466), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n477), .A2(G138), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n484), .A2(KEYINPUT4), .A3(G138), .ZN(new_n496));
  NAND2_X1  g071(.A1(G102), .A2(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n494), .A2(new_n495), .B1(new_n473), .B2(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT71), .B1(new_n502), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(new_n500), .A3(KEYINPUT5), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT70), .B1(new_n509), .B2(G651), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(new_n507), .A3(KEYINPUT6), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n508), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n519), .A2(new_n507), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n518), .A2(new_n520), .ZN(G166));
  NAND2_X1  g096(.A1(G63), .A2(G651), .ZN(new_n522));
  INV_X1    g097(.A(new_n501), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n504), .B1(KEYINPUT5), .B2(new_n500), .ZN(new_n524));
  NOR3_X1   g099(.A1(new_n502), .A2(KEYINPUT71), .A3(G543), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT72), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n506), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n522), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n506), .A2(new_n513), .A3(G89), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n513), .A2(G51), .A3(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NOR3_X1   g111(.A1(new_n530), .A2(new_n533), .A3(new_n536), .ZN(G168));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n538), .B1(new_n527), .B2(new_n529), .ZN(new_n539));
  INV_X1    g114(.A(G77), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n500), .ZN(new_n541));
  OAI21_X1  g116(.A(G651), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n516), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n506), .A2(new_n513), .ZN(new_n544));
  XOR2_X1   g119(.A(KEYINPUT74), .B(G90), .Z(new_n545));
  AOI22_X1  g120(.A1(G52), .A2(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n542), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  AOI211_X1 g123(.A(KEYINPUT72), .B(new_n501), .C1(new_n503), .C2(new_n505), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n503), .A2(new_n505), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n528), .B1(new_n550), .B2(new_n523), .ZN(new_n551));
  OAI21_X1  g126(.A(G56), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(G68), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n500), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n507), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(G81), .ZN(new_n557));
  INV_X1    g132(.A(G43), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n514), .A2(new_n557), .B1(new_n516), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G188));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  INV_X1    g142(.A(G53), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n516), .B2(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n513), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G91), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n572), .A2(new_n507), .B1(new_n514), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G299));
  INV_X1    g151(.A(new_n522), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n577), .B1(new_n549), .B2(new_n551), .ZN(new_n578));
  INV_X1    g153(.A(new_n536), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n578), .A2(new_n532), .A3(new_n531), .A4(new_n579), .ZN(G286));
  INV_X1    g155(.A(G166), .ZN(G303));
  NAND2_X1  g156(.A1(new_n527), .A2(new_n529), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n582), .B2(G74), .ZN(new_n583));
  AOI22_X1  g158(.A1(G49), .A2(new_n543), .B1(new_n544), .B2(G87), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G288));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  INV_X1    g161(.A(G48), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n514), .A2(new_n586), .B1(new_n516), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n506), .A2(G61), .ZN(new_n589));
  AND2_X1   g164(.A1(G73), .A2(G543), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT75), .Z(new_n591));
  AOI21_X1  g166(.A(new_n507), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(G47), .A2(new_n543), .B1(new_n544), .B2(G85), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n582), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(new_n507), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT76), .B1(new_n514), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT76), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n506), .A2(new_n513), .A3(new_n601), .A4(G92), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n600), .A2(KEYINPUT10), .A3(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(KEYINPUT10), .B1(new_n600), .B2(new_n602), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g181(.A(KEYINPUT79), .B(G66), .Z(new_n607));
  NAND2_X1  g182(.A1(new_n506), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT78), .Z(new_n610));
  AOI21_X1  g185(.A(new_n507), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT77), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n516), .B(new_n612), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n611), .B1(new_n613), .B2(G54), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n606), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n598), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n598), .B1(new_n616), .B2(G868), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n575), .ZN(G297));
  OAI21_X1  g195(.A(new_n619), .B1(G868), .B2(new_n575), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n616), .B1(new_n622), .B2(G860), .ZN(G148));
  NOR2_X1   g198(.A1(new_n560), .A2(G868), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n616), .A2(new_n622), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT80), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g203(.A1(new_n488), .A2(G123), .B1(G135), .B2(new_n477), .ZN(new_n629));
  NOR2_X1   g204(.A1(G99), .A2(G2105), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(new_n473), .B2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT81), .B(G2096), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n473), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2100), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n634), .A2(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2435), .ZN(new_n641));
  XOR2_X1   g216(.A(G2427), .B(G2438), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT14), .ZN(new_n644));
  XOR2_X1   g219(.A(G2451), .B(G2454), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n644), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G1341), .B(G1348), .Z(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT82), .Z(new_n652));
  INV_X1    g227(.A(G14), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n649), .B2(new_n650), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2067), .B(G2678), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT83), .ZN(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n658), .A2(new_n659), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n659), .B(KEYINPUT17), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n664), .B(new_n661), .C1(new_n658), .C2(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n658), .A2(new_n665), .A3(new_n660), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT86), .ZN(new_n676));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT20), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n673), .A2(new_n674), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT87), .ZN(new_n683));
  INV_X1    g258(.A(new_n681), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(new_n675), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n680), .B(new_n683), .C1(new_n678), .C2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1991), .B(G1996), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT88), .B(G1986), .ZN(new_n691));
  INV_X1    g266(.A(G1981), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n690), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  NOR2_X1   g271(.A1(G16), .A2(G22), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G166), .B2(G16), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1971), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G6), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n593), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT32), .B(G1981), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n700), .A2(G23), .ZN(new_n706));
  INV_X1    g281(.A(G288), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(new_n700), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT91), .B(KEYINPUT92), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT33), .B(G1976), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n708), .A2(new_n710), .ZN(new_n713));
  AND3_X1   g288(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n712), .B1(new_n711), .B2(new_n713), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n705), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(KEYINPUT34), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G25), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n477), .A2(G131), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT89), .Z(new_n721));
  OAI21_X1  g296(.A(KEYINPUT90), .B1(G95), .B2(G2105), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(G2104), .B1(new_n473), .B2(G107), .ZN(new_n724));
  NOR3_X1   g299(.A1(KEYINPUT90), .A2(G95), .A3(G2105), .ZN(new_n725));
  NOR3_X1   g300(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n488), .B2(G119), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n721), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n719), .B1(new_n729), .B2(new_n718), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT35), .B(G1991), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n730), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n700), .A2(G24), .ZN(new_n734));
  INV_X1    g309(.A(G290), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n700), .ZN(new_n736));
  INV_X1    g311(.A(G1986), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n733), .B(new_n738), .C1(new_n716), .C2(KEYINPUT34), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n739), .A2(KEYINPUT93), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(KEYINPUT93), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n717), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(KEYINPUT36), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT36), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n744), .B(new_n717), .C1(new_n740), .C2(new_n741), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n718), .A2(G35), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G162), .B2(new_n718), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2090), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT105), .B(KEYINPUT29), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n700), .A2(G4), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n615), .B2(G16), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1348), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT28), .ZN(new_n755));
  INV_X1    g330(.A(G26), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(G29), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(G29), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n488), .A2(G128), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(KEYINPUT94), .ZN(new_n760));
  OR2_X1    g335(.A1(G104), .A2(G2105), .ZN(new_n761));
  INV_X1    g336(.A(G116), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n462), .B1(new_n762), .B2(G2105), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n477), .A2(G140), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT94), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n488), .A2(new_n765), .A3(G128), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n760), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n758), .B1(new_n767), .B2(G29), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n757), .B1(new_n768), .B2(new_n755), .ZN(new_n769));
  INV_X1    g344(.A(G2067), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n700), .A2(G19), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n560), .B2(new_n700), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(G1341), .Z(new_n774));
  NAND3_X1  g349(.A1(new_n754), .A2(new_n771), .A3(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT95), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n754), .A2(new_n771), .A3(KEYINPUT95), .A4(new_n774), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n718), .A2(G33), .ZN(new_n780));
  NAND2_X1  g355(.A1(G115), .A2(G2104), .ZN(new_n781));
  INV_X1    g356(.A(G127), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n466), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G2105), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT96), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n477), .A2(G139), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT25), .Z(new_n789));
  NAND3_X1  g364(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT97), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n780), .B1(new_n792), .B2(new_n718), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(G2072), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT98), .Z(new_n795));
  NOR2_X1   g370(.A1(G164), .A2(new_n718), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G27), .B2(new_n718), .ZN(new_n797));
  INV_X1    g372(.A(G2078), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT99), .ZN(new_n799));
  NOR2_X1   g374(.A1(KEYINPUT24), .A2(G34), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(KEYINPUT24), .A2(G34), .ZN(new_n802));
  AOI21_X1  g377(.A(G29), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI22_X1  g378(.A1(G160), .A2(G29), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n799), .B2(new_n803), .ZN(new_n805));
  INV_X1    g380(.A(G2084), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI22_X1  g382(.A1(new_n797), .A2(new_n798), .B1(KEYINPUT104), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n798), .B2(new_n797), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n700), .A2(KEYINPUT23), .A3(G20), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT23), .ZN(new_n811));
  INV_X1    g386(.A(G20), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(G16), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n810), .B(new_n813), .C1(new_n575), .C2(new_n700), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(G1956), .Z(new_n815));
  NAND4_X1  g390(.A1(new_n779), .A2(new_n795), .A3(new_n809), .A4(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT102), .B1(G5), .B2(G16), .ZN(new_n817));
  OR3_X1    g392(.A1(KEYINPUT102), .A2(G5), .A3(G16), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n817), .B(new_n818), .C1(G301), .C2(new_n700), .ZN(new_n819));
  INV_X1    g394(.A(G1961), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n805), .A2(new_n806), .ZN(new_n823));
  NOR2_X1   g398(.A1(G29), .A2(G32), .ZN(new_n824));
  NAND3_X1  g399(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT26), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(new_n488), .B2(G129), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n473), .A2(G105), .A3(G2104), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n477), .A2(G141), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n824), .B1(new_n831), .B2(G29), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT27), .B(G1996), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(KEYINPUT104), .B2(new_n807), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NOR4_X1   g412(.A1(new_n816), .A2(new_n822), .A3(new_n823), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n793), .A2(G2072), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT100), .Z(new_n840));
  NAND4_X1  g415(.A1(new_n746), .A2(new_n751), .A3(new_n838), .A4(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT30), .B(G28), .ZN(new_n842));
  OR2_X1    g417(.A1(KEYINPUT31), .A2(G11), .ZN(new_n843));
  NAND2_X1  g418(.A1(KEYINPUT31), .A2(G11), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n842), .A2(new_n718), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n632), .B2(new_n718), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT101), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n700), .A2(G21), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(G168), .B2(new_n700), .ZN(new_n849));
  INV_X1    g424(.A(G1966), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n847), .B(new_n851), .C1(new_n820), .C2(new_n819), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT103), .Z(new_n853));
  NOR2_X1   g428(.A1(new_n841), .A2(new_n853), .ZN(G311));
  NOR3_X1   g429(.A1(new_n816), .A2(new_n823), .A3(new_n837), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n821), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n743), .B2(new_n745), .ZN(new_n857));
  INV_X1    g432(.A(new_n853), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n857), .A2(new_n858), .A3(new_n751), .A4(new_n840), .ZN(G150));
  OAI21_X1  g434(.A(G67), .B1(new_n549), .B2(new_n551), .ZN(new_n860));
  INV_X1    g435(.A(G80), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n861), .A2(new_n500), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n507), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(G93), .ZN(new_n865));
  INV_X1    g440(.A(G55), .ZN(new_n866));
  OAI22_X1  g441(.A1(new_n514), .A2(new_n865), .B1(new_n516), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(G860), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT37), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n616), .A2(G559), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT39), .ZN(new_n873));
  XNOR2_X1  g448(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G56), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(new_n527), .B2(new_n529), .ZN(new_n877));
  OAI21_X1  g452(.A(G651), .B1(new_n877), .B2(new_n554), .ZN(new_n878));
  INV_X1    g453(.A(new_n559), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n878), .B(new_n879), .C1(new_n864), .C2(new_n867), .ZN(new_n880));
  INV_X1    g455(.A(G67), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n881), .B1(new_n527), .B2(new_n529), .ZN(new_n882));
  OAI21_X1  g457(.A(G651), .B1(new_n882), .B2(new_n862), .ZN(new_n883));
  INV_X1    g458(.A(new_n867), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n883), .B(new_n884), .C1(new_n556), .C2(new_n559), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n875), .B(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n871), .B1(new_n887), .B2(G860), .ZN(G145));
  AOI22_X1  g463(.A1(new_n488), .A2(G130), .B1(G142), .B2(new_n477), .ZN(new_n889));
  NOR2_X1   g464(.A1(G106), .A2(G2105), .ZN(new_n890));
  OAI21_X1  g465(.A(G2104), .B1(new_n473), .B2(G118), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n636), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT107), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n767), .A2(G164), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n494), .A2(new_n495), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n498), .A2(new_n473), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n899), .A2(new_n764), .A3(new_n760), .A4(new_n766), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n831), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n896), .A2(new_n900), .A3(new_n831), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n895), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n903), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n905), .A2(KEYINPUT107), .A3(new_n901), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n792), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT108), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n902), .A2(new_n790), .A3(new_n903), .ZN(new_n910));
  OAI211_X1 g485(.A(KEYINPUT108), .B(new_n792), .C1(new_n906), .C2(new_n904), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n729), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n632), .B(G160), .ZN(new_n914));
  XNOR2_X1  g489(.A(G162), .B(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n909), .A2(new_n728), .A3(new_n910), .A4(new_n911), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n916), .B1(new_n913), .B2(new_n917), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n894), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n913), .A2(new_n917), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n915), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n923), .A2(new_n893), .A3(new_n918), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n921), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT40), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT40), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n921), .A2(new_n924), .A3(new_n928), .A4(new_n925), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(G395));
  INV_X1    g505(.A(G868), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n735), .A2(G288), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n707), .A2(G290), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT109), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n932), .A2(KEYINPUT109), .A3(new_n933), .ZN(new_n937));
  XNOR2_X1  g512(.A(G166), .B(new_n593), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n934), .A2(new_n935), .A3(new_n938), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT42), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n941), .A2(KEYINPUT42), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT110), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n941), .A2(KEYINPUT42), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(new_n947), .A3(new_n942), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n625), .B(new_n886), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n575), .B1(new_n606), .B2(new_n614), .ZN(new_n950));
  INV_X1    g525(.A(new_n605), .ZN(new_n951));
  AND4_X1   g526(.A1(new_n575), .A2(new_n614), .A3(new_n603), .A4(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n949), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n615), .A2(G299), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n606), .A2(new_n575), .A3(new_n614), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(KEYINPUT41), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT41), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(new_n950), .B2(new_n952), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n949), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n945), .A2(new_n948), .A3(new_n954), .A4(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n954), .ZN(new_n964));
  OAI221_X1 g539(.A(KEYINPUT110), .B1(new_n964), .B2(new_n961), .C1(new_n943), .C2(new_n944), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n931), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n869), .A2(G868), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(G295));
  OR3_X1    g543(.A1(new_n966), .A2(KEYINPUT111), .A3(new_n967), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT111), .B1(new_n966), .B2(new_n967), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(G331));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n972));
  OAI21_X1  g547(.A(G64), .B1(new_n549), .B2(new_n551), .ZN(new_n973));
  INV_X1    g548(.A(new_n541), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n507), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n544), .A2(new_n545), .ZN(new_n976));
  INV_X1    g551(.A(G52), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n976), .B1(new_n977), .B2(new_n516), .ZN(new_n978));
  OAI21_X1  g553(.A(G168), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n542), .A2(G286), .A3(new_n546), .ZN(new_n980));
  AND4_X1   g555(.A1(new_n880), .A2(new_n885), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n880), .A2(new_n885), .B1(new_n979), .B2(new_n980), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT112), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT112), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n979), .A2(new_n980), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n984), .B1(new_n886), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n983), .A2(new_n953), .A3(new_n986), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n957), .B(new_n959), .C1(new_n981), .C2(new_n982), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n987), .A2(KEYINPUT113), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT113), .B1(new_n987), .B2(new_n988), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n989), .A2(new_n990), .A3(new_n941), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n972), .B1(new_n991), .B2(G37), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n941), .A2(new_n988), .A3(new_n987), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n987), .A2(new_n988), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n939), .A2(new_n940), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n987), .A2(new_n988), .A3(KEYINPUT113), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n999), .A2(KEYINPUT114), .A3(new_n925), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n992), .A2(KEYINPUT43), .A3(new_n993), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n960), .B1(new_n983), .B2(new_n986), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n981), .A2(new_n982), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1003), .B1(new_n953), .B2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n925), .B(new_n993), .C1(new_n1005), .C2(new_n941), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1001), .A2(new_n1002), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT115), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1001), .A2(new_n1011), .A3(new_n1002), .A4(new_n1008), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n992), .A2(new_n1007), .A3(new_n993), .A4(new_n1000), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1006), .A2(KEYINPUT43), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(KEYINPUT44), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1013), .A2(new_n1016), .ZN(G397));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(G164), .B2(G1384), .ZN(new_n1019));
  NAND2_X1  g594(.A1(G160), .A2(G40), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1996), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g598(.A(new_n1023), .B(KEYINPUT46), .Z(new_n1024));
  XNOR2_X1  g599(.A(new_n767), .B(G2067), .ZN(new_n1025));
  OR2_X1    g600(.A1(new_n1025), .A2(new_n830), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1024), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1027), .B(KEYINPUT126), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1028), .B(KEYINPUT47), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n830), .B(G1996), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n728), .A2(new_n731), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  OAI22_X1  g608(.A1(new_n1031), .A2(new_n1033), .B1(G2067), .B2(new_n767), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n1021), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1035), .B(KEYINPUT125), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n735), .A2(new_n737), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1037), .B(KEYINPUT116), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1021), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1039), .B(KEYINPUT48), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1021), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n729), .A2(new_n732), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1031), .A2(new_n1042), .A3(new_n1032), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1040), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1029), .A2(new_n1036), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  NOR2_X1   g622(.A1(G166), .A2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1048), .B(KEYINPUT55), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT118), .ZN(new_n1051));
  INV_X1    g626(.A(G1384), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n899), .A2(KEYINPUT45), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1020), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1019), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G1971), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(G164), .B2(G1384), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NOR3_X1   g635(.A1(G164), .A2(new_n1058), .A3(G1384), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1054), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1057), .B1(new_n1062), .B2(G2090), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1049), .A2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1051), .A2(G8), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1384), .B1(new_n897), .B2(new_n898), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1047), .B1(new_n1054), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n707), .A2(G1976), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT52), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n588), .A2(new_n592), .A3(G1981), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(G1981), .B1(new_n588), .B2(new_n592), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1073), .A2(KEYINPUT49), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT49), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1074), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1076), .B1(new_n1077), .B2(new_n1072), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1068), .A2(new_n1075), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1976), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT52), .B1(G288), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1068), .A2(new_n1069), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1071), .A2(new_n1079), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1068), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G288), .A2(G1976), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(KEYINPUT119), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1072), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n1066), .A2(new_n1083), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1348), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1062), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1054), .A2(new_n1067), .A3(new_n770), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n615), .A2(KEYINPUT60), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1053), .A2(new_n1019), .A3(new_n1022), .A4(new_n1054), .ZN(new_n1095));
  XOR2_X1   g670(.A(KEYINPUT58), .B(G1341), .Z(new_n1096));
  NAND2_X1  g671(.A1(new_n899), .A2(new_n1052), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1096), .B1(new_n1097), .B2(new_n1020), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT59), .B1(new_n1099), .B2(new_n560), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1099), .A2(KEYINPUT59), .A3(new_n560), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1094), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n575), .B(KEYINPUT57), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT56), .B(G2072), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1053), .A2(new_n1019), .A3(new_n1054), .A4(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n899), .A2(KEYINPUT50), .A3(new_n1052), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1020), .B1(new_n1106), .B2(new_n1059), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1103), .B(new_n1105), .C1(new_n1107), .C2(G1956), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1108), .A2(new_n1109), .A3(KEYINPUT61), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n1108), .B2(KEYINPUT61), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1108), .A2(KEYINPUT61), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n615), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n615), .B(new_n1092), .C1(new_n1107), .C2(G1348), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT60), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1102), .A2(new_n1112), .A3(new_n1113), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1114), .A2(new_n1108), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1105), .B1(new_n1107), .B2(G1956), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1103), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1118), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT51), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1020), .B1(new_n1097), .B2(new_n1018), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1067), .A2(KEYINPUT120), .A3(KEYINPUT45), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1053), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n850), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1107), .A2(new_n806), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1130), .A2(G168), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1124), .B1(new_n1132), .B2(G8), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(G286), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT51), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1132), .A2(G8), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1133), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1063), .A2(G8), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1083), .B1(new_n1139), .B2(new_n1050), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1062), .A2(new_n820), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT53), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1055), .B2(G2078), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1142), .A2(G2078), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1141), .B(new_n1143), .C1(new_n1145), .C2(new_n1129), .ZN(new_n1146));
  XOR2_X1   g721(.A(G301), .B(KEYINPUT54), .Z(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1125), .A2(new_n1053), .A3(new_n1144), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1141), .A2(new_n1143), .A3(new_n1147), .A4(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1140), .A2(new_n1149), .A3(new_n1066), .A4(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1138), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1089), .B1(new_n1123), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1047), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1140), .A2(G168), .A3(new_n1066), .A4(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1158), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1154), .A2(new_n1155), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1155), .B1(new_n1154), .B2(new_n1164), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT124), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1167), .B1(new_n1138), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1132), .A2(G8), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(KEYINPUT51), .B2(new_n1135), .ZN(new_n1171));
  OAI211_X1 g746(.A(KEYINPUT124), .B(KEYINPUT62), .C1(new_n1171), .C2(new_n1133), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1169), .A2(new_n1172), .A3(new_n1066), .A4(new_n1140), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1138), .A2(new_n1168), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1174), .A2(G171), .A3(new_n1146), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1165), .A2(new_n1166), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(G290), .A2(G1986), .ZN(new_n1178));
  XOR2_X1   g753(.A(new_n1178), .B(KEYINPUT117), .Z(new_n1179));
  NOR2_X1   g754(.A1(new_n1038), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1041), .B1(new_n1043), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1046), .B1(new_n1177), .B2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g757(.A1(new_n1001), .A2(new_n1008), .ZN(new_n1184));
  NOR2_X1   g758(.A1(G227), .A2(new_n459), .ZN(new_n1185));
  NAND3_X1  g759(.A1(new_n695), .A2(new_n655), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n1187));
  OR2_X1    g761(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1189));
  AND4_X1   g763(.A1(new_n926), .A2(new_n1184), .A3(new_n1188), .A4(new_n1189), .ZN(G308));
  NAND4_X1  g764(.A1(new_n926), .A2(new_n1184), .A3(new_n1188), .A4(new_n1189), .ZN(G225));
endmodule


