

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767;

  NOR2_X1 U374 ( .A1(n544), .A2(n543), .ZN(n690) );
  AND2_X1 U375 ( .A1(n417), .A2(n416), .ZN(n415) );
  INV_X2 U376 ( .A(G953), .ZN(n759) );
  XOR2_X1 U377 ( .A(n408), .B(n407), .Z(n354) );
  NAND2_X2 U378 ( .A1(n415), .A2(n411), .ZN(n660) );
  NAND2_X2 U379 ( .A1(n387), .A2(n386), .ZN(n385) );
  XNOR2_X2 U380 ( .A(n495), .B(n482), .ZN(n464) );
  XNOR2_X2 U381 ( .A(n563), .B(n562), .ZN(n612) );
  AND2_X1 U382 ( .A1(n393), .A2(n605), .ZN(n392) );
  AND2_X1 U383 ( .A1(n607), .A2(n634), .ZN(n613) );
  OR2_X1 U384 ( .A1(n537), .A2(n546), .ZN(n472) );
  NOR2_X1 U385 ( .A1(n537), .A2(n575), .ZN(n576) );
  XNOR2_X1 U386 ( .A(n354), .B(n465), .ZN(n645) );
  OR2_X2 U387 ( .A1(n758), .A2(KEYINPUT72), .ZN(n355) );
  AND2_X1 U388 ( .A1(n371), .A2(n370), .ZN(n600) );
  AND2_X1 U389 ( .A1(n372), .A2(n598), .ZN(n371) );
  XNOR2_X1 U390 ( .A(n428), .B(G137), .ZN(n437) );
  INV_X1 U391 ( .A(G140), .ZN(n428) );
  OR2_X1 U392 ( .A1(n674), .A2(G902), .ZN(n436) );
  XNOR2_X1 U393 ( .A(n423), .B(KEYINPUT68), .ZN(n422) );
  INV_X1 U394 ( .A(KEYINPUT10), .ZN(n423) );
  AND2_X1 U395 ( .A1(n473), .A2(n718), .ZN(n424) );
  OR2_X1 U396 ( .A1(n549), .A2(n546), .ZN(n584) );
  XNOR2_X1 U397 ( .A(n532), .B(n531), .ZN(n539) );
  XNOR2_X1 U398 ( .A(KEYINPUT93), .B(KEYINPUT20), .ZN(n405) );
  NOR2_X1 U399 ( .A1(G953), .A2(G237), .ZN(n474) );
  XNOR2_X1 U400 ( .A(n603), .B(KEYINPUT48), .ZN(n399) );
  NOR2_X1 U401 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U402 ( .A(n382), .B(n381), .ZN(n500) );
  XNOR2_X1 U403 ( .A(G116), .B(G113), .ZN(n382) );
  XNOR2_X1 U404 ( .A(G119), .B(KEYINPUT3), .ZN(n381) );
  XNOR2_X1 U405 ( .A(n369), .B(n368), .ZN(n494) );
  INV_X1 U406 ( .A(KEYINPUT8), .ZN(n368) );
  NAND2_X1 U407 ( .A1(n759), .A2(G234), .ZN(n369) );
  INV_X1 U408 ( .A(G122), .ZN(n481) );
  XNOR2_X1 U409 ( .A(KEYINPUT69), .B(G131), .ZN(n482) );
  NAND2_X1 U410 ( .A1(n355), .A2(n425), .ZN(n388) );
  XNOR2_X1 U411 ( .A(n555), .B(n554), .ZN(n727) );
  XNOR2_X1 U412 ( .A(n527), .B(n357), .ZN(n556) );
  XNOR2_X1 U413 ( .A(n439), .B(n441), .ZN(n420) );
  XNOR2_X1 U414 ( .A(G116), .B(G107), .ZN(n493) );
  XNOR2_X1 U415 ( .A(G122), .B(KEYINPUT7), .ZN(n490) );
  XOR2_X1 U416 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n491) );
  INV_X1 U417 ( .A(G134), .ZN(n427) );
  XNOR2_X1 U418 ( .A(G104), .B(KEYINPUT89), .ZN(n429) );
  XNOR2_X1 U419 ( .A(n464), .B(n437), .ZN(n756) );
  AND2_X1 U420 ( .A1(n379), .A2(n553), .ZN(n545) );
  AND2_X1 U421 ( .A1(n690), .A2(n380), .ZN(n379) );
  INV_X1 U422 ( .A(n575), .ZN(n380) );
  OR2_X1 U423 ( .A1(n651), .A2(n513), .ZN(n518) );
  NAND2_X1 U424 ( .A1(n667), .A2(n496), .ZN(n498) );
  XNOR2_X1 U425 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U426 ( .A(n445), .B(n401), .ZN(n400) );
  XNOR2_X1 U427 ( .A(n444), .B(n446), .ZN(n401) );
  INV_X1 U428 ( .A(KEYINPUT1), .ZN(n367) );
  AND2_X1 U429 ( .A1(n539), .A2(n538), .ZN(n567) );
  INV_X1 U430 ( .A(G237), .ZN(n470) );
  XNOR2_X1 U431 ( .A(n406), .B(n403), .ZN(n447) );
  XNOR2_X1 U432 ( .A(n405), .B(n404), .ZN(n403) );
  INV_X1 U433 ( .A(KEYINPUT92), .ZN(n404) );
  NAND2_X1 U434 ( .A1(n395), .A2(n394), .ZN(n393) );
  INV_X1 U435 ( .A(KEYINPUT79), .ZN(n394) );
  INV_X1 U436 ( .A(n604), .ZN(n395) );
  AND2_X1 U437 ( .A1(n604), .A2(KEYINPUT79), .ZN(n397) );
  XOR2_X1 U438 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n475) );
  XNOR2_X1 U439 ( .A(G143), .B(G113), .ZN(n477) );
  XOR2_X1 U440 ( .A(KEYINPUT97), .B(G140), .Z(n478) );
  XNOR2_X1 U441 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n503) );
  NAND2_X1 U442 ( .A1(G234), .A2(G237), .ZN(n449) );
  XNOR2_X1 U443 ( .A(n549), .B(KEYINPUT38), .ZN(n718) );
  OR2_X1 U444 ( .A1(n706), .A2(n705), .ZN(n620) );
  INV_X1 U445 ( .A(G902), .ZN(n496) );
  XNOR2_X1 U446 ( .A(n383), .B(n500), .ZN(n748) );
  XNOR2_X1 U447 ( .A(n502), .B(n499), .ZN(n383) );
  NAND2_X1 U448 ( .A1(n389), .A2(n361), .ZN(n386) );
  NAND2_X1 U449 ( .A1(n758), .A2(n366), .ZN(n389) );
  INV_X1 U450 ( .A(KEYINPUT34), .ZN(n557) );
  BUF_X1 U451 ( .A(n556), .Z(n623) );
  XNOR2_X1 U452 ( .A(n420), .B(n419), .ZN(n418) );
  XNOR2_X1 U453 ( .A(n442), .B(n754), .ZN(n421) );
  XNOR2_X1 U454 ( .A(n438), .B(n440), .ZN(n419) );
  XNOR2_X1 U455 ( .A(n377), .B(n375), .ZN(n667) );
  XNOR2_X1 U456 ( .A(n378), .B(n492), .ZN(n377) );
  XNOR2_X1 U457 ( .A(n493), .B(KEYINPUT9), .ZN(n376) );
  XNOR2_X1 U458 ( .A(n756), .B(n434), .ZN(n674) );
  NAND2_X1 U459 ( .A1(n414), .A2(n412), .ZN(n411) );
  AND2_X1 U460 ( .A1(n690), .A2(n413), .ZN(n412) );
  XNOR2_X1 U461 ( .A(n374), .B(n587), .ZN(n696) );
  AND2_X1 U462 ( .A1(n567), .A2(n356), .ZN(n540) );
  AND2_X1 U463 ( .A1(n702), .A2(n701), .ZN(n551) );
  AND2_X1 U464 ( .A1(n706), .A2(n702), .ZN(n356) );
  XNOR2_X1 U465 ( .A(n642), .B(n641), .ZN(n743) );
  INV_X1 U466 ( .A(n743), .ZN(n366) );
  XOR2_X1 U467 ( .A(n526), .B(KEYINPUT0), .Z(n357) );
  XOR2_X1 U468 ( .A(n651), .B(n650), .Z(n358) );
  XNOR2_X1 U469 ( .A(n657), .B(KEYINPUT59), .ZN(n359) );
  XNOR2_X1 U470 ( .A(KEYINPUT62), .B(n645), .ZN(n360) );
  XNOR2_X1 U471 ( .A(n421), .B(n418), .ZN(n663) );
  AND2_X1 U472 ( .A1(n513), .A2(KEYINPUT2), .ZN(n361) );
  XNOR2_X1 U473 ( .A(KEYINPUT15), .B(G902), .ZN(n644) );
  XOR2_X1 U474 ( .A(KEYINPUT120), .B(KEYINPUT60), .Z(n362) );
  XOR2_X1 U475 ( .A(n649), .B(KEYINPUT82), .Z(n363) );
  XNOR2_X1 U476 ( .A(n364), .B(n362), .ZN(G60) );
  NAND2_X1 U477 ( .A1(n659), .A2(n647), .ZN(n364) );
  XNOR2_X1 U478 ( .A(n365), .B(n363), .ZN(G57) );
  NAND2_X1 U479 ( .A1(n648), .A2(n647), .ZN(n365) );
  NAND2_X1 U480 ( .A1(n399), .A2(n397), .ZN(n396) );
  NOR2_X2 U481 ( .A1(n398), .A2(n391), .ZN(n758) );
  INV_X1 U482 ( .A(n389), .ZN(n700) );
  NAND2_X1 U483 ( .A1(n396), .A2(n392), .ZN(n391) );
  XNOR2_X1 U484 ( .A(n577), .B(n367), .ZN(n706) );
  XNOR2_X2 U485 ( .A(n436), .B(n435), .ZN(n577) );
  NOR2_X1 U486 ( .A1(n743), .A2(n644), .ZN(n390) );
  NAND2_X1 U487 ( .A1(n388), .A2(n390), .ZN(n387) );
  NAND2_X1 U488 ( .A1(n696), .A2(n695), .ZN(n370) );
  NAND2_X1 U489 ( .A1(n373), .A2(KEYINPUT47), .ZN(n372) );
  NAND2_X1 U490 ( .A1(n688), .A2(n721), .ZN(n373) );
  NAND2_X1 U491 ( .A1(n586), .A2(n585), .ZN(n374) );
  XNOR2_X1 U492 ( .A(n495), .B(n376), .ZN(n375) );
  NAND2_X1 U493 ( .A1(n494), .A2(G217), .ZN(n378) );
  INV_X1 U494 ( .A(n690), .ZN(n591) );
  NAND2_X1 U495 ( .A1(n384), .A2(n424), .ZN(n536) );
  AND2_X1 U496 ( .A1(n384), .A2(n473), .ZN(n520) );
  XNOR2_X1 U497 ( .A(n458), .B(KEYINPUT73), .ZN(n384) );
  XNOR2_X2 U498 ( .A(n385), .B(KEYINPUT66), .ZN(n662) );
  NOR2_X1 U499 ( .A1(n399), .A2(KEYINPUT79), .ZN(n398) );
  XNOR2_X2 U500 ( .A(n402), .B(n400), .ZN(n702) );
  NAND2_X1 U501 ( .A1(n663), .A2(n496), .ZN(n402) );
  NAND2_X1 U502 ( .A1(n644), .A2(G234), .ZN(n406) );
  NAND2_X1 U503 ( .A1(n758), .A2(n606), .ZN(n425) );
  XNOR2_X1 U504 ( .A(n462), .B(KEYINPUT5), .ZN(n407) );
  NAND2_X1 U505 ( .A1(n410), .A2(n409), .ZN(n408) );
  NAND2_X1 U506 ( .A1(n500), .A2(n461), .ZN(n409) );
  NAND2_X1 U507 ( .A1(n460), .A2(n459), .ZN(n410) );
  XNOR2_X1 U508 ( .A(n558), .B(n557), .ZN(n561) );
  INV_X1 U509 ( .A(n572), .ZN(n413) );
  INV_X1 U510 ( .A(n570), .ZN(n414) );
  NAND2_X1 U511 ( .A1(n591), .A2(n572), .ZN(n416) );
  NAND2_X1 U512 ( .A1(n570), .A2(n572), .ZN(n417) );
  NAND2_X1 U513 ( .A1(n660), .A2(n767), .ZN(n583) );
  XNOR2_X2 U514 ( .A(n505), .B(n422), .ZN(n754) );
  XNOR2_X2 U515 ( .A(n443), .B(G125), .ZN(n505) );
  AND2_X1 U516 ( .A1(n610), .A2(KEYINPUT44), .ZN(n426) );
  NOR2_X1 U517 ( .A1(n759), .A2(G952), .ZN(n677) );
  NAND2_X1 U518 ( .A1(n577), .A2(n551), .ZN(n624) );
  XNOR2_X1 U519 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U520 ( .A(n489), .B(n488), .ZN(n544) );
  INV_X1 U521 ( .A(n677), .ZN(n647) );
  XNOR2_X2 U522 ( .A(G143), .B(G128), .ZN(n507) );
  XNOR2_X2 U523 ( .A(n507), .B(n427), .ZN(n495) );
  XNOR2_X2 U524 ( .A(G110), .B(G107), .ZN(n501) );
  XNOR2_X1 U525 ( .A(n501), .B(n429), .ZN(n432) );
  NAND2_X1 U526 ( .A1(n759), .A2(G227), .ZN(n430) );
  XNOR2_X1 U527 ( .A(n430), .B(KEYINPUT75), .ZN(n431) );
  XNOR2_X1 U528 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X2 U529 ( .A(KEYINPUT4), .B(G101), .ZN(n504) );
  XNOR2_X1 U530 ( .A(n504), .B(G146), .ZN(n462) );
  XNOR2_X1 U531 ( .A(n433), .B(n462), .ZN(n434) );
  XNOR2_X1 U532 ( .A(KEYINPUT70), .B(G469), .ZN(n435) );
  INV_X1 U533 ( .A(n437), .ZN(n439) );
  XNOR2_X1 U534 ( .A(G128), .B(G119), .ZN(n438) );
  XOR2_X1 U535 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n441) );
  XNOR2_X1 U536 ( .A(G110), .B(KEYINPUT90), .ZN(n440) );
  NAND2_X1 U537 ( .A1(G221), .A2(n494), .ZN(n442) );
  INV_X1 U538 ( .A(G146), .ZN(n443) );
  NAND2_X1 U539 ( .A1(n447), .A2(G217), .ZN(n445) );
  XOR2_X1 U540 ( .A(KEYINPUT25), .B(KEYINPUT74), .Z(n444) );
  INV_X1 U541 ( .A(KEYINPUT91), .ZN(n446) );
  AND2_X1 U542 ( .A1(n447), .A2(G221), .ZN(n448) );
  XNOR2_X1 U543 ( .A(n448), .B(KEYINPUT21), .ZN(n701) );
  XNOR2_X1 U544 ( .A(n624), .B(KEYINPUT105), .ZN(n457) );
  XNOR2_X1 U545 ( .A(n449), .B(KEYINPUT14), .ZN(n453) );
  NAND2_X1 U546 ( .A1(G902), .A2(n453), .ZN(n450) );
  XNOR2_X1 U547 ( .A(KEYINPUT87), .B(n450), .ZN(n451) );
  NAND2_X1 U548 ( .A1(n451), .A2(G953), .ZN(n521) );
  XOR2_X1 U549 ( .A(KEYINPUT103), .B(n521), .Z(n452) );
  NOR2_X1 U550 ( .A1(n452), .A2(G900), .ZN(n455) );
  NAND2_X1 U551 ( .A1(n453), .A2(G952), .ZN(n454) );
  XNOR2_X1 U552 ( .A(n454), .B(KEYINPUT86), .ZN(n733) );
  NOR2_X1 U553 ( .A1(n733), .A2(G953), .ZN(n523) );
  NOR2_X1 U554 ( .A1(n455), .A2(n523), .ZN(n541) );
  INV_X1 U555 ( .A(n541), .ZN(n456) );
  NAND2_X1 U556 ( .A1(n457), .A2(n456), .ZN(n458) );
  INV_X1 U557 ( .A(n500), .ZN(n460) );
  NAND2_X1 U558 ( .A1(n474), .A2(G210), .ZN(n461) );
  INV_X1 U559 ( .A(n461), .ZN(n459) );
  XNOR2_X1 U560 ( .A(G137), .B(KEYINPUT94), .ZN(n463) );
  NAND2_X1 U561 ( .A1(n645), .A2(n496), .ZN(n469) );
  XNOR2_X1 U562 ( .A(KEYINPUT71), .B(KEYINPUT95), .ZN(n467) );
  INV_X1 U563 ( .A(G472), .ZN(n466) );
  XNOR2_X1 U564 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X2 U565 ( .A(n469), .B(n468), .ZN(n537) );
  NAND2_X1 U566 ( .A1(n496), .A2(n470), .ZN(n514) );
  AND2_X1 U567 ( .A1(n514), .A2(G214), .ZN(n546) );
  INV_X1 U568 ( .A(KEYINPUT30), .ZN(n471) );
  XNOR2_X1 U569 ( .A(n472), .B(n471), .ZN(n473) );
  NAND2_X1 U570 ( .A1(G214), .A2(n474), .ZN(n476) );
  XNOR2_X1 U571 ( .A(n476), .B(n475), .ZN(n480) );
  XNOR2_X1 U572 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U573 ( .A(n480), .B(n479), .Z(n484) );
  XNOR2_X1 U574 ( .A(n481), .B(G104), .ZN(n499) );
  XOR2_X1 U575 ( .A(n482), .B(n499), .Z(n483) );
  XNOR2_X1 U576 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U577 ( .A(n485), .B(n754), .ZN(n657) );
  NOR2_X1 U578 ( .A1(G902), .A2(n657), .ZN(n489) );
  XNOR2_X1 U579 ( .A(KEYINPUT13), .B(KEYINPUT98), .ZN(n487) );
  INV_X1 U580 ( .A(G475), .ZN(n486) );
  XNOR2_X1 U581 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U582 ( .A(KEYINPUT101), .B(G478), .Z(n497) );
  XNOR2_X1 U583 ( .A(n498), .B(n497), .ZN(n543) );
  INV_X1 U584 ( .A(n543), .ZN(n528) );
  OR2_X1 U585 ( .A1(n544), .A2(n528), .ZN(n559) );
  XNOR2_X1 U586 ( .A(n501), .B(KEYINPUT16), .ZN(n502) );
  XNOR2_X1 U587 ( .A(n504), .B(n503), .ZN(n506) );
  XNOR2_X1 U588 ( .A(n506), .B(n505), .ZN(n511) );
  NAND2_X1 U589 ( .A1(n759), .A2(G224), .ZN(n508) );
  XNOR2_X1 U590 ( .A(n508), .B(KEYINPUT76), .ZN(n509) );
  XNOR2_X1 U591 ( .A(n507), .B(n509), .ZN(n510) );
  XNOR2_X1 U592 ( .A(n510), .B(n511), .ZN(n512) );
  XNOR2_X1 U593 ( .A(n748), .B(n512), .ZN(n651) );
  INV_X1 U594 ( .A(n644), .ZN(n513) );
  NAND2_X1 U595 ( .A1(n514), .A2(G210), .ZN(n516) );
  INV_X1 U596 ( .A(KEYINPUT85), .ZN(n515) );
  XNOR2_X1 U597 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X2 U598 ( .A(n518), .B(n517), .ZN(n549) );
  NOR2_X1 U599 ( .A1(n559), .A2(n549), .ZN(n519) );
  NAND2_X1 U600 ( .A1(n520), .A2(n519), .ZN(n599) );
  XNOR2_X1 U601 ( .A(n599), .B(G143), .ZN(G45) );
  XNOR2_X2 U602 ( .A(n584), .B(KEYINPUT19), .ZN(n588) );
  NOR2_X1 U603 ( .A1(G898), .A2(n521), .ZN(n522) );
  OR2_X1 U604 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U605 ( .A(n524), .B(KEYINPUT88), .ZN(n525) );
  NAND2_X1 U606 ( .A1(n588), .A2(n525), .ZN(n527) );
  INV_X1 U607 ( .A(KEYINPUT83), .ZN(n526) );
  NAND2_X1 U608 ( .A1(n544), .A2(n528), .ZN(n720) );
  INV_X1 U609 ( .A(n701), .ZN(n529) );
  NOR2_X1 U610 ( .A1(n720), .A2(n529), .ZN(n530) );
  NAND2_X1 U611 ( .A1(n556), .A2(n530), .ZN(n532) );
  INV_X1 U612 ( .A(KEYINPUT22), .ZN(n531) );
  INV_X1 U613 ( .A(n702), .ZN(n565) );
  NAND2_X1 U614 ( .A1(n537), .A2(n565), .ZN(n533) );
  INV_X1 U615 ( .A(n706), .ZN(n695) );
  NOR2_X1 U616 ( .A1(n533), .A2(n695), .ZN(n534) );
  NAND2_X1 U617 ( .A1(n539), .A2(n534), .ZN(n634) );
  XNOR2_X1 U618 ( .A(n634), .B(G110), .ZN(G12) );
  INV_X1 U619 ( .A(KEYINPUT39), .ZN(n535) );
  XNOR2_X2 U620 ( .A(n536), .B(n535), .ZN(n570) );
  AND2_X1 U621 ( .A1(n544), .A2(n543), .ZN(n692) );
  INV_X1 U622 ( .A(n692), .ZN(n592) );
  OR2_X1 U623 ( .A1(n570), .A2(n592), .ZN(n605) );
  XNOR2_X1 U624 ( .A(n605), .B(G134), .ZN(G36) );
  XNOR2_X1 U625 ( .A(n537), .B(KEYINPUT6), .ZN(n553) );
  INV_X1 U626 ( .A(n553), .ZN(n538) );
  XNOR2_X1 U627 ( .A(n540), .B(KEYINPUT102), .ZN(n630) );
  XOR2_X1 U628 ( .A(G101), .B(n630), .Z(G3) );
  NOR2_X1 U629 ( .A1(n541), .A2(n702), .ZN(n542) );
  NAND2_X1 U630 ( .A1(n542), .A2(n701), .ZN(n575) );
  XNOR2_X1 U631 ( .A(n545), .B(KEYINPUT104), .ZN(n586) );
  INV_X1 U632 ( .A(n546), .ZN(n717) );
  AND2_X1 U633 ( .A1(n586), .A2(n717), .ZN(n547) );
  NAND2_X1 U634 ( .A1(n547), .A2(n706), .ZN(n548) );
  XNOR2_X1 U635 ( .A(n548), .B(KEYINPUT43), .ZN(n550) );
  NAND2_X1 U636 ( .A1(n550), .A2(n549), .ZN(n604) );
  XNOR2_X1 U637 ( .A(n604), .B(G140), .ZN(G42) );
  XNOR2_X1 U638 ( .A(G122), .B(KEYINPUT126), .ZN(n564) );
  INV_X1 U639 ( .A(n551), .ZN(n705) );
  INV_X1 U640 ( .A(n620), .ZN(n552) );
  NAND2_X1 U641 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U642 ( .A(KEYINPUT84), .B(KEYINPUT33), .ZN(n554) );
  NAND2_X1 U643 ( .A1(n727), .A2(n623), .ZN(n558) );
  INV_X1 U644 ( .A(n559), .ZN(n560) );
  NAND2_X1 U645 ( .A1(n561), .A2(n560), .ZN(n563) );
  XOR2_X1 U646 ( .A(KEYINPUT77), .B(KEYINPUT35), .Z(n562) );
  XOR2_X1 U647 ( .A(n564), .B(n612), .Z(G24) );
  XNOR2_X1 U648 ( .A(G119), .B(KEYINPUT127), .ZN(n569) );
  AND2_X1 U649 ( .A1(n695), .A2(n565), .ZN(n566) );
  NAND2_X1 U650 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X2 U651 ( .A(n568), .B(KEYINPUT32), .ZN(n607) );
  XOR2_X1 U652 ( .A(n569), .B(n607), .Z(G21) );
  INV_X1 U653 ( .A(KEYINPUT107), .ZN(n571) );
  XNOR2_X1 U654 ( .A(n571), .B(KEYINPUT40), .ZN(n572) );
  NAND2_X1 U655 ( .A1(n718), .A2(n717), .ZN(n722) );
  NOR2_X1 U656 ( .A1(n720), .A2(n722), .ZN(n574) );
  XNOR2_X1 U657 ( .A(KEYINPUT41), .B(KEYINPUT108), .ZN(n573) );
  XNOR2_X1 U658 ( .A(n574), .B(n573), .ZN(n735) );
  XNOR2_X1 U659 ( .A(KEYINPUT28), .B(n576), .ZN(n578) );
  NAND2_X1 U660 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U661 ( .A(n579), .B(KEYINPUT106), .ZN(n590) );
  NOR2_X1 U662 ( .A1(n735), .A2(n590), .ZN(n581) );
  INV_X1 U663 ( .A(KEYINPUT42), .ZN(n580) );
  XNOR2_X1 U664 ( .A(n581), .B(n580), .ZN(n767) );
  XNOR2_X1 U665 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n582) );
  XNOR2_X1 U666 ( .A(n583), .B(n582), .ZN(n602) );
  INV_X1 U667 ( .A(n584), .ZN(n585) );
  INV_X1 U668 ( .A(KEYINPUT36), .ZN(n587) );
  INV_X1 U669 ( .A(n588), .ZN(n589) );
  NOR2_X2 U670 ( .A1(n590), .A2(n589), .ZN(n688) );
  NAND2_X1 U671 ( .A1(n592), .A2(n591), .ZN(n721) );
  INV_X1 U672 ( .A(KEYINPUT47), .ZN(n593) );
  AND2_X1 U673 ( .A1(n593), .A2(KEYINPUT78), .ZN(n594) );
  NAND2_X1 U674 ( .A1(n721), .A2(n594), .ZN(n596) );
  OR2_X1 U675 ( .A1(KEYINPUT78), .A2(n721), .ZN(n595) );
  NAND2_X1 U676 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U677 ( .A1(n688), .A2(n597), .ZN(n598) );
  NAND2_X1 U678 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X2 U679 ( .A1(n602), .A2(n601), .ZN(n603) );
  INV_X1 U680 ( .A(KEYINPUT2), .ZN(n643) );
  AND2_X1 U681 ( .A1(n643), .A2(KEYINPUT72), .ZN(n606) );
  NOR2_X1 U682 ( .A1(n613), .A2(KEYINPUT67), .ZN(n608) );
  INV_X1 U683 ( .A(n608), .ZN(n611) );
  INV_X1 U684 ( .A(KEYINPUT81), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n612), .A2(n609), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n611), .A2(n426), .ZN(n618) );
  INV_X1 U687 ( .A(n612), .ZN(n619) );
  NAND2_X1 U688 ( .A1(n619), .A2(n613), .ZN(n616) );
  OR2_X1 U689 ( .A1(KEYINPUT81), .A2(KEYINPUT67), .ZN(n614) );
  NOR2_X1 U690 ( .A1(n614), .A2(KEYINPUT44), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n640) );
  NAND2_X1 U693 ( .A1(n619), .A2(KEYINPUT81), .ZN(n633) );
  NOR2_X1 U694 ( .A1(n620), .A2(n537), .ZN(n621) );
  XNOR2_X1 U695 ( .A(n621), .B(KEYINPUT96), .ZN(n713) );
  NAND2_X1 U696 ( .A1(n713), .A2(n623), .ZN(n622) );
  XNOR2_X1 U697 ( .A(n622), .B(KEYINPUT31), .ZN(n693) );
  INV_X1 U698 ( .A(n623), .ZN(n627) );
  INV_X1 U699 ( .A(n624), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n537), .A2(n625), .ZN(n626) );
  NOR2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n683) );
  NOR2_X1 U702 ( .A1(n693), .A2(n683), .ZN(n629) );
  XOR2_X1 U703 ( .A(KEYINPUT78), .B(n721), .Z(n628) );
  NOR2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n631) );
  NOR2_X1 U705 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U706 ( .A1(n633), .A2(n632), .ZN(n638) );
  INV_X1 U707 ( .A(n607), .ZN(n636) );
  NAND2_X1 U708 ( .A1(n634), .A2(KEYINPUT67), .ZN(n635) );
  NOR2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n642) );
  XNOR2_X1 U711 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n641) );
  NAND2_X1 U712 ( .A1(n662), .A2(G472), .ZN(n646) );
  XNOR2_X1 U713 ( .A(n646), .B(n360), .ZN(n648) );
  XNOR2_X1 U714 ( .A(KEYINPUT109), .B(KEYINPUT63), .ZN(n649) );
  NAND2_X1 U715 ( .A1(n662), .A2(G210), .ZN(n652) );
  XOR2_X1 U716 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n650) );
  XNOR2_X1 U717 ( .A(n652), .B(n358), .ZN(n653) );
  AND2_X2 U718 ( .A1(n653), .A2(n647), .ZN(n656) );
  XNOR2_X1 U719 ( .A(KEYINPUT118), .B(KEYINPUT56), .ZN(n654) );
  XNOR2_X1 U720 ( .A(n654), .B(KEYINPUT80), .ZN(n655) );
  XNOR2_X1 U721 ( .A(n656), .B(n655), .ZN(G51) );
  NAND2_X1 U722 ( .A1(n662), .A2(G475), .ZN(n658) );
  XNOR2_X1 U723 ( .A(n658), .B(n359), .ZN(n659) );
  BUF_X1 U724 ( .A(n660), .Z(n661) );
  XNOR2_X1 U725 ( .A(n661), .B(G131), .ZN(G33) );
  BUF_X1 U726 ( .A(n662), .Z(n671) );
  NAND2_X1 U727 ( .A1(n671), .A2(G217), .ZN(n665) );
  XOR2_X1 U728 ( .A(n663), .B(KEYINPUT122), .Z(n664) );
  XNOR2_X1 U729 ( .A(n665), .B(n664), .ZN(n666) );
  NOR2_X1 U730 ( .A1(n666), .A2(n677), .ZN(G66) );
  NAND2_X1 U731 ( .A1(n671), .A2(G478), .ZN(n669) );
  XNOR2_X1 U732 ( .A(n667), .B(KEYINPUT121), .ZN(n668) );
  XNOR2_X1 U733 ( .A(n669), .B(n668), .ZN(n670) );
  NOR2_X1 U734 ( .A1(n670), .A2(n677), .ZN(G63) );
  NAND2_X1 U735 ( .A1(n671), .A2(G469), .ZN(n676) );
  XNOR2_X1 U736 ( .A(KEYINPUT119), .B(KEYINPUT57), .ZN(n672) );
  XNOR2_X1 U737 ( .A(n672), .B(KEYINPUT58), .ZN(n673) );
  XNOR2_X1 U738 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U739 ( .A(n676), .B(n675), .ZN(n678) );
  NOR2_X1 U740 ( .A1(n678), .A2(n677), .ZN(G54) );
  NAND2_X1 U741 ( .A1(n683), .A2(n690), .ZN(n679) );
  XNOR2_X1 U742 ( .A(n679), .B(G104), .ZN(G6) );
  XOR2_X1 U743 ( .A(KEYINPUT27), .B(KEYINPUT111), .Z(n681) );
  XNOR2_X1 U744 ( .A(G107), .B(KEYINPUT26), .ZN(n680) );
  XNOR2_X1 U745 ( .A(n681), .B(n680), .ZN(n682) );
  XOR2_X1 U746 ( .A(KEYINPUT110), .B(n682), .Z(n685) );
  NAND2_X1 U747 ( .A1(n683), .A2(n692), .ZN(n684) );
  XNOR2_X1 U748 ( .A(n685), .B(n684), .ZN(G9) );
  XOR2_X1 U749 ( .A(G128), .B(KEYINPUT29), .Z(n687) );
  NAND2_X1 U750 ( .A1(n688), .A2(n692), .ZN(n686) );
  XNOR2_X1 U751 ( .A(n687), .B(n686), .ZN(G30) );
  NAND2_X1 U752 ( .A1(n688), .A2(n690), .ZN(n689) );
  XNOR2_X1 U753 ( .A(n689), .B(G146), .ZN(G48) );
  NAND2_X1 U754 ( .A1(n693), .A2(n690), .ZN(n691) );
  XNOR2_X1 U755 ( .A(n691), .B(G113), .ZN(G15) );
  NAND2_X1 U756 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U757 ( .A(n694), .B(G116), .ZN(G18) );
  NAND2_X1 U758 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U759 ( .A(KEYINPUT37), .B(n697), .Z(n698) );
  XNOR2_X1 U760 ( .A(n698), .B(KEYINPUT112), .ZN(n699) );
  XNOR2_X1 U761 ( .A(G125), .B(n699), .ZN(G27) );
  XNOR2_X1 U762 ( .A(n700), .B(KEYINPUT2), .ZN(n740) );
  NOR2_X1 U763 ( .A1(n702), .A2(n701), .ZN(n704) );
  XNOR2_X1 U764 ( .A(KEYINPUT113), .B(KEYINPUT49), .ZN(n703) );
  XNOR2_X1 U765 ( .A(n704), .B(n703), .ZN(n710) );
  NAND2_X1 U766 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U767 ( .A(n707), .B(KEYINPUT50), .ZN(n708) );
  NAND2_X1 U768 ( .A1(n708), .A2(n537), .ZN(n709) );
  NOR2_X1 U769 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U770 ( .A(n711), .B(KEYINPUT114), .ZN(n712) );
  NOR2_X1 U771 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U772 ( .A(n714), .B(KEYINPUT51), .ZN(n715) );
  XNOR2_X1 U773 ( .A(KEYINPUT115), .B(n715), .ZN(n716) );
  NOR2_X1 U774 ( .A1(n735), .A2(n716), .ZN(n730) );
  NOR2_X1 U775 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U776 ( .A1(n720), .A2(n719), .ZN(n726) );
  INV_X1 U777 ( .A(n721), .ZN(n723) );
  NOR2_X1 U778 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U779 ( .A(n724), .B(KEYINPUT116), .ZN(n725) );
  NOR2_X1 U780 ( .A1(n726), .A2(n725), .ZN(n728) );
  INV_X1 U781 ( .A(n727), .ZN(n734) );
  NOR2_X1 U782 ( .A1(n728), .A2(n734), .ZN(n729) );
  NOR2_X1 U783 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U784 ( .A(n731), .B(KEYINPUT52), .ZN(n732) );
  NOR2_X1 U785 ( .A1(n733), .A2(n732), .ZN(n737) );
  NOR2_X1 U786 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U787 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U788 ( .A(KEYINPUT117), .B(n738), .Z(n739) );
  NAND2_X1 U789 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U790 ( .A1(n741), .A2(G953), .ZN(n742) );
  XNOR2_X1 U791 ( .A(n742), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U792 ( .A1(n366), .A2(n759), .ZN(n747) );
  NAND2_X1 U793 ( .A1(G953), .A2(G224), .ZN(n744) );
  XNOR2_X1 U794 ( .A(KEYINPUT61), .B(n744), .ZN(n745) );
  NAND2_X1 U795 ( .A1(n745), .A2(G898), .ZN(n746) );
  NAND2_X1 U796 ( .A1(n747), .A2(n746), .ZN(n752) );
  XOR2_X1 U797 ( .A(n748), .B(G101), .Z(n750) );
  NOR2_X1 U798 ( .A1(n759), .A2(G898), .ZN(n749) );
  NOR2_X1 U799 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U800 ( .A(n752), .B(n751), .ZN(n753) );
  XOR2_X1 U801 ( .A(KEYINPUT123), .B(n753), .Z(G69) );
  XNOR2_X1 U802 ( .A(KEYINPUT124), .B(n754), .ZN(n755) );
  XNOR2_X1 U803 ( .A(n755), .B(KEYINPUT4), .ZN(n757) );
  XNOR2_X1 U804 ( .A(n756), .B(n757), .ZN(n761) );
  XOR2_X1 U805 ( .A(n761), .B(n758), .Z(n760) );
  NAND2_X1 U806 ( .A1(n760), .A2(n759), .ZN(n765) );
  XNOR2_X1 U807 ( .A(G227), .B(n761), .ZN(n762) );
  NAND2_X1 U808 ( .A1(n762), .A2(G900), .ZN(n763) );
  NAND2_X1 U809 ( .A1(n763), .A2(G953), .ZN(n764) );
  NAND2_X1 U810 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U811 ( .A(KEYINPUT125), .B(n766), .Z(G72) );
  XNOR2_X1 U812 ( .A(n767), .B(G137), .ZN(G39) );
endmodule

