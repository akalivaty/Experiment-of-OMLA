//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940;
  INV_X1    g000(.A(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G217), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT71), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G128), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n192), .B(new_n194), .C1(G119), .C2(new_n193), .ZN(new_n195));
  XNOR2_X1  g009(.A(G119), .B(G128), .ZN(new_n196));
  XOR2_X1   g010(.A(KEYINPUT24), .B(G110), .Z(new_n197));
  OAI22_X1  g011(.A1(new_n195), .A2(G110), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT16), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G125), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G140), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OAI211_X1 g019(.A(G146), .B(new_n201), .C1(new_n205), .C2(new_n199), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(KEYINPUT74), .ZN(new_n207));
  XNOR2_X1  g021(.A(G125), .B(G140), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT74), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n198), .A2(new_n206), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(KEYINPUT16), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n201), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(new_n211), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n206), .A2(KEYINPUT73), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT73), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n214), .A2(new_n218), .A3(G146), .A4(new_n201), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n197), .A2(new_n196), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n195), .A2(KEYINPUT72), .A3(G110), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT72), .B1(new_n195), .B2(G110), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n213), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT22), .B(G137), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n226), .B(KEYINPUT75), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT68), .B(G953), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(G221), .A3(G234), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n227), .B(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n230), .B(new_n213), .C1(new_n224), .C2(new_n220), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G902), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(KEYINPUT25), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT25), .B1(new_n234), .B2(new_n235), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n189), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n189), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n235), .ZN(new_n241));
  XOR2_X1   g055(.A(new_n241), .B(KEYINPUT76), .Z(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n234), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n239), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G472), .ZN(new_n246));
  INV_X1    g060(.A(G116), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(G119), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT66), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(new_n247), .B2(G119), .ZN(new_n251));
  NOR3_X1   g065(.A1(new_n191), .A2(KEYINPUT66), .A3(G116), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n249), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT2), .B(G113), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT66), .B1(new_n191), .B2(G116), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n250), .A2(new_n247), .A3(G119), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n248), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n254), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n211), .A2(G143), .ZN(new_n262));
  INV_X1    g076(.A(G143), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G146), .ZN(new_n264));
  AND2_X1   g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G143), .B(G146), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT0), .B(G128), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G137), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(G134), .ZN(new_n272));
  INV_X1    g086(.A(G134), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT11), .B1(new_n273), .B2(G137), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT11), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n271), .A3(G134), .ZN(new_n276));
  AOI211_X1 g090(.A(G131), .B(new_n272), .C1(new_n274), .C2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G131), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n274), .A2(new_n276), .ZN(new_n279));
  INV_X1    g093(.A(new_n272), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n270), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n278), .A3(new_n280), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT65), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n284), .B1(new_n271), .B2(G134), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n271), .A2(G134), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n273), .A2(KEYINPUT65), .A3(G137), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G131), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n262), .B(new_n264), .C1(KEYINPUT1), .C2(new_n193), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT1), .B1(new_n263), .B2(G146), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n263), .A2(G146), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n211), .A2(G143), .ZN(new_n293));
  OAI211_X1 g107(.A(G128), .B(new_n291), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n283), .A2(new_n289), .A3(new_n290), .A4(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n282), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT30), .B1(new_n296), .B2(KEYINPUT64), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT64), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT30), .ZN(new_n299));
  AOI211_X1 g113(.A(new_n298), .B(new_n299), .C1(new_n282), .C2(new_n295), .ZN(new_n300));
  OAI211_X1 g114(.A(KEYINPUT67), .B(new_n261), .C1(new_n297), .C2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n261), .ZN(new_n302));
  AND4_X1   g116(.A1(new_n283), .A2(new_n289), .A3(new_n290), .A4(new_n294), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n275), .B1(G134), .B2(new_n271), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n273), .A2(KEYINPUT11), .A3(G137), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n280), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G131), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n269), .B1(new_n307), .B2(new_n283), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT64), .B1(new_n303), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n299), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n296), .A2(KEYINPUT64), .A3(KEYINPUT30), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n302), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n302), .A2(new_n282), .A3(new_n295), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT67), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n301), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT31), .ZN(new_n317));
  INV_X1    g131(.A(G237), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n228), .A2(G210), .A3(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(KEYINPUT70), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT26), .B(G101), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n320), .B(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n316), .A2(new_n317), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n324), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n296), .B(new_n302), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT28), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n313), .A2(new_n328), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n326), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n317), .B1(new_n316), .B2(new_n324), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n246), .B(new_n235), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT32), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n316), .A2(new_n324), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT31), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(new_n331), .A3(new_n325), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT32), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n338), .A2(new_n339), .A3(new_n246), .A4(new_n235), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n316), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n326), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n344));
  OR3_X1    g158(.A1(new_n329), .A2(new_n326), .A3(new_n330), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n346), .B(new_n235), .C1(new_n344), .C2(new_n345), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G472), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n245), .B1(new_n341), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(G214), .B1(G237), .B2(G902), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n269), .A2(G125), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n294), .A2(new_n290), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n351), .B1(new_n352), .B2(G125), .ZN(new_n353));
  INV_X1    g167(.A(G224), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(G953), .ZN(new_n355));
  XOR2_X1   g169(.A(new_n353), .B(new_n355), .Z(new_n356));
  XNOR2_X1  g170(.A(G110), .B(G122), .ZN(new_n357));
  INV_X1    g171(.A(G104), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT3), .B1(new_n358), .B2(G107), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n360));
  INV_X1    g174(.A(G107), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n361), .A3(G104), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(G107), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n359), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G101), .ZN(new_n365));
  INV_X1    g179(.A(G101), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n359), .A2(new_n362), .A3(new_n366), .A4(new_n363), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(KEYINPUT4), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n364), .A2(new_n369), .A3(G101), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n261), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(KEYINPUT5), .B(new_n249), .C1(new_n251), .C2(new_n252), .ZN(new_n372));
  INV_X1    g186(.A(G113), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT5), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n373), .B1(new_n248), .B2(new_n374), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n372), .A2(new_n375), .B1(new_n258), .B2(new_n259), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n358), .A2(G107), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n361), .A2(G104), .ZN(new_n378));
  OAI21_X1  g192(.A(G101), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n367), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT78), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT78), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n367), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n376), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n371), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT82), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n357), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n371), .A2(new_n384), .A3(KEYINPUT82), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n371), .A2(new_n384), .A3(new_n357), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT6), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n387), .A2(KEYINPUT6), .A3(new_n388), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n356), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(G210), .B1(G237), .B2(G902), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT7), .B1(new_n354), .B2(G953), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n353), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n353), .A2(new_n397), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n390), .A3(new_n399), .ZN(new_n400));
  XOR2_X1   g214(.A(new_n357), .B(KEYINPUT8), .Z(new_n401));
  INV_X1    g215(.A(new_n380), .ZN(new_n402));
  OR2_X1    g216(.A1(new_n376), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n401), .B1(new_n403), .B2(new_n384), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n235), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n394), .A2(new_n396), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n356), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n387), .A2(KEYINPUT6), .A3(new_n388), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n387), .A2(new_n388), .B1(KEYINPUT6), .B2(new_n390), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n405), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n395), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n350), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT83), .ZN(new_n414));
  INV_X1    g228(.A(new_n350), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n396), .B1(new_n394), .B2(new_n405), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n410), .A2(new_n395), .A3(new_n411), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT83), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n414), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n422));
  INV_X1    g236(.A(G953), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT68), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT68), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G953), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n424), .A2(new_n426), .A3(G214), .A4(new_n318), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n263), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n228), .A2(G143), .A3(G214), .A4(new_n318), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G131), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT17), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n428), .A2(new_n429), .A3(new_n278), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AND4_X1   g248(.A1(KEYINPUT85), .A2(new_n430), .A3(KEYINPUT17), .A4(G131), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n278), .B1(new_n428), .B2(new_n429), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT85), .B1(new_n436), .B2(KEYINPUT17), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n220), .B(new_n434), .C1(new_n435), .C2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G113), .B(G122), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(new_n358), .ZN(new_n440));
  OR3_X1    g254(.A1(new_n208), .A2(KEYINPUT84), .A3(new_n211), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT84), .B1(new_n208), .B2(new_n211), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n212), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AND2_X1   g257(.A1(KEYINPUT18), .A2(G131), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n428), .A2(new_n429), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n444), .B1(new_n428), .B2(new_n429), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n438), .A2(new_n440), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT19), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n207), .A2(new_n210), .A3(new_n449), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n450), .B(new_n211), .C1(new_n449), .C2(new_n208), .ZN(new_n451));
  INV_X1    g265(.A(new_n433), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n451), .B(new_n206), .C1(new_n436), .C2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n447), .ZN(new_n454));
  INV_X1    g268(.A(new_n440), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n448), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(G475), .A2(G902), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(KEYINPUT86), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n422), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  AOI211_X1 g275(.A(KEYINPUT20), .B(new_n459), .C1(new_n448), .C2(new_n456), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n438), .A2(new_n447), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n455), .ZN(new_n464));
  AOI21_X1  g278(.A(G902), .B1(new_n464), .B2(new_n448), .ZN(new_n465));
  INV_X1    g279(.A(G475), .ZN(new_n466));
  OAI22_X1  g280(.A1(new_n461), .A2(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G952), .ZN(new_n468));
  AOI211_X1 g282(.A(G953), .B(new_n468), .C1(G234), .C2(G237), .ZN(new_n469));
  AOI211_X1 g283(.A(new_n235), .B(new_n228), .C1(G234), .C2(G237), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(G898), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT9), .B(G234), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(G217), .A3(new_n423), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT13), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n193), .B2(G143), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n263), .A2(KEYINPUT13), .A3(G128), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n193), .A2(G143), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G134), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n263), .A2(G128), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n479), .A3(new_n273), .ZN(new_n484));
  INV_X1    g298(.A(G122), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G116), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n247), .A2(G122), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n486), .A2(new_n487), .A3(new_n361), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n361), .B1(new_n486), .B2(new_n487), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n484), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(G116), .B(G122), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n361), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n483), .A2(new_n479), .A3(new_n273), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n273), .B1(new_n483), .B2(new_n479), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n247), .A2(KEYINPUT14), .A3(G122), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G107), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT14), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n497), .B1(new_n498), .B2(new_n491), .ZN(new_n499));
  OAI22_X1  g313(.A1(new_n482), .A2(new_n490), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n475), .B1(new_n500), .B2(KEYINPUT87), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(KEYINPUT87), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT87), .ZN(new_n504));
  OAI221_X1 g318(.A(new_n504), .B1(new_n495), .B2(new_n499), .C1(new_n482), .C2(new_n490), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n475), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n235), .ZN(new_n509));
  INV_X1    g323(.A(G478), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(KEYINPUT15), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n508), .B(new_n235), .C1(KEYINPUT15), .C2(new_n510), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n467), .A2(new_n472), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(G221), .B1(new_n473), .B2(G902), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n277), .A2(new_n281), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n352), .B1(new_n381), .B2(new_n383), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n294), .A2(new_n290), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(new_n380), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n518), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT12), .B1(new_n518), .B2(KEYINPUT79), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI221_X1 g338(.A(new_n518), .B1(KEYINPUT79), .B2(KEYINPUT12), .C1(new_n519), .C2(new_n521), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n381), .A2(new_n352), .A3(KEYINPUT10), .A4(new_n383), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n368), .A2(new_n270), .A3(new_n370), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT77), .B(KEYINPUT10), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n529), .B1(new_n520), .B2(new_n380), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n527), .A2(new_n528), .A3(new_n517), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n228), .A2(G227), .ZN(new_n532));
  XOR2_X1   g346(.A(G110), .B(G140), .Z(new_n533));
  XOR2_X1   g347(.A(new_n532), .B(new_n533), .Z(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT80), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT80), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n531), .A2(new_n537), .A3(new_n534), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n526), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n518), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n531), .ZN(new_n542));
  INV_X1    g356(.A(new_n534), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G469), .ZN(new_n546));
  AND4_X1   g360(.A1(KEYINPUT81), .A2(new_n545), .A3(new_n546), .A4(new_n235), .ZN(new_n547));
  AOI21_X1  g361(.A(G902), .B1(new_n539), .B2(new_n544), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT81), .B1(new_n548), .B2(new_n546), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n541), .A2(new_n531), .A3(new_n534), .ZN(new_n551));
  AND4_X1   g365(.A1(new_n517), .A2(new_n527), .A3(new_n528), .A4(new_n530), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n524), .B2(new_n525), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n551), .B1(new_n553), .B2(new_n534), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n546), .B1(new_n554), .B2(new_n235), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n515), .B(new_n516), .C1(new_n550), .C2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n421), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n349), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(G101), .ZN(G3));
  INV_X1    g373(.A(KEYINPUT90), .ZN(new_n560));
  INV_X1    g374(.A(new_n472), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n418), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT33), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n507), .B1(new_n503), .B2(new_n505), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n563), .B1(new_n564), .B2(new_n501), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n500), .A2(KEYINPUT88), .A3(new_n507), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n507), .B1(new_n500), .B2(KEYINPUT88), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT33), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n510), .A2(G902), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n565), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT89), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n509), .A2(new_n510), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT89), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n565), .A2(new_n573), .A3(new_n568), .A4(new_n569), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n467), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n560), .B1(new_n562), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n576), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n578), .A2(new_n418), .A3(KEYINPUT90), .A4(new_n561), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n235), .B1(new_n332), .B2(new_n333), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G472), .ZN(new_n582));
  INV_X1    g396(.A(new_n245), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n334), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n516), .B1(new_n550), .B2(new_n555), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT34), .B(G104), .Z(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(G6));
  INV_X1    g403(.A(new_n448), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n440), .B1(new_n438), .B2(new_n447), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n235), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G475), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n514), .B(new_n593), .C1(new_n461), .C2(new_n462), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n562), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n586), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT35), .B(G107), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G9));
  NOR2_X1   g412(.A1(new_n230), .A2(KEYINPUT36), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(new_n225), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n242), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n239), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n582), .A2(new_n334), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT91), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT91), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n582), .A2(new_n605), .A3(new_n334), .A4(new_n602), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n557), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT37), .B(G110), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G12));
  INV_X1    g423(.A(new_n516), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n545), .A2(new_n546), .A3(new_n235), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT81), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n548), .A2(KEYINPUT81), .A3(new_n546), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n554), .A2(new_n235), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(G469), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n610), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n418), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n341), .A2(new_n348), .ZN(new_n621));
  INV_X1    g435(.A(new_n594), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT92), .B(G900), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n470), .A2(new_n623), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n624), .A2(new_n469), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n620), .A2(new_n621), .A3(new_n602), .A4(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G128), .ZN(G30));
  XNOR2_X1  g442(.A(new_n625), .B(KEYINPUT39), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n618), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n630), .B(KEYINPUT40), .Z(new_n631));
  OR2_X1    g445(.A1(new_n631), .A2(KEYINPUT95), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(KEYINPUT95), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n342), .A2(new_n324), .ZN(new_n634));
  AOI21_X1  g448(.A(G902), .B1(new_n327), .B2(new_n326), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n246), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n335), .B2(new_n340), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n416), .A2(new_n417), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT93), .B(KEYINPUT38), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT94), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n638), .B(new_n640), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n512), .A2(new_n513), .ZN(new_n642));
  OR2_X1    g456(.A1(new_n461), .A2(new_n462), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n642), .B1(new_n643), .B2(new_n593), .ZN(new_n644));
  INV_X1    g458(.A(new_n602), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n645), .A3(new_n350), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n637), .A2(new_n641), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n632), .A2(new_n633), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G143), .ZN(G45));
  NAND3_X1  g463(.A1(new_n467), .A2(new_n575), .A3(new_n625), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n620), .A2(new_n621), .A3(new_n602), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G146), .ZN(G48));
  INV_X1    g467(.A(new_n548), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(G469), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n516), .B(new_n655), .C1(new_n547), .C2(new_n549), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT96), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n349), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n580), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT41), .B(G113), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G15));
  AND2_X1   g475(.A1(new_n658), .A2(new_n595), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(new_n247), .ZN(G18));
  INV_X1    g477(.A(KEYINPUT97), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n664), .B1(new_n656), .B2(new_n413), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n613), .A2(new_n614), .B1(G469), .B2(new_n654), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n666), .A2(KEYINPUT97), .A3(new_n418), .A4(new_n516), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n668), .A2(new_n621), .A3(new_n515), .A4(new_n602), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT98), .B(G119), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G21));
  INV_X1    g485(.A(KEYINPUT99), .ZN(new_n672));
  AOI22_X1  g486(.A1(new_n582), .A2(new_n334), .B1(new_n672), .B2(new_n581), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n581), .A2(new_n672), .A3(new_n246), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n644), .A2(new_n418), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n677), .A2(new_n561), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n676), .A2(new_n657), .A3(new_n678), .A4(new_n583), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT100), .B(G122), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G24));
  INV_X1    g495(.A(new_n668), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n581), .A2(new_n672), .ZN(new_n683));
  INV_X1    g497(.A(new_n334), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n246), .B1(new_n338), .B2(new_n235), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n650), .B(KEYINPUT101), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n686), .A2(new_n687), .A3(new_n602), .A4(new_n674), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n203), .ZN(G27));
  NAND3_X1  g504(.A1(new_n416), .A2(new_n417), .A3(new_n350), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n546), .A2(KEYINPUT102), .A3(G902), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n551), .B(new_n692), .C1(new_n553), .C2(new_n534), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n617), .B2(KEYINPUT102), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n516), .B1(new_n550), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n691), .B1(new_n696), .B2(KEYINPUT103), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT102), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n693), .B1(new_n555), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n610), .B1(new_n615), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n349), .A2(new_n697), .A3(new_n687), .A4(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT42), .B1(new_n703), .B2(KEYINPUT104), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n696), .A2(KEYINPUT103), .ZN(new_n705));
  INV_X1    g519(.A(new_n691), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n702), .A3(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n708), .A2(new_n709), .A3(new_n349), .A4(new_n687), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n704), .A2(KEYINPUT105), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT42), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n712), .B1(new_n703), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n710), .B2(new_n704), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G131), .ZN(G33));
  AND4_X1   g531(.A1(new_n349), .A2(new_n697), .A3(new_n626), .A4(new_n702), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT106), .B(G134), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G36));
  INV_X1    g534(.A(new_n575), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n467), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI22_X1  g538(.A1(new_n724), .A2(KEYINPUT108), .B1(KEYINPUT43), .B2(new_n722), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(KEYINPUT108), .B2(new_n724), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n726), .A2(KEYINPUT109), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(KEYINPUT109), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n645), .B1(new_n582), .B2(new_n334), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n554), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n546), .B1(new_n554), .B2(new_n734), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n546), .A2(new_n235), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n550), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(new_n740), .B2(new_n739), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n742), .A2(new_n516), .A3(new_n629), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n732), .A2(new_n706), .A3(new_n733), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G137), .ZN(G39));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n516), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT47), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n335), .A2(new_n340), .B1(new_n347), .B2(G472), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(new_n245), .A3(new_n651), .A4(new_n706), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G140), .ZN(G42));
  NOR3_X1   g565(.A1(new_n245), .A2(new_n415), .A3(new_n610), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT110), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n753), .A2(new_n641), .A3(new_n722), .ZN(new_n754));
  INV_X1    g568(.A(new_n666), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT49), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n755), .A2(KEYINPUT49), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n754), .A2(new_n637), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n637), .ZN(new_n759));
  INV_X1    g573(.A(new_n656), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n469), .A3(new_n706), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n759), .A2(new_n761), .A3(new_n245), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n578), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(G952), .A3(new_n423), .ZN(new_n764));
  INV_X1    g578(.A(new_n761), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n726), .A2(new_n349), .A3(new_n765), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(KEYINPUT48), .Z(new_n767));
  AND4_X1   g581(.A1(new_n583), .A2(new_n726), .A3(new_n469), .A4(new_n676), .ZN(new_n768));
  AOI211_X1 g582(.A(new_n764), .B(new_n767), .C1(new_n668), .C2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n350), .B1(KEYINPUT114), .B2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n768), .A2(new_n641), .A3(new_n760), .A4(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n770), .A2(KEYINPUT114), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n772), .B(new_n773), .Z(new_n774));
  NAND4_X1  g588(.A1(new_n762), .A2(new_n593), .A3(new_n643), .A4(new_n721), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n726), .A2(new_n765), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n673), .A2(new_n645), .A3(new_n675), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n775), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n747), .B1(new_n516), .B2(new_n755), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n706), .A3(new_n768), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n774), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n779), .B(KEYINPUT115), .Z(new_n784));
  NAND2_X1  g598(.A1(new_n774), .A2(new_n784), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT116), .Z(new_n786));
  NAND2_X1  g600(.A1(new_n782), .A2(KEYINPUT51), .ZN(new_n787));
  OAI221_X1 g601(.A(new_n769), .B1(KEYINPUT51), .B2(new_n783), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n349), .B(new_n657), .C1(new_n580), .C2(new_n595), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n790), .A2(new_n679), .A3(new_n669), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n643), .A2(new_n642), .A3(new_n593), .A4(new_n625), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n691), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n621), .A2(new_n618), .A3(new_n602), .A4(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(new_n688), .B2(new_n707), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n718), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n472), .B1(new_n576), .B2(new_n594), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n414), .A2(new_n797), .A3(new_n420), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n586), .A2(new_n798), .ZN(new_n799));
  AND4_X1   g613(.A1(KEYINPUT111), .A2(new_n607), .A3(new_n558), .A4(new_n799), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n349), .A2(new_n557), .B1(new_n586), .B2(new_n798), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT111), .B1(new_n801), .B2(new_n607), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n791), .B(new_n796), .C1(new_n800), .C2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n688), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n748), .A2(new_n619), .A3(new_n645), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n668), .A2(new_n805), .B1(new_n806), .B2(new_n626), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT113), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n239), .A2(new_n601), .A3(new_n625), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT112), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT112), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n239), .A2(new_n813), .A3(new_n601), .A4(new_n625), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n677), .A2(new_n700), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n810), .B1(new_n815), .B2(new_n637), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n812), .A2(new_n644), .A3(new_n418), .A4(new_n814), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n696), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n759), .A2(new_n818), .A3(KEYINPUT113), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n807), .A2(KEYINPUT52), .A3(new_n652), .A4(new_n820), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n627), .B(new_n652), .C1(new_n682), .C2(new_n688), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n816), .A2(new_n819), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n808), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n716), .A2(new_n804), .A3(new_n809), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n716), .A2(new_n804), .A3(KEYINPUT53), .A4(new_n825), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n789), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n826), .A2(KEYINPUT53), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n716), .A2(new_n804), .A3(new_n827), .A4(new_n825), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT54), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n788), .A2(new_n830), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(G952), .A2(G953), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n758), .B1(new_n834), .B2(new_n835), .ZN(G75));
  AND2_X1   g650(.A1(new_n831), .A2(new_n832), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(G210), .A3(G902), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n392), .A2(new_n356), .A3(new_n393), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n840), .A2(new_n410), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT55), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n838), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n842), .B1(new_n838), .B2(new_n839), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n228), .A2(G952), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(G51));
  INV_X1    g660(.A(new_n845), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n738), .B(KEYINPUT57), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n831), .A2(KEYINPUT54), .A3(new_n832), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n849), .B2(new_n833), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n851), .A3(new_n545), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n837), .A2(G902), .A3(new_n737), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n851), .B1(new_n850), .B2(new_n545), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n847), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT118), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI211_X1 g672(.A(KEYINPUT118), .B(new_n847), .C1(new_n854), .C2(new_n855), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(G54));
  NAND4_X1  g674(.A1(new_n837), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n861));
  INV_X1    g675(.A(new_n457), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n863), .A2(new_n864), .A3(new_n845), .ZN(G60));
  NAND2_X1  g679(.A1(G478), .A2(G902), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(KEYINPUT59), .Z(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n868), .B1(new_n830), .B2(new_n833), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n565), .A2(new_n568), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n869), .A2(KEYINPUT119), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n849), .A2(new_n833), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n872), .A2(new_n870), .A3(new_n867), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT119), .B1(new_n869), .B2(new_n870), .ZN(new_n874));
  NOR4_X1   g688(.A1(new_n871), .A2(new_n873), .A3(new_n874), .A4(new_n845), .ZN(G63));
  NAND2_X1  g689(.A1(G217), .A2(G902), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT60), .Z(new_n877));
  NAND2_X1  g691(.A1(new_n837), .A2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n837), .A2(KEYINPUT120), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n600), .B(KEYINPUT121), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n880), .A2(new_n244), .A3(new_n881), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n847), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n884), .A2(KEYINPUT61), .A3(new_n847), .A4(new_n885), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(G66));
  OAI21_X1  g704(.A(G953), .B1(new_n471), .B2(new_n354), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT122), .Z(new_n892));
  OAI21_X1  g706(.A(new_n791), .B1(new_n800), .B2(new_n802), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n228), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n392), .B(new_n393), .C1(G898), .C2(new_n228), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n896), .B(new_n897), .ZN(G69));
  INV_X1    g712(.A(new_n718), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n743), .A2(new_n349), .A3(new_n677), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n750), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n822), .ZN(new_n902));
  AND4_X1   g716(.A1(new_n716), .A2(new_n901), .A3(new_n744), .A4(new_n902), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n903), .A2(KEYINPUT124), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(KEYINPUT124), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n228), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n310), .A2(new_n311), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n450), .B1(new_n449), .B2(new_n208), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n907), .B(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(G900), .B2(new_n895), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  AOI211_X1 g725(.A(new_n691), .B(new_n630), .C1(new_n576), .C2(new_n594), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n349), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT123), .Z(new_n914));
  AND3_X1   g728(.A1(new_n744), .A2(new_n750), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n648), .A2(new_n902), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n916), .A2(KEYINPUT62), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(KEYINPUT62), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n909), .B1(new_n919), .B2(new_n895), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n911), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n228), .B1(G227), .B2(G900), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(G72));
  NAND3_X1  g737(.A1(new_n904), .A2(new_n894), .A3(new_n905), .ZN(new_n924));
  XNOR2_X1  g738(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n246), .A2(new_n235), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n925), .B(new_n926), .Z(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AOI211_X1 g742(.A(new_n324), .B(new_n342), .C1(new_n924), .C2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n930), .B2(new_n893), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n931), .A2(KEYINPUT126), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(KEYINPUT126), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n932), .A2(new_n933), .A3(new_n634), .ZN(new_n934));
  INV_X1    g748(.A(new_n343), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n336), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n927), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n935), .B2(new_n937), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n828), .B2(new_n829), .ZN(new_n940));
  NOR4_X1   g754(.A1(new_n929), .A2(new_n934), .A3(new_n845), .A4(new_n940), .ZN(G57));
endmodule


