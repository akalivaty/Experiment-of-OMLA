//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n538, new_n539, new_n540, new_n541, new_n542, new_n544,
    new_n546, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(KEYINPUT66), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n462), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n459), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n464), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n465), .B2(new_n467), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n471), .A2(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n474), .A2(G136), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n459), .B1(new_n465), .B2(new_n467), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  OAI211_X1 g060(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n489), .A3(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n492), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n462), .A2(new_n468), .A3(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n491), .B1(new_n494), .B2(new_n496), .ZN(G164));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT67), .B1(new_n498), .B2(KEYINPUT6), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(G651), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n499), .A2(new_n502), .B1(KEYINPUT6), .B2(new_n498), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT68), .B1(new_n506), .B2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(new_n504), .A3(G543), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n505), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n503), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n516), .A2(new_n498), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n515), .A2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT70), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n503), .A2(new_n510), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n503), .A2(G543), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT69), .B(G51), .Z(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n522), .A2(new_n524), .A3(new_n527), .A4(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  XOR2_X1   g105(.A(KEYINPUT71), .B(G90), .Z(new_n531));
  NAND2_X1  g106(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n525), .A2(G52), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n498), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(G171));
  NAND2_X1  g112(.A1(new_n525), .A2(G43), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n523), .A2(G81), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n538), .B(new_n539), .C1(new_n498), .C2(new_n540), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT72), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  AND3_X1   g118(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT73), .ZN(G188));
  NAND2_X1  g124(.A1(new_n510), .A2(G65), .ZN(new_n550));
  NAND2_X1  g125(.A1(G78), .A2(G543), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g127(.A(KEYINPUT74), .B1(new_n552), .B2(G651), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n554));
  AOI211_X1 g129(.A(new_n554), .B(new_n498), .C1(new_n550), .C2(new_n551), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT9), .B1(new_n513), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n503), .A2(new_n559), .A3(G53), .A4(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n523), .A2(G91), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n556), .A2(new_n563), .ZN(G299));
  OAI21_X1  g139(.A(KEYINPUT75), .B1(new_n534), .B2(new_n536), .ZN(new_n565));
  INV_X1    g140(.A(new_n536), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT75), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n566), .A2(new_n567), .A3(new_n533), .A4(new_n532), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n565), .A2(new_n568), .ZN(G301));
  NAND2_X1  g144(.A1(new_n525), .A2(G49), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n523), .A2(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  AND2_X1   g149(.A1(G73), .A2(G543), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n510), .B2(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n574), .B1(new_n576), .B2(new_n498), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  AOI211_X1 g153(.A(new_n578), .B(new_n505), .C1(new_n507), .C2(new_n509), .ZN(new_n579));
  OAI211_X1 g154(.A(KEYINPUT76), .B(G651), .C1(new_n579), .C2(new_n575), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n503), .A2(new_n510), .A3(G86), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n503), .A2(G48), .A3(G543), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n581), .A2(new_n585), .ZN(G305));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  XOR2_X1   g162(.A(KEYINPUT77), .B(G47), .Z(new_n588));
  OAI22_X1  g163(.A1(new_n587), .A2(new_n511), .B1(new_n513), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n498), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  NAND3_X1  g168(.A1(new_n523), .A2(KEYINPUT10), .A3(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n511), .B2(new_n596), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n510), .A2(G66), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G651), .ZN(new_n602));
  INV_X1    g177(.A(G54), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n513), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  MUX2_X1   g181(.A(new_n606), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g182(.A(new_n606), .B(G301), .S(G868), .Z(G321));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(G299), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n609), .B2(G168), .ZN(G297));
  OAI21_X1  g186(.A(new_n610), .B1(new_n609), .B2(G168), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n605), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n605), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g193(.A1(new_n462), .A2(new_n468), .A3(new_n472), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT78), .B(G2100), .Z(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT79), .ZN(new_n626));
  INV_X1    g201(.A(G111), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n625), .A2(new_n626), .B1(new_n627), .B2(G2105), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n626), .B2(new_n625), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n474), .A2(G135), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n480), .A2(G123), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2096), .Z(new_n633));
  NAND3_X1  g208(.A1(new_n623), .A2(new_n624), .A3(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G1341), .B(G1348), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT81), .ZN(new_n649));
  OAI21_X1  g224(.A(G14), .B1(new_n646), .B2(new_n647), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n654), .A2(KEYINPUT17), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n652), .A2(new_n653), .ZN(new_n656));
  AOI21_X1  g231(.A(KEYINPUT18), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n654), .B2(KEYINPUT18), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n657), .B(new_n659), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2100), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT82), .B(G2096), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  AND2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n669), .A2(new_n670), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n668), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n668), .A2(new_n671), .A3(new_n675), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1991), .B(G1996), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G229));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G32), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n472), .A2(G105), .ZN(new_n690));
  NAND3_X1  g265(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT26), .ZN(new_n692));
  AOI211_X1 g267(.A(new_n690), .B(new_n692), .C1(G129), .C2(new_n480), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n474), .A2(G141), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT90), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n689), .B1(new_n696), .B2(G29), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT27), .B(G1996), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(G27), .A2(G29), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G164), .B2(G29), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G2078), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT31), .B(G11), .ZN(new_n706));
  INV_X1    g281(.A(G28), .ZN(new_n707));
  AOI21_X1  g282(.A(G29), .B1(new_n707), .B2(KEYINPUT30), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(KEYINPUT93), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(KEYINPUT93), .ZN(new_n710));
  OR3_X1    g285(.A1(new_n707), .A2(KEYINPUT92), .A3(KEYINPUT30), .ZN(new_n711));
  OAI21_X1  g286(.A(KEYINPUT92), .B1(new_n707), .B2(KEYINPUT30), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  OAI221_X1 g288(.A(new_n706), .B1(new_n709), .B2(new_n713), .C1(new_n632), .C2(new_n687), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n702), .B2(new_n703), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT94), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT24), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n687), .B1(new_n717), .B2(G34), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(KEYINPUT89), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(KEYINPUT89), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n717), .B2(G34), .ZN(new_n721));
  AOI22_X1  g296(.A1(G160), .A2(G29), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(G2084), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n705), .B(new_n715), .C1(new_n716), .C2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n725), .A2(G21), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G286), .B2(G16), .ZN(new_n727));
  INV_X1    g302(.A(G1966), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G171), .A2(new_n725), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G5), .B2(new_n725), .ZN(new_n731));
  INV_X1    g306(.A(G1961), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n729), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n474), .A2(G140), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n480), .A2(G128), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n459), .A2(G116), .ZN(new_n736));
  OAI21_X1  g311(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n734), .B(new_n735), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G29), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT87), .ZN(new_n740));
  INV_X1    g315(.A(G26), .ZN(new_n741));
  OAI21_X1  g316(.A(KEYINPUT28), .B1(new_n741), .B2(G29), .ZN(new_n742));
  OR3_X1    g317(.A1(new_n741), .A2(KEYINPUT28), .A3(G29), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n740), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT88), .B(G2067), .ZN(new_n745));
  OAI22_X1  g320(.A1(new_n744), .A2(new_n745), .B1(new_n727), .B2(new_n728), .ZN(new_n746));
  NOR3_X1   g321(.A1(new_n724), .A2(new_n733), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n605), .A2(G16), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G4), .B2(G16), .ZN(new_n749));
  INV_X1    g324(.A(G1348), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n749), .A2(new_n750), .B1(new_n716), .B2(new_n723), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n747), .B(new_n751), .C1(new_n750), .C2(new_n749), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n542), .A2(new_n725), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n725), .B2(G19), .ZN(new_n754));
  INV_X1    g329(.A(G1341), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n731), .A2(new_n732), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n687), .A2(G35), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G162), .B2(new_n687), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT29), .Z(new_n761));
  INV_X1    g336(.A(G2090), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n744), .A2(new_n745), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n756), .A2(new_n757), .A3(new_n758), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n687), .A2(G33), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT25), .Z(new_n767));
  INV_X1    g342(.A(G139), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n475), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n462), .A2(new_n468), .A3(G127), .ZN(new_n770));
  INV_X1    g345(.A(G115), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(new_n464), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n769), .B1(new_n772), .B2(G2105), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n765), .B1(new_n773), .B2(new_n687), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(G2072), .Z(new_n775));
  AOI22_X1  g350(.A1(new_n697), .A2(new_n698), .B1(new_n722), .B2(G2084), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT91), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n752), .A2(new_n764), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n725), .A2(G20), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT23), .Z(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G299), .B2(G16), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT95), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G1956), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n761), .A2(new_n762), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT96), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n779), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT97), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n725), .A2(G23), .ZN(new_n797));
  INV_X1    g372(.A(G288), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n725), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT33), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1976), .ZN(new_n801));
  MUX2_X1   g376(.A(G6), .B(G305), .S(G16), .Z(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT32), .B(G1981), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n725), .A2(G22), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT86), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G166), .B2(new_n725), .ZN(new_n808));
  INV_X1    g383(.A(G1971), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n801), .A2(new_n804), .A3(new_n805), .A4(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n687), .A2(G25), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n474), .A2(G131), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n480), .A2(G119), .ZN(new_n816));
  OR2_X1    g391(.A1(G95), .A2(G2105), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n817), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n814), .B1(new_n820), .B2(new_n687), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT35), .B(G1991), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n725), .A2(G24), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT84), .Z(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n592), .B2(new_n725), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT85), .B(G1986), .Z(new_n827));
  OAI21_X1  g402(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n826), .B2(new_n827), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n812), .A2(new_n813), .A3(new_n829), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(KEYINPUT36), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(KEYINPUT36), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n795), .A2(new_n796), .B1(new_n831), .B2(new_n832), .ZN(G311));
  NAND2_X1  g408(.A1(new_n795), .A2(new_n796), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n831), .A2(new_n832), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(G150));
  NAND2_X1  g411(.A1(new_n605), .A2(G559), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT38), .Z(new_n838));
  AOI22_X1  g413(.A1(G93), .A2(new_n523), .B1(new_n525), .B2(G55), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n498), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(new_n541), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n542), .A2(new_n841), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n838), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n848));
  AOI21_X1  g423(.A(G860), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n848), .B2(new_n847), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT99), .ZN(new_n851));
  INV_X1    g426(.A(new_n843), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(G860), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n851), .A2(new_n854), .ZN(G145));
  NAND2_X1  g430(.A1(new_n480), .A2(G130), .ZN(new_n856));
  OR2_X1    g431(.A1(G106), .A2(G2105), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n857), .B(G2104), .C1(G118), .C2(new_n459), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(G142), .B2(new_n474), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n620), .B(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n861), .A2(new_n819), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n819), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n773), .B(new_n696), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n865), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n862), .A2(new_n867), .A3(new_n863), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n494), .A2(new_n496), .ZN(new_n870));
  INV_X1    g445(.A(new_n491), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n738), .ZN(new_n873));
  XNOR2_X1  g448(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n873), .B(new_n874), .Z(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n866), .A2(new_n875), .A3(new_n868), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(G160), .B(G162), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n632), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(G37), .ZN(new_n883));
  INV_X1    g458(.A(new_n881), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n877), .A2(new_n884), .A3(new_n878), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n886), .A2(KEYINPUT102), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(KEYINPUT102), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g465(.A1(new_n852), .A2(new_n609), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n846), .B(new_n615), .ZN(new_n892));
  XNOR2_X1  g467(.A(G299), .B(new_n605), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n893), .B(KEYINPUT103), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n898), .B1(new_n892), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(G290), .B(G305), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n798), .B(G303), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n901), .B(new_n902), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n903), .B(KEYINPUT42), .Z(new_n904));
  XNOR2_X1  g479(.A(new_n900), .B(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n891), .B1(new_n905), .B2(new_n609), .ZN(G295));
  OAI21_X1  g481(.A(new_n891), .B1(new_n905), .B2(new_n609), .ZN(G331));
  NOR2_X1   g482(.A1(G301), .A2(G286), .ZN(new_n908));
  NOR2_X1   g483(.A1(G168), .A2(G171), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n844), .B(new_n845), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n846), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n899), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n896), .A2(KEYINPUT105), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT105), .B1(new_n895), .B2(new_n896), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n913), .B(new_n903), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n914), .A2(new_n897), .ZN(new_n919));
  INV_X1    g494(.A(new_n903), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n912), .A2(new_n893), .A3(new_n910), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n918), .A2(new_n883), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n923), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n924));
  XOR2_X1   g499(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  AOI22_X1  g501(.A1(new_n910), .A2(new_n912), .B1(new_n895), .B2(new_n896), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n912), .A2(new_n893), .A3(new_n910), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n903), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n922), .A3(new_n883), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n924), .B(KEYINPUT44), .C1(new_n926), .C2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT106), .B1(new_n923), .B2(KEYINPUT43), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n930), .A2(new_n926), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n923), .A2(new_n926), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI22_X1  g510(.A1(new_n931), .A2(new_n932), .B1(new_n935), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g511(.A(KEYINPUT50), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n938));
  INV_X1    g513(.A(G1384), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n872), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT110), .B1(G164), .B2(G1384), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n872), .A2(new_n937), .A3(new_n939), .ZN(new_n943));
  INV_X1    g518(.A(G40), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n471), .A2(new_n477), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n785), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n872), .A2(KEYINPUT45), .A3(new_n939), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n948), .A2(new_n945), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT45), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n950), .B1(G164), .B2(G1384), .ZN(new_n951));
  XNOR2_X1  g526(.A(KEYINPUT56), .B(G2072), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT118), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n949), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n955));
  NAND2_X1  g530(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n556), .A2(new_n563), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n553), .A2(new_n555), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n561), .A2(new_n562), .ZN(new_n959));
  OAI211_X1 g534(.A(KEYINPUT117), .B(KEYINPUT57), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n947), .A2(new_n954), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n947), .A2(new_n957), .A3(new_n954), .A4(new_n960), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n945), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n940), .A2(new_n941), .A3(new_n937), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n750), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n940), .A2(new_n945), .A3(new_n941), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(G2067), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n606), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n961), .B1(new_n962), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT61), .ZN(new_n973));
  AND4_X1   g548(.A1(new_n947), .A2(new_n957), .A3(new_n954), .A4(new_n960), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(new_n961), .ZN(new_n975));
  AOI21_X1  g550(.A(G1348), .B1(new_n964), .B2(new_n965), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n976), .A2(new_n969), .A3(new_n605), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT60), .B1(new_n971), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT120), .ZN(new_n980));
  XOR2_X1   g555(.A(KEYINPUT58), .B(G1341), .Z(new_n981));
  AND3_X1   g556(.A1(new_n968), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n980), .B1(new_n968), .B2(new_n981), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n948), .A2(new_n945), .A3(new_n951), .ZN(new_n984));
  XNOR2_X1  g559(.A(KEYINPUT119), .B(G1996), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n982), .A2(new_n983), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n542), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n979), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n979), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n542), .A2(new_n988), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n983), .A2(new_n986), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n991), .B(new_n992), .C1(new_n993), .C2(new_n982), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n975), .A2(new_n978), .A3(new_n990), .A4(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n961), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n996), .A2(KEYINPUT61), .A3(new_n962), .ZN(new_n997));
  OR4_X1    g572(.A1(KEYINPUT60), .A2(new_n976), .A3(new_n606), .A4(new_n969), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n972), .B1(new_n995), .B2(new_n999), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n940), .A2(new_n941), .A3(new_n937), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n945), .A2(new_n963), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n732), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n938), .B1(new_n872), .B2(new_n939), .ZN(new_n1004));
  NOR3_X1   g579(.A1(G164), .A2(KEYINPUT110), .A3(G1384), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n950), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1007), .A2(G2078), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n949), .A3(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n948), .A2(new_n945), .A3(new_n951), .A4(new_n703), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n1007), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1003), .A2(new_n1009), .A3(G301), .A4(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT124), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n966), .A2(new_n732), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1015), .A2(KEYINPUT124), .A3(G301), .A4(new_n1009), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT123), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n949), .A2(new_n1019), .A3(new_n951), .A4(new_n1008), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1008), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT123), .B1(new_n984), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1015), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1018), .B1(new_n1024), .B2(G171), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1017), .A2(new_n1025), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1001), .A2(G2084), .A3(new_n1002), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1966), .B1(new_n1006), .B2(new_n949), .ZN(new_n1028));
  OAI21_X1  g603(.A(G8), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(G286), .A2(G8), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT122), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT51), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1029), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT45), .B1(new_n940), .B2(new_n941), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n948), .A2(new_n945), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n728), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(G2084), .B2(new_n966), .ZN(new_n1038));
  OAI211_X1 g613(.A(G8), .B(new_n1032), .C1(new_n1038), .C2(G286), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(G8), .A3(G286), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1034), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1015), .A2(new_n1023), .A3(G301), .ZN(new_n1042));
  AOI21_X1  g617(.A(G301), .B1(new_n1015), .B2(new_n1009), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1018), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1026), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G303), .A2(G8), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n984), .A2(new_n809), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT50), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n943), .A2(new_n945), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(G2090), .B1(new_n1054), .B2(KEYINPUT115), .ZN(new_n1055));
  OR3_X1    g630(.A1(new_n942), .A2(KEYINPUT115), .A3(new_n946), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1051), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G8), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1049), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n964), .A2(new_n965), .A3(new_n762), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT111), .B1(new_n1060), .B2(new_n1050), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1060), .A2(KEYINPUT111), .A3(new_n1050), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1062), .A2(G8), .A3(new_n1048), .A4(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n1065));
  INV_X1    g640(.A(G1981), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n581), .B2(new_n585), .ZN(new_n1067));
  AOI211_X1 g642(.A(G1981), .B(new_n584), .C1(new_n577), .C2(new_n580), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1065), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT49), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n968), .A2(G8), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT49), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1065), .B(new_n1072), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n798), .A2(G1976), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1075), .A2(G8), .A3(new_n968), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(KEYINPUT112), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1075), .A2(new_n968), .A3(G8), .A4(new_n1078), .ZN(new_n1081));
  OR3_X1    g656(.A1(new_n798), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1074), .A2(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1059), .A2(new_n1064), .A3(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1000), .A2(new_n1045), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1063), .A2(G8), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1048), .B1(new_n1088), .B2(new_n1062), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1074), .A2(new_n1083), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1087), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1063), .A2(G8), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1049), .B1(new_n1092), .B2(new_n1061), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1084), .A2(new_n1093), .A3(KEYINPUT116), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1029), .A2(G286), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1064), .A2(new_n1095), .A3(KEYINPUT63), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1091), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1059), .A2(new_n1084), .A3(new_n1064), .A4(new_n1095), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT63), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(G288), .A2(G1976), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1103), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1071), .B1(new_n1104), .B2(new_n1068), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1064), .B2(new_n1090), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1105), .B(KEYINPUT114), .C1(new_n1064), .C2(new_n1090), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1086), .A2(new_n1101), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1086), .A2(new_n1101), .A3(KEYINPUT125), .A4(new_n1110), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1041), .A2(KEYINPUT62), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1041), .A2(KEYINPUT62), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1115), .A2(new_n1085), .A3(new_n1043), .A4(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n477), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n469), .A2(new_n470), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1119), .B(G40), .C1(new_n1120), .C2(new_n459), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(new_n951), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1122), .B(KEYINPUT107), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1123), .A2(G1996), .A3(new_n696), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT108), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1127));
  INV_X1    g702(.A(G2067), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n738), .B(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(G1996), .B2(new_n696), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1123), .A2(new_n1130), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1126), .A2(new_n1127), .A3(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n819), .B(new_n822), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n1133), .B(KEYINPUT109), .Z(new_n1134));
  NAND2_X1  g709(.A1(new_n1123), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(G1986), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n592), .B(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1136), .B1(new_n1123), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1118), .A2(new_n1139), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1132), .A2(new_n822), .A3(new_n820), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n738), .A2(G2067), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1123), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(G1996), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1123), .A2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT46), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1129), .A2(new_n695), .A3(new_n693), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1123), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT47), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1123), .A2(new_n1137), .A3(new_n592), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT48), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1132), .A2(new_n1135), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1143), .A2(new_n1150), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT126), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1143), .A2(new_n1153), .A3(new_n1156), .A4(new_n1150), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1140), .A2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n1161));
  INV_X1    g735(.A(G227), .ZN(new_n1162));
  AND2_X1   g736(.A1(new_n1162), .A2(G319), .ZN(new_n1163));
  NAND2_X1  g737(.A1(new_n685), .A2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g738(.A(new_n1161), .B1(new_n1164), .B2(G401), .ZN(new_n1165));
  INV_X1    g739(.A(G401), .ZN(new_n1166));
  NAND4_X1  g740(.A1(new_n1166), .A2(KEYINPUT127), .A3(new_n685), .A4(new_n1163), .ZN(new_n1167));
  AOI22_X1  g741(.A1(new_n1165), .A2(new_n1167), .B1(new_n887), .B2(new_n888), .ZN(new_n1168));
  OR2_X1    g742(.A1(new_n933), .A2(new_n934), .ZN(new_n1169));
  AND2_X1   g743(.A1(new_n1168), .A2(new_n1169), .ZN(G308));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(G225));
endmodule


