//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n191), .A3(new_n195), .A4(new_n192), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT70), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(KEYINPUT70), .A3(new_n196), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT10), .ZN(new_n203));
  INV_X1    g017(.A(G107), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT79), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT79), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G107), .ZN(new_n207));
  AOI21_X1  g021(.A(G104), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT82), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G107), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n204), .A2(KEYINPUT82), .A3(G104), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(G101), .B1(new_n208), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n210), .A2(KEYINPUT3), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n205), .A3(new_n207), .ZN(new_n216));
  INV_X1    g030(.A(G101), .ZN(new_n217));
  OAI21_X1  g031(.A(G107), .B1(new_n210), .B2(KEYINPUT3), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n210), .A2(KEYINPUT3), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT65), .A2(G146), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(G143), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n224), .A2(G143), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n227), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n227), .A2(KEYINPUT67), .A3(new_n229), .A4(new_n231), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(KEYINPUT65), .A2(G146), .ZN(new_n237));
  NOR2_X1   g051(.A1(KEYINPUT65), .A2(G146), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n228), .B1(new_n239), .B2(G143), .ZN(new_n240));
  INV_X1    g054(.A(G143), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT1), .B1(new_n241), .B2(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G128), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT83), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n227), .A2(new_n229), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT83), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(new_n243), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n203), .B(new_n222), .C1(new_n236), .C2(new_n249), .ZN(new_n250));
  NOR3_X1   g064(.A1(new_n237), .A2(new_n238), .A3(new_n241), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT1), .ZN(new_n252));
  OAI21_X1  g066(.A(G128), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(new_n241), .B2(G146), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n224), .A2(KEYINPUT64), .A3(G143), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n255), .B(new_n256), .C1(new_n239), .C2(G143), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n234), .A2(new_n235), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT10), .B1(new_n258), .B2(new_n221), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n250), .A2(new_n259), .ZN(new_n260));
  AND2_X1   g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  NOR2_X1   g075(.A1(KEYINPUT0), .A2(G128), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(G143), .B1(new_n225), .B2(new_n226), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n255), .A2(new_n256), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n227), .A2(new_n229), .A3(new_n261), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n220), .A2(KEYINPUT4), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G101), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n268), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT4), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n270), .A2(new_n273), .A3(G101), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT80), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT80), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n270), .A2(new_n276), .A3(new_n273), .A4(G101), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n272), .A2(new_n278), .A3(KEYINPUT81), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT81), .B1(new_n272), .B2(new_n278), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n260), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT86), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n202), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n260), .B(KEYINPUT86), .C1(new_n279), .C2(new_n280), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n260), .B(new_n202), .C1(new_n279), .C2(new_n280), .ZN(new_n286));
  XNOR2_X1  g100(.A(G110), .B(G140), .ZN(new_n287));
  INV_X1    g101(.A(G227), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(G953), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n287), .B(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT85), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n286), .A2(KEYINPUT85), .A3(new_n291), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n285), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  AOI221_X4 g110(.A(KEYINPUT83), .B1(new_n242), .B2(G128), .C1(new_n227), .C2(new_n229), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n247), .B1(new_n246), .B2(new_n243), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n234), .A2(new_n235), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n221), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n253), .A2(new_n257), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n300), .A2(new_n302), .A3(new_n221), .ZN(new_n303));
  OAI211_X1 g117(.A(KEYINPUT12), .B(new_n197), .C1(new_n301), .C2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT84), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n222), .B1(new_n236), .B2(new_n249), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n258), .A2(new_n221), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n202), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n306), .B1(new_n309), .B2(KEYINPUT12), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n201), .B1(new_n301), .B2(new_n303), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT12), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(KEYINPUT84), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n305), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n286), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n290), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n296), .A2(G469), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G469), .ZN(new_n318));
  INV_X1    g132(.A(G902), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT87), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n314), .B2(new_n292), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n309), .A2(new_n306), .A3(KEYINPUT12), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT84), .B1(new_n311), .B2(new_n312), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n304), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n286), .A2(new_n291), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT87), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n315), .B1(new_n283), .B2(new_n284), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n324), .B(new_n329), .C1(new_n330), .C2(new_n291), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n318), .A3(new_n319), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n322), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G113), .B(G122), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(new_n210), .ZN(new_n335));
  INV_X1    g149(.A(G140), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G125), .ZN(new_n337));
  INV_X1    g151(.A(G125), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G140), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(new_n339), .A3(KEYINPUT16), .ZN(new_n340));
  OR3_X1    g154(.A1(new_n338), .A2(KEYINPUT16), .A3(G140), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(G146), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(G146), .B1(new_n340), .B2(new_n341), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G237), .ZN(new_n346));
  INV_X1    g160(.A(G953), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n347), .A3(G214), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n241), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n346), .A2(new_n347), .A3(G143), .A4(G214), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n195), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(KEYINPUT89), .A3(KEYINPUT17), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT89), .B1(new_n351), .B2(KEYINPUT17), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n345), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT90), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n351), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT17), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n349), .A2(new_n195), .A3(new_n350), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(KEYINPUT90), .B(new_n345), .C1(new_n353), .C2(new_n354), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n357), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n337), .A2(new_n339), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT88), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G146), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n239), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n349), .A2(new_n350), .ZN(new_n369));
  NAND2_X1  g183(.A1(KEYINPUT18), .A2(G131), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n369), .B(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n335), .B1(new_n363), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n362), .A2(new_n361), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n369), .A2(KEYINPUT17), .A3(G131), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT89), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n352), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT90), .B1(new_n378), .B2(new_n345), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n335), .B(new_n372), .C1(new_n374), .C2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT91), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n363), .A2(KEYINPUT91), .A3(new_n335), .A4(new_n372), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n373), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(G475), .B1(new_n384), .B2(G902), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n205), .A2(new_n207), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT92), .B(G122), .ZN(new_n387));
  INV_X1    g201(.A(G116), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(G122), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n386), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n386), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n393), .B(new_n390), .C1(new_n388), .C2(new_n387), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT93), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n396), .B1(new_n230), .B2(G143), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n241), .A2(KEYINPUT93), .A3(G128), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n230), .A2(G143), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n188), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n395), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT13), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n399), .A2(new_n403), .B1(new_n230), .B2(G143), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n397), .A2(KEYINPUT13), .A3(new_n398), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n188), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT94), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n406), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT94), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n408), .A2(new_n395), .A3(new_n409), .A4(new_n401), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n399), .A2(new_n400), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G134), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n401), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n390), .B(KEYINPUT14), .ZN(new_n414));
  OAI21_X1  g228(.A(G107), .B1(new_n414), .B2(new_n389), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n394), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n407), .A2(new_n410), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT9), .B(G234), .ZN(new_n418));
  INV_X1    g232(.A(G217), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n418), .A2(new_n419), .A3(G953), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n407), .A2(new_n410), .A3(new_n416), .A4(new_n420), .ZN(new_n423));
  AOI21_X1  g237(.A(G902), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G478), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(KEYINPUT15), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n424), .B(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n382), .A2(new_n383), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n343), .B1(new_n358), .B2(new_n360), .ZN(new_n430));
  MUX2_X1   g244(.A(new_n364), .B(new_n365), .S(KEYINPUT19), .Z(new_n431));
  INV_X1    g245(.A(new_n239), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n335), .B1(new_n433), .B2(new_n372), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(G475), .A2(G902), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n428), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n434), .B1(new_n382), .B2(new_n383), .ZN(new_n439));
  INV_X1    g253(.A(new_n437), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n439), .A2(KEYINPUT20), .A3(new_n440), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n385), .B(new_n427), .C1(new_n438), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(G234), .A2(G237), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(G952), .A3(new_n347), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(G898), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n443), .A2(G902), .A3(G953), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n444), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G214), .B1(G237), .B2(G902), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n268), .A2(G125), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n300), .A2(new_n302), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n450), .B1(new_n451), .B2(G125), .ZN(new_n452));
  INV_X1    g266(.A(G224), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT7), .B1(new_n453), .B2(G953), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n452), .B(new_n454), .Z(new_n455));
  XNOR2_X1  g269(.A(G110), .B(G122), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(KEYINPUT8), .ZN(new_n457));
  INV_X1    g271(.A(G113), .ZN(new_n458));
  INV_X1    g272(.A(G119), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G116), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT5), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n388), .A2(G119), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n463), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(KEYINPUT2), .A2(G113), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT68), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT68), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(KEYINPUT2), .A3(G113), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT2), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n468), .A2(new_n470), .B1(new_n471), .B2(new_n458), .ZN(new_n472));
  XNOR2_X1  g286(.A(G116), .B(G119), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n466), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n457), .B1(new_n475), .B2(new_n221), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n465), .A2(KEYINPUT69), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT69), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT5), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n481), .A2(new_n463), .B1(new_n472), .B2(new_n473), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n476), .B1(new_n221), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n269), .A2(new_n271), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n468), .A2(new_n470), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n471), .A2(new_n458), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n477), .A3(new_n479), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n474), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n490), .A2(new_n278), .B1(new_n222), .B2(new_n482), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n483), .B1(new_n491), .B2(new_n456), .ZN(new_n492));
  AOI21_X1  g306(.A(G902), .B1(new_n455), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n482), .A2(new_n222), .ZN(new_n494));
  INV_X1    g308(.A(new_n278), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n484), .A2(new_n489), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n456), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n494), .B(new_n456), .C1(new_n495), .C2(new_n496), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(KEYINPUT6), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n497), .A2(new_n502), .A3(new_n498), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n453), .A2(G953), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n452), .B(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n501), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(G210), .B1(G237), .B2(G902), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n493), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n507), .B1(new_n493), .B2(new_n506), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n448), .B(new_n449), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n442), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(G221), .B1(new_n418), .B2(G902), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n333), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT32), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT71), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n190), .A2(G134), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT66), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n192), .A3(new_n517), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n518), .B(G131), .C1(new_n517), .C2(new_n516), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n196), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n451), .A2(new_n515), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT71), .B1(new_n258), .B2(new_n520), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT72), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n488), .A2(new_n524), .A3(new_n474), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n524), .B1(new_n488), .B2(new_n474), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n268), .ZN(new_n528));
  INV_X1    g342(.A(new_n200), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT70), .B1(new_n194), .B2(new_n196), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n522), .A2(new_n523), .A3(new_n527), .A4(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n346), .A2(new_n347), .A3(G210), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(KEYINPUT27), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT26), .B(G101), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n534), .B(new_n535), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT31), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n197), .A2(new_n267), .A3(new_n266), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n539), .B(new_n540), .C1(new_n258), .C2(new_n520), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n522), .A2(new_n523), .A3(new_n531), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n542), .B1(new_n543), .B2(KEYINPUT30), .ZN(new_n544));
  INV_X1    g358(.A(new_n489), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n537), .B(new_n538), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n536), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT28), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n520), .B1(new_n300), .B2(new_n302), .ZN(new_n549));
  INV_X1    g363(.A(new_n540), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n489), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n548), .B1(new_n532), .B2(new_n551), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n525), .A2(new_n526), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(new_n549), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT28), .B1(new_n554), .B2(new_n531), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n547), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n546), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n543), .A2(KEYINPUT30), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n545), .B1(new_n558), .B2(new_n541), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n532), .A2(new_n536), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT31), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT73), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n537), .B1(new_n544), .B2(new_n545), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT73), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT31), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n557), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(G472), .A2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n514), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n546), .A2(new_n556), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT31), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n564), .B1(new_n563), .B2(KEYINPUT31), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(KEYINPUT32), .A3(new_n567), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n543), .A2(new_n553), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n532), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n555), .B1(new_n576), .B2(KEYINPUT28), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT29), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n547), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(G902), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n532), .B1(new_n544), .B2(new_n545), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n547), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n532), .A2(new_n551), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT28), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT74), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n527), .B1(new_n258), .B2(new_n520), .ZN(new_n586));
  INV_X1    g400(.A(new_n531), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n548), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n584), .A2(new_n585), .A3(new_n536), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n582), .A2(new_n578), .A3(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n552), .A2(new_n555), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n585), .B1(new_n591), .B2(new_n536), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n580), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G472), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n569), .A2(new_n574), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT78), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT75), .B1(new_n230), .B2(G119), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT23), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n598), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n459), .A2(G128), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(G119), .B(G128), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT24), .B(G110), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n602), .A2(G110), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(new_n344), .B2(new_n343), .ZN(new_n607));
  OAI22_X1  g421(.A1(new_n602), .A2(G110), .B1(new_n603), .B2(new_n605), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(new_n342), .A3(new_n367), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT22), .B(G137), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n347), .A2(G221), .A3(G234), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT76), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n607), .A2(new_n609), .A3(new_n613), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(KEYINPUT25), .A3(new_n319), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT25), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n618), .B2(G902), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n620), .A2(KEYINPUT77), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n419), .B1(G234), .B2(new_n319), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n624), .B1(new_n622), .B2(KEYINPUT77), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n624), .A2(G902), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n626), .B1(new_n619), .B2(new_n627), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n595), .A2(new_n596), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n596), .B1(new_n595), .B2(new_n628), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n513), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G101), .ZN(G3));
  INV_X1    g446(.A(KEYINPUT95), .ZN(new_n633));
  INV_X1    g447(.A(G472), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n566), .A2(G902), .A3(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n635), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n573), .B2(new_n319), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n512), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n322), .B2(new_n332), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n639), .A2(new_n641), .A3(new_n628), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n385), .B1(new_n438), .B2(new_n441), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n422), .A2(new_n423), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT33), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT33), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n422), .A2(new_n646), .A3(new_n423), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n645), .A2(G478), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n425), .A2(new_n319), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(new_n424), .B2(new_n425), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n643), .A2(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n642), .A2(new_n510), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT34), .B(G104), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  NOR4_X1   g470(.A1(new_n439), .A2(KEYINPUT97), .A3(KEYINPUT20), .A4(new_n440), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n436), .A2(new_n428), .A3(new_n437), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT97), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT96), .ZN(new_n661));
  OAI21_X1  g475(.A(KEYINPUT20), .B1(new_n439), .B2(new_n440), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n658), .A2(new_n660), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n661), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT97), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n441), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n664), .B1(new_n666), .B2(new_n657), .ZN(new_n667));
  INV_X1    g481(.A(new_n385), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n427), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n663), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n642), .A2(new_n510), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT98), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT35), .B(G107), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  OR2_X1    g488(.A1(new_n623), .A2(new_n625), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT36), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n614), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n610), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n610), .A2(new_n677), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n627), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n680), .B(KEYINPUT99), .Z(new_n681));
  NAND2_X1  g495(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n639), .A2(new_n641), .A3(new_n511), .A4(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  INV_X1    g499(.A(new_n449), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n493), .A2(new_n506), .ZN(new_n687));
  INV_X1    g501(.A(new_n507), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n493), .A2(new_n506), .A3(new_n507), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n686), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  OR2_X1    g506(.A1(new_n447), .A2(G900), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n444), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n670), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n595), .A2(new_n682), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n697), .A3(new_n641), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G128), .ZN(G30));
  NOR2_X1   g513(.A1(new_n508), .A2(new_n509), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT38), .Z(new_n701));
  INV_X1    g515(.A(new_n581), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n547), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n319), .B1(new_n576), .B2(new_n536), .ZN(new_n704));
  OAI21_X1  g518(.A(G472), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n569), .A2(new_n574), .A3(new_n705), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n682), .A2(new_n686), .A3(new_n427), .ZN(new_n707));
  AND4_X1   g521(.A1(new_n643), .A2(new_n701), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n694), .B(KEYINPUT39), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n641), .A2(new_n709), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n708), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G143), .ZN(G45));
  NAND4_X1  g528(.A1(new_n691), .A2(new_n643), .A3(new_n652), .A4(new_n694), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT100), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n659), .A2(new_n662), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n651), .B1(new_n718), .B2(new_n385), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(KEYINPUT100), .A3(new_n691), .A4(new_n694), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n697), .A3(new_n641), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  AND2_X1   g537(.A1(new_n595), .A2(new_n628), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n331), .A2(new_n319), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(G469), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n512), .A3(new_n332), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT101), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n653), .A2(new_n510), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n726), .A2(KEYINPUT101), .A3(new_n512), .A4(new_n332), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n724), .A2(new_n729), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT41), .B(G113), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G15));
  INV_X1    g548(.A(new_n510), .ZN(new_n735));
  AND4_X1   g549(.A1(new_n735), .A2(new_n663), .A3(new_n667), .A4(new_n669), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n724), .A2(new_n729), .A3(new_n736), .A4(new_n731), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G116), .ZN(G18));
  AND3_X1   g552(.A1(new_n331), .A2(new_n318), .A3(new_n319), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n318), .B1(new_n331), .B2(new_n319), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n739), .A2(new_n740), .A3(new_n640), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(new_n595), .A3(new_n511), .A4(new_n682), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  INV_X1    g557(.A(KEYINPUT103), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n561), .A2(new_n546), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n549), .A2(new_n515), .B1(new_n201), .B2(new_n528), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n527), .B1(new_n746), .B2(new_n523), .ZN(new_n747));
  INV_X1    g561(.A(new_n532), .ZN(new_n748));
  OAI21_X1  g562(.A(KEYINPUT28), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n588), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT102), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n536), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n577), .A2(KEYINPUT102), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n745), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n744), .B1(new_n754), .B2(new_n568), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n750), .A2(new_n751), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n547), .B1(new_n577), .B2(KEYINPUT102), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI211_X1 g572(.A(KEYINPUT103), .B(new_n567), .C1(new_n758), .C2(new_n745), .ZN(new_n759));
  OAI21_X1  g573(.A(G472), .B1(new_n566), .B2(G902), .ZN(new_n760));
  AND4_X1   g574(.A1(new_n628), .A2(new_n755), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n427), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n643), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n510), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n729), .A2(new_n761), .A3(new_n731), .A4(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G122), .ZN(G24));
  NOR2_X1   g580(.A1(new_n727), .A2(new_n692), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n653), .A2(new_n695), .ZN(new_n768));
  AND4_X1   g582(.A1(new_n682), .A2(new_n755), .A3(new_n759), .A4(new_n760), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G125), .ZN(G27));
  NAND4_X1  g585(.A1(new_n689), .A2(new_n512), .A3(new_n449), .A4(new_n690), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n317), .A2(new_n321), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n773), .B1(new_n739), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT104), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n772), .B1(new_n322), .B2(new_n332), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT104), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n724), .A2(new_n776), .A3(new_n768), .A4(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT105), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(KEYINPUT42), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n777), .A2(new_n778), .ZN(new_n784));
  AOI211_X1 g598(.A(KEYINPUT104), .B(new_n772), .C1(new_n322), .C2(new_n332), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n782), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n786), .A2(new_n724), .A3(new_n768), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G131), .ZN(G33));
  AND4_X1   g604(.A1(new_n663), .A2(new_n667), .A3(new_n669), .A4(new_n694), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n724), .A2(new_n776), .A3(new_n791), .A4(new_n779), .ZN(new_n792));
  XNOR2_X1  g606(.A(KEYINPUT106), .B(G134), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(G36));
  INV_X1    g608(.A(new_n682), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n639), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n718), .A2(new_n652), .A3(new_n385), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT43), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT44), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT107), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT107), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n796), .A2(new_n799), .A3(new_n803), .A4(KEYINPUT44), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT45), .B1(new_n296), .B2(new_n316), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n318), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n296), .A2(KEYINPUT45), .A3(new_n316), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n320), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n809), .A2(KEYINPUT46), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n332), .B1(new_n809), .B2(KEYINPUT46), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n512), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n700), .A2(new_n449), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n814), .B(KEYINPUT108), .Z(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n800), .B2(new_n801), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n805), .A2(new_n709), .A3(new_n813), .A4(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G137), .ZN(G39));
  NOR2_X1   g632(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n812), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n822));
  OAI221_X1 g636(.A(new_n512), .B1(new_n822), .B2(new_n819), .C1(new_n810), .C2(new_n811), .ZN(new_n823));
  INV_X1    g637(.A(new_n768), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n824), .A2(new_n595), .A3(new_n628), .A4(new_n814), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n821), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G140), .ZN(G42));
  NAND2_X1  g641(.A1(new_n512), .A2(new_n449), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n701), .A2(new_n643), .A3(new_n651), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n739), .A2(new_n740), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT49), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n830), .B1(KEYINPUT110), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT110), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n832), .B1(new_n833), .B2(KEYINPUT49), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n830), .A2(KEYINPUT110), .A3(new_n831), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n829), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n628), .A2(new_n569), .A3(new_n574), .A4(new_n705), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n772), .A2(new_n444), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n830), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n797), .B(KEYINPUT43), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n724), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT48), .Z(new_n844));
  OR2_X1    g658(.A1(new_n840), .A2(new_n837), .ZN(new_n845));
  OAI211_X1 g659(.A(G952), .B(new_n347), .C1(new_n845), .C2(new_n653), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n841), .A2(new_n444), .ZN(new_n847));
  INV_X1    g661(.A(new_n761), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n849), .A2(new_n767), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n844), .A2(new_n846), .A3(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n845), .A2(new_n643), .A3(new_n652), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(new_n769), .B2(new_n842), .ZN(new_n853));
  INV_X1    g667(.A(new_n849), .ZN(new_n854));
  OR3_X1    g668(.A1(new_n701), .A2(new_n727), .A3(new_n449), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(KEYINPUT50), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT50), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n854), .A2(new_n858), .A3(new_n855), .ZN(new_n859));
  OAI211_X1 g673(.A(KEYINPUT51), .B(new_n853), .C1(new_n857), .C2(new_n859), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n854), .A2(new_n815), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n821), .A2(new_n823), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n830), .A2(new_n640), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n851), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT114), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n821), .A2(new_n823), .A3(KEYINPUT114), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n868), .A2(new_n869), .A3(new_n863), .ZN(new_n870));
  OAI221_X1 g684(.A(new_n853), .B1(new_n857), .B2(new_n859), .C1(new_n870), .C2(new_n861), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n865), .B1(new_n866), .B2(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n732), .A2(new_n737), .A3(new_n765), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n776), .A2(new_n769), .A3(new_n779), .A4(new_n768), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n762), .A2(new_n668), .A3(new_n695), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n663), .A2(new_n667), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n697), .A2(new_n777), .A3(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n792), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n641), .A2(new_n511), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n595), .A2(new_n628), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT78), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n595), .A2(new_n596), .A3(new_n628), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n718), .A2(new_n762), .A3(new_n385), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n510), .B1(new_n653), .B2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(new_n639), .A3(new_n641), .A4(new_n628), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n742), .A2(new_n886), .A3(new_n683), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n789), .A2(new_n873), .A3(new_n878), .A4(new_n888), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n641), .B(new_n697), .C1(new_n696), .C2(new_n721), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n681), .B(new_n694), .C1(new_n623), .C2(new_n625), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT111), .Z(new_n893));
  NOR2_X1   g707(.A1(new_n763), .A2(new_n692), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n893), .A2(new_n641), .A3(new_n706), .A4(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n890), .A2(new_n891), .A3(new_n770), .A4(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n698), .A2(new_n722), .A3(new_n770), .A4(new_n895), .ZN(new_n897));
  XNOR2_X1  g711(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n889), .A2(KEYINPUT53), .A3(new_n896), .A4(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n792), .A2(new_n874), .A3(new_n877), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n788), .B2(new_n783), .ZN(new_n902));
  INV_X1    g716(.A(new_n511), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n727), .A2(new_n903), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n795), .A2(new_n636), .A3(new_n638), .ZN(new_n905));
  AOI22_X1  g719(.A1(new_n904), .A2(new_n697), .B1(new_n513), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n631), .A3(new_n886), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n732), .A2(new_n737), .A3(new_n765), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n897), .A2(KEYINPUT52), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n902), .A2(new_n909), .A3(new_n896), .A4(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT53), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT54), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n900), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n889), .A2(KEYINPUT53), .A3(new_n896), .A4(new_n910), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n902), .A2(new_n909), .A3(new_n896), .A4(new_n899), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n912), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n914), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT113), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n917), .A2(new_n912), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n911), .A2(new_n912), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT54), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT113), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n900), .A2(new_n913), .A3(new_n914), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n872), .A2(new_n920), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT115), .ZN(new_n928));
  OR2_X1    g742(.A1(G952), .A2(G953), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n927), .A2(KEYINPUT115), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n838), .B1(new_n930), .B2(new_n931), .ZN(G75));
  NOR2_X1   g746(.A1(new_n347), .A2(G952), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n319), .B1(new_n900), .B2(new_n913), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT56), .B1(new_n935), .B2(G210), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n501), .A2(new_n503), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(new_n505), .Z(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT55), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n934), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n936), .B2(new_n940), .ZN(G51));
  NAND2_X1  g756(.A1(new_n900), .A2(new_n913), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT54), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n925), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n320), .B(KEYINPUT57), .Z(new_n947));
  OAI21_X1  g761(.A(new_n331), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n807), .A2(new_n808), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT116), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n935), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n933), .B1(new_n948), .B2(new_n951), .ZN(G54));
  NAND2_X1  g766(.A1(KEYINPUT58), .A2(G475), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT117), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n935), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n439), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n935), .A2(new_n436), .A3(new_n954), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n956), .A2(new_n934), .A3(new_n957), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT118), .Z(G60));
  NAND2_X1  g773(.A1(new_n645), .A2(new_n647), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n920), .A2(new_n926), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n649), .B(KEYINPUT59), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n960), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n962), .B1(new_n645), .B2(new_n647), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n933), .B1(new_n945), .B2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(KEYINPUT119), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT119), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n962), .B1(new_n920), .B2(new_n926), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n969), .B(new_n966), .C1(new_n970), .C2(new_n960), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n968), .A2(new_n971), .ZN(G63));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT60), .Z(new_n974));
  NAND2_X1  g788(.A1(new_n678), .A2(new_n679), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT120), .Z(new_n976));
  NAND3_X1  g790(.A1(new_n943), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n943), .A2(new_n974), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n934), .B(new_n977), .C1(new_n978), .C2(new_n619), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g794(.A(G953), .B1(new_n445), .B2(new_n453), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n909), .B2(G953), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n937), .B1(G898), .B2(new_n347), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(G69));
  INV_X1    g798(.A(new_n710), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n814), .B1(new_n653), .B2(new_n884), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n985), .B(new_n986), .C1(new_n629), .C2(new_n630), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n817), .A2(new_n826), .A3(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT62), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n890), .A2(new_n770), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(new_n713), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n990), .A2(new_n989), .A3(new_n713), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n988), .A2(KEYINPUT122), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT122), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n993), .A2(new_n817), .A3(new_n826), .A4(new_n987), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n995), .B1(new_n996), .B2(new_n991), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n347), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n431), .B(KEYINPUT121), .Z(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(new_n544), .Z(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n999), .A2(KEYINPUT123), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT123), .ZN(new_n1004));
  AOI21_X1  g818(.A(G953), .B1(new_n994), .B2(new_n997), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1004), .B1(new_n1005), .B2(new_n1001), .ZN(new_n1006));
  NAND2_X1  g820(.A1(G900), .A2(G953), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1001), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n813), .A2(new_n724), .A3(new_n709), .A4(new_n894), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n1009), .A2(KEYINPUT125), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1009), .A2(KEYINPUT125), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n817), .B(new_n826), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n990), .A2(new_n789), .A3(new_n792), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1008), .B1(new_n1014), .B2(new_n347), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1003), .A2(new_n1006), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(G900), .ZN(new_n1018));
  OAI21_X1  g832(.A(G953), .B1(new_n288), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT124), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1019), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1017), .B(new_n1021), .ZN(G72));
  NAND2_X1  g836(.A1(G472), .A2(G902), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT63), .Z(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1025), .B1(new_n1014), .B2(new_n909), .ZN(new_n1026));
  INV_X1    g840(.A(KEYINPUT126), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n547), .B(new_n702), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  NOR3_X1   g844(.A1(new_n998), .A2(new_n908), .A3(new_n907), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n703), .B1(new_n1031), .B2(new_n1025), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n916), .A2(new_n918), .ZN(new_n1033));
  INV_X1    g847(.A(new_n563), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT127), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1034), .B1(new_n582), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n581), .A2(KEYINPUT127), .A3(new_n547), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1025), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n933), .B1(new_n1033), .B2(new_n1038), .ZN(new_n1039));
  AND3_X1   g853(.A1(new_n1030), .A2(new_n1032), .A3(new_n1039), .ZN(G57));
endmodule


