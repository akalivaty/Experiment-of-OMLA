//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058;
  INV_X1    g000(.A(KEYINPUT78), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G140), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  AND2_X1   g003(.A1(new_n189), .A2(G227), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT73), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G131), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(KEYINPUT67), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G137), .ZN(new_n199));
  OR2_X1    g013(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n197), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n202), .A2(KEYINPUT66), .A3(KEYINPUT11), .A4(G134), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n198), .A2(G137), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n195), .B1(new_n201), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(G134), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n196), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n195), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n209), .A2(new_n210), .A3(new_n204), .A4(new_n203), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(KEYINPUT3), .A2(G107), .ZN(new_n213));
  NOR2_X1   g027(.A1(KEYINPUT3), .A2(G107), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n213), .B1(G104), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n216));
  INV_X1    g030(.A(G107), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT74), .ZN(new_n219));
  INV_X1    g033(.A(G104), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT74), .A2(G104), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G101), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n215), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n217), .A3(new_n222), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n224), .B1(G104), .B2(G107), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT64), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT64), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G146), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n231), .A2(new_n233), .A3(G143), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n230), .A2(G143), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(KEYINPUT1), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n234), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n237), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n230), .A2(G143), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n231), .A2(new_n233), .ZN(new_n243));
  INV_X1    g057(.A(G143), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n239), .B1(new_n240), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n229), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n225), .A2(new_n228), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n234), .A2(new_n236), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT76), .B1(new_n241), .B2(KEYINPUT1), .ZN(new_n250));
  OAI211_X1 g064(.A(KEYINPUT76), .B(KEYINPUT1), .C1(new_n244), .C2(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G128), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n249), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n248), .B1(new_n239), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n212), .B1(new_n247), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT12), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n252), .A2(new_n250), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT64), .B(G146), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n235), .B1(new_n259), .B2(G143), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n239), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n229), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n241), .B1(new_n259), .B2(G143), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n264), .B1(new_n259), .B2(G143), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n263), .B1(new_n265), .B2(new_n237), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n248), .A3(new_n239), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(KEYINPUT12), .A3(new_n212), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n257), .A2(new_n269), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n234), .A2(new_n236), .A3(new_n238), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G128), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n271), .B1(new_n273), .B2(new_n263), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT77), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n225), .A2(KEYINPUT10), .A3(new_n228), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n276), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT77), .B1(new_n278), .B2(new_n246), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n224), .A2(KEYINPUT75), .ZN(new_n281));
  INV_X1    g095(.A(new_n222), .ZN(new_n282));
  NOR2_X1   g096(.A1(KEYINPUT74), .A2(G104), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n282), .A2(new_n214), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(KEYINPUT3), .A2(G107), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n218), .B2(new_n220), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n281), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(KEYINPUT4), .A3(new_n225), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n215), .A2(new_n223), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT75), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT4), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .A4(G101), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g107(.A1(KEYINPUT0), .A2(G128), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n234), .A2(new_n236), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT65), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT65), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n234), .A2(new_n297), .A3(new_n236), .A4(new_n294), .ZN(new_n298));
  NOR2_X1   g112(.A1(KEYINPUT0), .A2(G128), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n296), .A2(new_n298), .B1(new_n263), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT10), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n293), .A2(new_n301), .B1(new_n302), .B2(new_n262), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n206), .A2(new_n211), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n280), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n193), .B1(new_n270), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n191), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n262), .A2(new_n302), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n275), .B1(new_n274), .B2(new_n276), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n296), .A2(new_n298), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n263), .A2(new_n300), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n310), .A2(new_n288), .A3(new_n292), .A4(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n278), .A2(KEYINPUT77), .A3(new_n246), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n308), .A2(new_n309), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n307), .B1(new_n314), .B2(new_n212), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n304), .B1(new_n280), .B2(new_n303), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n187), .B1(new_n306), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G902), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n314), .A2(new_n212), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n305), .A2(new_n320), .A3(new_n307), .ZN(new_n321));
  AND4_X1   g135(.A1(new_n308), .A2(new_n309), .A3(new_n312), .A4(new_n313), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n322), .A2(new_n304), .B1(new_n257), .B2(new_n269), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n321), .B(KEYINPUT78), .C1(new_n323), .C2(new_n193), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n318), .A2(new_n319), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G469), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT79), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT79), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(new_n328), .A3(G469), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT81), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n257), .A2(new_n330), .A3(new_n269), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT12), .B1(new_n268), .B2(new_n212), .ZN(new_n332));
  AOI211_X1 g146(.A(new_n256), .B(new_n304), .C1(new_n262), .C2(new_n267), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT81), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n331), .A2(new_n334), .A3(new_n305), .A4(new_n307), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n314), .A2(new_n212), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n191), .B1(new_n316), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT80), .B(G469), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n319), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n327), .A2(new_n329), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT9), .B(G234), .ZN(new_n343));
  OAI21_X1  g157(.A(G221), .B1(new_n343), .B2(G902), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n244), .A2(G128), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n237), .A2(G143), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(G134), .ZN(new_n349));
  XNOR2_X1  g163(.A(G116), .B(G122), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G107), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n217), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n349), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT13), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n346), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n244), .A2(KEYINPUT13), .A3(G128), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(new_n347), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n358), .A2(KEYINPUT91), .A3(G134), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT91), .B1(new_n358), .B2(G134), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n354), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n198), .B1(new_n346), .B2(new_n347), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n353), .B1(new_n349), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G116), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(KEYINPUT14), .A3(G122), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G107), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT14), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n366), .B1(new_n367), .B2(new_n350), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT92), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n348), .B(G134), .ZN(new_n370));
  OAI211_X1 g184(.A(G107), .B(new_n365), .C1(new_n351), .C2(KEYINPUT14), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT92), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .A4(new_n353), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n361), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G217), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n343), .A2(new_n375), .A3(G953), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n361), .A2(new_n369), .A3(new_n373), .A4(new_n376), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n319), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT93), .ZN(new_n382));
  INV_X1    g196(.A(G478), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT94), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(KEYINPUT15), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(KEYINPUT15), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n383), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT93), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n380), .A2(new_n389), .A3(new_n319), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n382), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(G234), .A2(G237), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(G952), .A3(new_n189), .ZN(new_n393));
  XOR2_X1   g207(.A(new_n393), .B(KEYINPUT95), .Z(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT21), .B(G898), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(G902), .A3(G953), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OR2_X1    g212(.A1(new_n381), .A2(new_n388), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n391), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G237), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n189), .A3(G214), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT86), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n244), .ZN(new_n404));
  NOR2_X1   g218(.A1(G237), .A2(G953), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n405), .B(G214), .C1(KEYINPUT86), .C2(G143), .ZN(new_n406));
  NAND2_X1  g220(.A1(KEYINPUT18), .A2(G131), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(new_n406), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(KEYINPUT18), .A3(G131), .ZN(new_n410));
  INV_X1    g224(.A(G140), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G125), .ZN(new_n412));
  INV_X1    g226(.A(G125), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G140), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT87), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G125), .B(G140), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT87), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n417), .A2(new_n419), .A3(G146), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n243), .A2(new_n415), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n408), .B(new_n410), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n417), .A2(new_n419), .A3(KEYINPUT19), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT19), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT88), .B1(new_n418), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n417), .A2(new_n419), .A3(KEYINPUT88), .A4(KEYINPUT19), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n243), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT16), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n411), .A3(G125), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n415), .B2(new_n429), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT71), .ZN(new_n432));
  INV_X1    g246(.A(new_n430), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(KEYINPUT71), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(G146), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n409), .A2(G131), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n404), .A2(new_n406), .A3(new_n194), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n422), .B1(new_n428), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT89), .ZN(new_n442));
  XNOR2_X1  g256(.A(G113), .B(G122), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(new_n220), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT89), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n446), .B(new_n422), .C1(new_n428), .C2(new_n440), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n442), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT90), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT71), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n418), .A2(KEYINPUT16), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n450), .B1(new_n451), .B2(new_n430), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n452), .A2(new_n230), .A3(new_n434), .ZN(new_n453));
  AOI21_X1  g267(.A(G146), .B1(new_n432), .B2(new_n435), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n449), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT17), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n437), .A2(new_n456), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n437), .A2(new_n438), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n457), .B1(new_n458), .B2(new_n456), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n230), .B1(new_n452), .B2(new_n434), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n436), .A3(KEYINPUT90), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n455), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n444), .A3(new_n422), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n448), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(G475), .A2(G902), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT20), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT20), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n464), .A2(new_n468), .A3(new_n465), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n462), .A2(new_n444), .A3(new_n422), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n444), .B1(new_n462), .B2(new_n422), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n319), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G475), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n400), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n345), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT29), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n405), .A2(G210), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n478), .B(KEYINPUT27), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT26), .B(G101), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n479), .B(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n209), .A2(new_n194), .A3(new_n204), .A4(new_n203), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n207), .A2(new_n204), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G131), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT68), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT68), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n483), .A2(new_n488), .A3(new_n485), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n489), .A3(new_n246), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n310), .A2(new_n212), .A3(new_n311), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(G116), .B(G119), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT2), .B(G113), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n495), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n493), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n492), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n486), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n301), .A2(new_n212), .B1(new_n501), .B2(new_n246), .ZN(new_n502));
  INV_X1    g316(.A(new_n499), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(KEYINPUT28), .A3(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n503), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT28), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n482), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n501), .A2(new_n246), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n491), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(new_n499), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n490), .A2(new_n513), .A3(new_n491), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n514), .B1(new_n513), .B2(new_n502), .ZN(new_n515));
  AOI211_X1 g329(.A(new_n481), .B(new_n512), .C1(new_n515), .C2(new_n499), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n477), .B1(new_n509), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT28), .B1(new_n502), .B2(new_n503), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n511), .A2(new_n499), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n507), .B1(new_n506), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT69), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n503), .B1(new_n491), .B2(new_n510), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n512), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT69), .B1(new_n524), .B2(new_n507), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n522), .A2(new_n525), .A3(KEYINPUT29), .A4(new_n481), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n517), .A2(new_n319), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(G472), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n490), .A2(new_n513), .A3(new_n491), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n513), .B1(new_n491), .B2(new_n510), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n499), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(new_n481), .A3(new_n506), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT31), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n512), .B1(new_n515), .B2(new_n499), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT31), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n535), .A3(new_n481), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n508), .A2(new_n500), .A3(new_n504), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n482), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n533), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(G472), .A2(G902), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT32), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n540), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n532), .A2(KEYINPUT31), .B1(new_n482), .B2(new_n537), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n544), .B1(new_n545), .B2(new_n536), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT32), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n528), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n375), .B1(G234), .B2(new_n319), .ZN(new_n549));
  INV_X1    g363(.A(G119), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT70), .B1(new_n550), .B2(G128), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT23), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(G128), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n237), .A2(G119), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT23), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(KEYINPUT70), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n552), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G110), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n554), .A2(new_n553), .ZN(new_n559));
  XOR2_X1   g373(.A(KEYINPUT24), .B(G110), .Z(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n562), .B1(new_n460), .B2(new_n436), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n421), .ZN(new_n565));
  OAI22_X1  g379(.A1(new_n557), .A2(G110), .B1(new_n559), .B2(new_n560), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n436), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT72), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT22), .B(G137), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n564), .A2(new_n567), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n571), .ZN(new_n573));
  INV_X1    g387(.A(new_n567), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n573), .B1(new_n574), .B2(new_n563), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT25), .B1(new_n576), .B2(new_n319), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT25), .ZN(new_n578));
  AOI211_X1 g392(.A(new_n578), .B(G902), .C1(new_n572), .C2(new_n575), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n549), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n549), .A2(G902), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n548), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n266), .A2(new_n413), .A3(new_n239), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n301), .B2(new_n413), .ZN(new_n587));
  INV_X1    g401(.A(G224), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(G953), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT7), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT85), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n587), .A2(KEYINPUT85), .A3(new_n591), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT82), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n493), .A2(KEYINPUT5), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT5), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(new_n550), .A3(G116), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(G113), .A3(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n229), .A2(new_n597), .A3(new_n498), .A4(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n288), .A2(new_n292), .A3(new_n499), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n498), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT82), .B1(new_n604), .B2(new_n248), .ZN(new_n605));
  XNOR2_X1  g419(.A(G110), .B(G122), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n602), .A2(new_n603), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(KEYINPUT8), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n604), .A2(new_n248), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n604), .A2(new_n248), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT7), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n590), .B(new_n586), .C1(new_n301), .C2(new_n413), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n607), .B(new_n611), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(G902), .B1(new_n596), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n606), .B(KEYINPUT83), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n618), .A2(KEYINPUT84), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT6), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n617), .A2(KEYINPUT6), .A3(new_n619), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n623), .A3(new_n607), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n587), .A2(new_n589), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n613), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(G210), .B1(G237), .B2(G902), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n616), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n628), .ZN(new_n630));
  INV_X1    g444(.A(new_n626), .ZN(new_n631));
  INV_X1    g445(.A(new_n607), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n621), .B2(new_n620), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n631), .B1(new_n633), .B2(new_n623), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n594), .A2(new_n595), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n319), .B1(new_n635), .B2(new_n614), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n630), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n629), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(G214), .B1(G237), .B2(G902), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n585), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n476), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G101), .ZN(G3));
  INV_X1    g457(.A(G472), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n539), .B2(new_n319), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n580), .A2(new_n583), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n645), .A2(new_n546), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n342), .A2(new_n647), .A3(new_n344), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT96), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n344), .ZN(new_n651));
  INV_X1    g465(.A(new_n341), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n326), .B2(KEYINPUT79), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n651), .B1(new_n653), .B2(new_n329), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(KEYINPUT96), .A3(new_n647), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n638), .A2(new_n398), .A3(new_n639), .ZN(new_n656));
  AOI22_X1  g470(.A1(new_n467), .A2(new_n469), .B1(G475), .B2(new_n473), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n382), .A2(new_n390), .ZN(new_n658));
  OAI21_X1  g472(.A(KEYINPUT33), .B1(new_n376), .B2(KEYINPUT97), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n380), .B(new_n659), .Z(new_n660));
  NOR2_X1   g474(.A1(new_n383), .A2(G902), .ZN(new_n661));
  AOI22_X1  g475(.A1(new_n658), .A2(new_n383), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n656), .A2(new_n657), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n650), .A2(new_n655), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT34), .B(G104), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G6));
  NAND2_X1  g480(.A1(new_n391), .A2(new_n399), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n470), .A2(new_n474), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n656), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n650), .A2(new_n655), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT35), .B(G107), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  NAND2_X1  g486(.A1(new_n564), .A2(new_n567), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n571), .A2(KEYINPUT36), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n581), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n580), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n638), .A2(new_n639), .A3(new_n677), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n678), .A2(new_n546), .A3(new_n645), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n476), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  INV_X1    g496(.A(new_n678), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n394), .B1(G900), .B2(new_n397), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n668), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n654), .A2(new_n548), .A3(new_n683), .A4(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT98), .B(G128), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G30));
  XNOR2_X1  g503(.A(new_n684), .B(KEYINPUT39), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  OR3_X1    g505(.A1(new_n345), .A2(KEYINPUT40), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(KEYINPUT40), .B1(new_n345), .B2(new_n691), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n638), .B(KEYINPUT38), .Z(new_n694));
  OR2_X1    g508(.A1(new_n534), .A2(new_n482), .ZN(new_n695));
  AOI21_X1  g509(.A(G902), .B1(new_n524), .B2(new_n482), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n644), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n541), .B2(new_n542), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n547), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n468), .B1(new_n464), .B2(new_n465), .ZN(new_n701));
  INV_X1    g515(.A(new_n465), .ZN(new_n702));
  AOI211_X1 g516(.A(KEYINPUT20), .B(new_n702), .C1(new_n448), .C2(new_n463), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n474), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n639), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n705), .B1(new_n391), .B2(new_n399), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NOR4_X1   g521(.A1(new_n694), .A2(new_n700), .A3(new_n677), .A4(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n692), .A2(new_n693), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G143), .ZN(G45));
  NOR3_X1   g524(.A1(new_n657), .A2(new_n662), .A3(new_n685), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n654), .A2(new_n548), .A3(new_n683), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G146), .ZN(G48));
  NAND2_X1  g527(.A1(new_n338), .A2(new_n319), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(G469), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(new_n584), .A3(new_n344), .A4(new_n341), .ZN(new_n716));
  AOI22_X1  g530(.A1(new_n527), .A2(G472), .B1(new_n546), .B2(KEYINPUT32), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n716), .B1(new_n717), .B2(new_n543), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n663), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT99), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n718), .A2(KEYINPUT99), .A3(new_n663), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT41), .B(G113), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  AND3_X1   g539(.A1(new_n715), .A2(new_n344), .A3(new_n341), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n669), .A2(new_n548), .A3(new_n584), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G116), .ZN(G18));
  INV_X1    g542(.A(new_n475), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n548), .A2(new_n683), .A3(new_n726), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  AOI21_X1  g545(.A(new_n481), .B1(new_n522), .B2(new_n525), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n535), .B1(new_n534), .B2(new_n481), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT100), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n521), .B(KEYINPUT28), .C1(new_n512), .C2(new_n523), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n508), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n520), .A2(new_n521), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n482), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT100), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n739), .A3(new_n533), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n734), .A2(new_n536), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n645), .B1(new_n741), .B2(new_n540), .ZN(new_n742));
  AND4_X1   g556(.A1(new_n344), .A2(new_n715), .A3(new_n341), .A4(new_n398), .ZN(new_n743));
  INV_X1    g557(.A(new_n638), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n707), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n742), .A2(new_n743), .A3(new_n584), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  NAND2_X1  g561(.A1(new_n715), .A2(new_n341), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n748), .A2(new_n640), .A3(new_n651), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(new_n742), .A3(new_n677), .A4(new_n711), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  OAI21_X1  g565(.A(KEYINPUT104), .B1(new_n546), .B2(KEYINPUT32), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n541), .A2(new_n753), .A3(new_n542), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n752), .A2(new_n754), .A3(new_n528), .A4(new_n547), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n755), .A2(new_n584), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT101), .B1(new_n323), .B2(new_n193), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT101), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n332), .A2(new_n333), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n758), .B(new_n192), .C1(new_n336), .C2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n757), .A2(G469), .A3(new_n321), .A4(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(G469), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n319), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n341), .A2(new_n761), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT102), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(G902), .B1(new_n335), .B2(new_n337), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n763), .B1(new_n768), .B2(new_n340), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(KEYINPUT102), .A3(new_n761), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n629), .A2(new_n637), .A3(new_n344), .A4(new_n639), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT103), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT103), .ZN(new_n775));
  AOI211_X1 g589(.A(new_n775), .B(new_n772), .C1(new_n767), .C2(new_n770), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n756), .B(new_n711), .C1(new_n774), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n765), .A2(new_n766), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT102), .B1(new_n769), .B2(new_n761), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n773), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n775), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n771), .A2(KEYINPUT103), .A3(new_n773), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n585), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR4_X1   g597(.A1(new_n657), .A2(new_n662), .A3(KEYINPUT42), .A4(new_n685), .ZN(new_n784));
  AOI22_X1  g598(.A1(KEYINPUT42), .A2(new_n777), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G131), .ZN(G33));
  INV_X1    g600(.A(new_n585), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n787), .B(new_n686), .C1(new_n774), .C2(new_n776), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G134), .ZN(G36));
  NOR2_X1   g603(.A1(new_n638), .A2(new_n705), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n645), .A2(new_n546), .ZN(new_n792));
  INV_X1    g606(.A(new_n677), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n660), .A2(new_n661), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n382), .A2(new_n390), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n795), .B1(new_n796), .B2(G478), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT43), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n657), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT43), .B1(new_n662), .B2(new_n704), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT105), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n801), .B1(new_n799), .B2(new_n800), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n794), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT44), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n791), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT106), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n807), .B1(new_n804), .B2(new_n805), .ZN(new_n808));
  INV_X1    g622(.A(new_n803), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(KEYINPUT106), .A3(KEYINPUT44), .A4(new_n794), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n806), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT107), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT45), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n318), .A2(new_n816), .A3(new_n324), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n757), .A2(new_n321), .A3(new_n760), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n817), .B(G469), .C1(new_n816), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n764), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT46), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n652), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(KEYINPUT46), .A3(new_n764), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n344), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n691), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n806), .A2(new_n808), .A3(new_n812), .A4(KEYINPUT107), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n815), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G137), .ZN(G39));
  XNOR2_X1  g643(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n825), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n824), .A2(new_n344), .A3(new_n830), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n711), .A2(new_n646), .A3(new_n790), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n548), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(G140), .ZN(G42));
  NAND2_X1  g652(.A1(new_n742), .A2(new_n584), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n394), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n799), .A2(new_n800), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n790), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT113), .Z(new_n846));
  INV_X1    g660(.A(new_n748), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n834), .B1(new_n651), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n748), .A2(new_n394), .A3(new_n772), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n700), .A2(new_n584), .A3(new_n851), .ZN(new_n852));
  XOR2_X1   g666(.A(new_n852), .B(KEYINPUT115), .Z(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n657), .A3(new_n662), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT114), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n694), .A2(new_n705), .A3(new_n726), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n855), .B1(new_n843), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT50), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n851), .A2(new_n800), .A3(new_n799), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n677), .A3(new_n742), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n854), .A2(new_n859), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  OR3_X1    g677(.A1(new_n849), .A2(new_n850), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n850), .B1(new_n849), .B2(new_n863), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n853), .A2(new_n704), .A3(new_n797), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n189), .A2(G952), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n844), .B2(new_n749), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n866), .A2(KEYINPUT116), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT116), .B1(new_n866), .B2(new_n868), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n861), .A2(new_n756), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT48), .Z(new_n872));
  NOR3_X1   g686(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n864), .A2(new_n865), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n777), .A2(KEYINPUT42), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n783), .A2(new_n784), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n391), .A2(KEYINPUT109), .A3(new_n399), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT109), .B1(new_n391), .B2(new_n399), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n657), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(new_n657), .B2(new_n797), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n656), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n650), .A2(new_n883), .A3(new_n655), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n654), .B(new_n729), .C1(new_n641), .C2(new_n679), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n875), .A2(new_n876), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n742), .A2(new_n677), .A3(new_n711), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n781), .A2(new_n782), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n654), .A2(new_n548), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT109), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n667), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n657), .A2(new_n684), .A3(new_n877), .A4(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT110), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n880), .A2(KEYINPUT110), .A3(new_n657), .A4(new_n684), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n793), .A2(new_n638), .A3(new_n705), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n887), .A2(new_n888), .B1(new_n889), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n746), .A2(new_n727), .A3(new_n730), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n721), .B2(new_n722), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n898), .A2(new_n900), .A3(new_n788), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n886), .A2(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n687), .A2(new_n750), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT52), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n685), .A2(new_n651), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n638), .A2(new_n704), .A3(new_n706), .A4(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n767), .B2(new_n770), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n677), .B1(new_n698), .B2(new_n547), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT112), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n907), .A2(KEYINPUT112), .A3(new_n908), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n903), .A2(new_n904), .A3(new_n712), .A4(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n687), .A2(new_n712), .A3(new_n750), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n907), .A2(KEYINPUT112), .A3(new_n908), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT112), .B1(new_n907), .B2(new_n908), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT52), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n687), .A2(new_n750), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT52), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n902), .A2(new_n920), .A3(KEYINPUT53), .A4(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT54), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT53), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n884), .A2(new_n885), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n887), .B1(new_n774), .B2(new_n776), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n897), .A2(new_n654), .A3(new_n548), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n788), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n926), .A2(new_n785), .A3(new_n929), .A4(new_n900), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n914), .A2(new_n919), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n925), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n923), .A2(new_n924), .A3(new_n932), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n930), .A2(new_n931), .A3(new_n925), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT111), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n886), .B2(new_n901), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n788), .A2(new_n928), .A3(new_n927), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n727), .A2(new_n730), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n718), .A2(KEYINPUT99), .A3(new_n663), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT99), .B1(new_n718), .B2(new_n663), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n938), .B(new_n746), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n942), .A2(KEYINPUT111), .A3(new_n785), .A4(new_n926), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n914), .A2(new_n919), .A3(new_n922), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n936), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n934), .B1(new_n945), .B2(new_n925), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n933), .B1(new_n946), .B2(new_n924), .ZN(new_n947));
  OAI22_X1  g761(.A1(new_n874), .A2(new_n947), .B1(G952), .B2(G953), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n748), .B(KEYINPUT49), .Z(new_n949));
  NAND3_X1  g763(.A1(new_n584), .A2(new_n344), .A3(new_n639), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n950), .A2(new_n704), .A3(new_n662), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n949), .A2(new_n694), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n948), .B1(new_n699), .B2(new_n952), .ZN(G75));
  NOR2_X1   g767(.A1(new_n189), .A2(G952), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n319), .B1(new_n923), .B2(new_n932), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT56), .B1(new_n956), .B2(G210), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n624), .A2(new_n626), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n958), .A2(new_n634), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT55), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n955), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(new_n957), .B2(new_n960), .ZN(G51));
  AOI211_X1 g776(.A(new_n319), .B(new_n819), .C1(new_n923), .C2(new_n932), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n763), .B(KEYINPUT57), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n923), .A2(new_n924), .A3(new_n932), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n924), .B1(new_n923), .B2(new_n932), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n963), .B1(new_n967), .B2(new_n338), .ZN(new_n968));
  OAI21_X1  g782(.A(KEYINPUT117), .B1(new_n968), .B2(new_n954), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT117), .ZN(new_n970));
  INV_X1    g784(.A(new_n338), .ZN(new_n971));
  INV_X1    g785(.A(new_n922), .ZN(new_n972));
  NOR4_X1   g786(.A1(new_n930), .A2(new_n931), .A3(new_n925), .A4(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(KEYINPUT53), .B1(new_n902), .B2(new_n920), .ZN(new_n974));
  OAI21_X1  g788(.A(KEYINPUT54), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n933), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n971), .B1(new_n976), .B2(new_n964), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n970), .B(new_n955), .C1(new_n977), .C2(new_n963), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n969), .A2(new_n978), .ZN(G54));
  AND2_X1   g793(.A1(KEYINPUT58), .A2(G475), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n956), .A2(new_n464), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n464), .B1(new_n956), .B2(new_n980), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n981), .A2(new_n982), .A3(new_n954), .ZN(G60));
  XOR2_X1   g797(.A(new_n660), .B(KEYINPUT118), .Z(new_n984));
  NAND2_X1  g798(.A1(G478), .A2(G902), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT59), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n954), .B1(new_n976), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n984), .B1(new_n947), .B2(new_n986), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n988), .B1(new_n989), .B2(KEYINPUT119), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT119), .ZN(new_n991));
  AOI211_X1 g805(.A(new_n991), .B(new_n984), .C1(new_n947), .C2(new_n986), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n990), .A2(new_n992), .ZN(G63));
  NAND2_X1  g807(.A1(G217), .A2(G902), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT120), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT60), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n973), .B2(new_n974), .ZN(new_n997));
  INV_X1    g811(.A(new_n576), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n675), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n999), .B(new_n955), .C1(new_n1000), .C2(new_n997), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT61), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(G66));
  OAI21_X1  g817(.A(G953), .B1(new_n395), .B2(new_n588), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n926), .A2(new_n900), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1004), .B1(new_n1006), .B2(G953), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n633), .B(new_n623), .C1(G898), .C2(new_n189), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT121), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1007), .B(new_n1009), .ZN(G69));
  AOI21_X1  g824(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n654), .A2(new_n690), .ZN(new_n1013));
  NOR4_X1   g827(.A1(new_n1013), .A2(new_n585), .A3(new_n791), .A4(new_n882), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1014), .B1(new_n834), .B2(new_n836), .ZN(new_n1015));
  INV_X1    g829(.A(new_n915), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT62), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n709), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(KEYINPUT122), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT122), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n709), .A2(new_n1016), .A3(new_n1020), .A4(new_n1017), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n828), .A2(new_n1015), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n709), .A2(new_n1016), .ZN(new_n1023));
  AND3_X1   g837(.A1(new_n1023), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n1024));
  AOI21_X1  g838(.A(KEYINPUT123), .B1(new_n1023), .B2(KEYINPUT62), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n189), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n426), .A2(new_n427), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n515), .B(new_n1028), .Z(new_n1029));
  INV_X1    g843(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g845(.A(KEYINPUT124), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n826), .A2(new_n745), .A3(new_n756), .ZN(new_n1033));
  AND3_X1   g847(.A1(new_n1033), .A2(new_n785), .A3(new_n788), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n915), .B1(new_n834), .B2(new_n836), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1034), .A2(new_n828), .A3(new_n189), .A4(new_n1035), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1030), .B1(G900), .B2(G953), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1031), .A2(new_n1032), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g853(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1032), .B1(new_n1031), .B2(new_n1038), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1012), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1031), .A2(new_n1038), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(KEYINPUT124), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1044), .A2(new_n1011), .A3(new_n1039), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1042), .A2(new_n1045), .ZN(G72));
  OR3_X1    g860(.A1(new_n1022), .A2(new_n1026), .A3(new_n1005), .ZN(new_n1047));
  NAND2_X1  g861(.A1(G472), .A2(G902), .ZN(new_n1048));
  XNOR2_X1  g862(.A(new_n1048), .B(KEYINPUT126), .ZN(new_n1049));
  XOR2_X1   g863(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1050));
  XNOR2_X1  g864(.A(new_n1049), .B(new_n1050), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n695), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g866(.A1(new_n1034), .A2(new_n828), .A3(new_n1035), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1051), .B1(new_n1053), .B2(new_n1005), .ZN(new_n1054));
  AND2_X1   g868(.A1(new_n1054), .A2(new_n516), .ZN(new_n1055));
  INV_X1    g869(.A(new_n516), .ZN(new_n1056));
  NAND3_X1  g870(.A1(new_n695), .A2(new_n1056), .A3(new_n1051), .ZN(new_n1057));
  NOR2_X1   g871(.A1(new_n946), .A2(new_n1057), .ZN(new_n1058));
  NOR4_X1   g872(.A1(new_n1052), .A2(new_n954), .A3(new_n1055), .A4(new_n1058), .ZN(G57));
endmodule


