

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780;

  BUF_X1 U375 ( .A(n665), .Z(n423) );
  NAND2_X1 U376 ( .A1(n734), .A2(n512), .ZN(n364) );
  INV_X1 U377 ( .A(G902), .ZN(n496) );
  XNOR2_X1 U378 ( .A(G116), .B(G113), .ZN(n531) );
  BUF_X1 U379 ( .A(G143), .Z(n720) );
  XNOR2_X1 U380 ( .A(n479), .B(n480), .ZN(n482) );
  XOR2_X2 U381 ( .A(KEYINPUT59), .B(n727), .Z(n728) );
  XNOR2_X2 U382 ( .A(n415), .B(n741), .ZN(n743) );
  AND2_X2 U383 ( .A1(n418), .A2(n694), .ZN(n416) );
  NAND2_X2 U384 ( .A1(n416), .A2(G472), .ZN(n697) );
  XNOR2_X2 U385 ( .A(n353), .B(KEYINPUT86), .ZN(n687) );
  NAND2_X1 U386 ( .A1(n686), .A2(n689), .ZN(n353) );
  XOR2_X2 U387 ( .A(n473), .B(KEYINPUT95), .Z(n381) );
  INV_X2 U388 ( .A(KEYINPUT0), .ZN(n646) );
  NOR2_X1 U389 ( .A1(n730), .A2(n745), .ZN(n732) );
  AND2_X2 U390 ( .A1(n390), .A2(n652), .ZN(n659) );
  NAND2_X1 U391 ( .A1(G237), .A2(G234), .ZN(n565) );
  XNOR2_X1 U392 ( .A(G146), .B(G125), .ZN(n481) );
  XOR2_X1 U393 ( .A(G122), .B(G134), .Z(n488) );
  XNOR2_X2 U394 ( .A(n419), .B(n646), .ZN(n649) );
  XNOR2_X2 U395 ( .A(G122), .B(G113), .ZN(n398) );
  INV_X16 U396 ( .A(G953), .ZN(n774) );
  XNOR2_X1 U397 ( .A(n670), .B(KEYINPUT32), .ZN(n719) );
  XNOR2_X1 U398 ( .A(n398), .B(G104), .ZN(n478) );
  NAND2_X1 U399 ( .A1(n512), .A2(G902), .ZN(n363) );
  INV_X1 U400 ( .A(G116), .ZN(n466) );
  INV_X1 U401 ( .A(G902), .ZN(n361) );
  INV_X1 U402 ( .A(KEYINPUT67), .ZN(n370) );
  INV_X1 U403 ( .A(KEYINPUT100), .ZN(n374) );
  XNOR2_X1 U404 ( .A(n677), .B(n676), .ZN(n679) );
  NAND2_X1 U405 ( .A1(n434), .A2(n719), .ZN(n672) );
  XNOR2_X1 U406 ( .A(n671), .B(n370), .ZN(n369) );
  NAND2_X1 U407 ( .A1(n452), .A2(n383), .ZN(n451) );
  XNOR2_X1 U408 ( .A(n602), .B(n424), .ZN(n452) );
  INV_X2 U409 ( .A(n750), .ZN(n395) );
  OR2_X2 U410 ( .A1(n362), .A2(n359), .ZN(n414) );
  NAND2_X1 U411 ( .A1(n364), .A2(n363), .ZN(n362) );
  XNOR2_X1 U412 ( .A(n476), .B(n421), .ZN(n420) );
  NAND2_X1 U413 ( .A1(G469), .A2(n361), .ZN(n360) );
  NOR2_X1 U414 ( .A1(n453), .A2(G953), .ZN(n486) );
  XNOR2_X1 U415 ( .A(G119), .B(G140), .ZN(n518) );
  INV_X1 U416 ( .A(G237), .ZN(n472) );
  XNOR2_X1 U417 ( .A(KEYINPUT71), .B(KEYINPUT3), .ZN(n465) );
  INV_X1 U418 ( .A(G234), .ZN(n453) );
  XNOR2_X1 U419 ( .A(G107), .B(G104), .ZN(n510) );
  XNOR2_X1 U420 ( .A(KEYINPUT75), .B(KEYINPUT34), .ZN(n648) );
  INV_X1 U421 ( .A(KEYINPUT81), .ZN(n676) );
  XNOR2_X2 U422 ( .A(n356), .B(n386), .ZN(n712) );
  NAND2_X1 U423 ( .A1(n649), .A2(n373), .ZN(n356) );
  NAND2_X1 U424 ( .A1(n357), .A2(n436), .ZN(n435) );
  NAND2_X1 U425 ( .A1(n722), .A2(KEYINPUT44), .ZN(n357) );
  XNOR2_X1 U426 ( .A(n358), .B(KEYINPUT69), .ZN(n625) );
  NAND2_X1 U427 ( .A1(n615), .A2(n616), .ZN(n358) );
  XNOR2_X1 U428 ( .A(n366), .B(KEYINPUT45), .ZN(n686) );
  NAND2_X1 U429 ( .A1(n663), .A2(n662), .ZN(n434) );
  OR2_X2 U430 ( .A1(n734), .A2(G902), .ZN(n365) );
  NOR2_X1 U431 ( .A1(n734), .A2(n360), .ZN(n359) );
  XNOR2_X1 U432 ( .A(n365), .B(G469), .ZN(n593) );
  NOR2_X1 U433 ( .A1(n746), .A2(n745), .ZN(n748) );
  NOR2_X1 U434 ( .A1(n703), .A2(n745), .ZN(n705) );
  NAND2_X1 U435 ( .A1(n371), .A2(n367), .ZN(n366) );
  NAND2_X1 U436 ( .A1(n369), .A2(n368), .ZN(n367) );
  INV_X1 U437 ( .A(n672), .ZN(n368) );
  XNOR2_X1 U438 ( .A(n372), .B(n454), .ZN(n371) );
  NAND2_X1 U439 ( .A1(n437), .A2(n438), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n560), .B(n559), .ZN(n621) );
  XNOR2_X2 U441 ( .A(n545), .B(n374), .ZN(n373) );
  INV_X1 U442 ( .A(n373), .ZN(n650) );
  BUF_X1 U443 ( .A(n591), .Z(n375) );
  BUF_X1 U444 ( .A(n701), .Z(n376) );
  NAND2_X2 U445 ( .A1(n586), .A2(n608), .ZN(n439) );
  XNOR2_X1 U446 ( .A(n607), .B(KEYINPUT38), .ZN(n377) );
  XNOR2_X1 U447 ( .A(n607), .B(KEYINPUT38), .ZN(n617) );
  BUF_X1 U448 ( .A(n508), .Z(n378) );
  BUF_X1 U449 ( .A(n696), .Z(n379) );
  XNOR2_X2 U450 ( .A(n380), .B(n381), .ZN(n586) );
  NOR2_X2 U451 ( .A1(n742), .A2(n689), .ZN(n380) );
  XNOR2_X1 U452 ( .A(n391), .B(n399), .ZN(n616) );
  INV_X1 U453 ( .A(KEYINPUT77), .ZN(n399) );
  NAND2_X1 U454 ( .A1(n392), .A2(n400), .ZN(n391) );
  XNOR2_X1 U455 ( .A(n393), .B(n401), .ZN(n392) );
  XNOR2_X1 U456 ( .A(n481), .B(KEYINPUT10), .ZN(n514) );
  NOR2_X2 U457 ( .A1(G953), .A2(G237), .ZN(n534) );
  INV_X1 U458 ( .A(KEYINPUT70), .ZN(n441) );
  XNOR2_X1 U459 ( .A(n623), .B(n388), .ZN(n624) );
  XNOR2_X1 U460 ( .A(G137), .B(G134), .ZN(n507) );
  NAND2_X1 U461 ( .A1(n593), .A2(n592), .ZN(n447) );
  XNOR2_X1 U462 ( .A(n419), .B(n646), .ZN(n413) );
  XNOR2_X1 U463 ( .A(n420), .B(n475), .ZN(n480) );
  XNOR2_X1 U464 ( .A(n510), .B(n511), .ZN(n450) );
  XNOR2_X1 U465 ( .A(n426), .B(n619), .ZN(n639) );
  INV_X1 U466 ( .A(KEYINPUT112), .ZN(n443) );
  XOR2_X1 U467 ( .A(n440), .B(G472), .Z(n410) );
  INV_X1 U468 ( .A(KEYINPUT78), .ZN(n401) );
  XNOR2_X1 U469 ( .A(G131), .B(KEYINPUT5), .ZN(n530) );
  INV_X1 U470 ( .A(KEYINPUT11), .ZN(n421) );
  XOR2_X1 U471 ( .A(KEYINPUT103), .B(KEYINPUT12), .Z(n475) );
  XNOR2_X1 U472 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n459) );
  OR2_X2 U473 ( .A1(n617), .A2(n597), .ZN(n397) );
  XNOR2_X1 U474 ( .A(n447), .B(n446), .ZN(n595) );
  INV_X1 U475 ( .A(KEYINPUT108), .ZN(n446) );
  XNOR2_X1 U476 ( .A(n579), .B(KEYINPUT6), .ZN(n666) );
  NOR2_X1 U477 ( .A1(n629), .A2(n395), .ZN(n630) );
  NOR2_X1 U478 ( .A1(n634), .A2(n395), .ZN(n609) );
  XNOR2_X1 U479 ( .A(n483), .B(KEYINPUT13), .ZN(n484) );
  INV_X1 U480 ( .A(G475), .ZN(n483) );
  NAND2_X1 U481 ( .A1(n445), .A2(n410), .ZN(n651) );
  BUF_X1 U482 ( .A(n666), .Z(n422) );
  XNOR2_X1 U483 ( .A(KEYINPUT76), .B(KEYINPUT16), .ZN(n467) );
  XNOR2_X1 U484 ( .A(n514), .B(n513), .ZN(n405) );
  XNOR2_X1 U485 ( .A(KEYINPUT98), .B(KEYINPUT80), .ZN(n513) );
  XNOR2_X1 U486 ( .A(n450), .B(n509), .ZN(n449) );
  NOR2_X1 U487 ( .A1(n774), .A2(G952), .ZN(n745) );
  INV_X1 U488 ( .A(n639), .ZN(n394) );
  AND2_X2 U489 ( .A1(n587), .A2(n417), .ZN(n400) );
  INV_X1 U490 ( .A(KEYINPUT110), .ZN(n424) );
  NAND2_X1 U491 ( .A1(n407), .A2(n607), .ZN(n602) );
  AND2_X1 U492 ( .A1(n400), .A2(n396), .ZN(n382) );
  AND2_X1 U493 ( .A1(n604), .A2(n603), .ZN(n383) );
  AND2_X1 U494 ( .A1(n654), .A2(n653), .ZN(n384) );
  AND2_X1 U495 ( .A1(n658), .A2(n422), .ZN(n385) );
  XNOR2_X1 U496 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n386) );
  AND2_X1 U497 ( .A1(n400), .A2(n750), .ZN(n387) );
  XOR2_X1 U498 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n388) );
  XOR2_X1 U499 ( .A(n379), .B(n695), .Z(n389) );
  NAND2_X1 U500 ( .A1(n712), .A2(n749), .ZN(n390) );
  NAND2_X1 U501 ( .A1(n652), .A2(n572), .ZN(n393) );
  NAND2_X1 U502 ( .A1(n638), .A2(n395), .ZN(n503) );
  NAND2_X1 U503 ( .A1(n394), .A2(n750), .ZN(n620) );
  NOR2_X1 U504 ( .A1(n712), .A2(n395), .ZN(n713) );
  AND2_X2 U505 ( .A1(n604), .A2(n501), .ZN(n750) );
  INV_X1 U506 ( .A(n757), .ZN(n396) );
  NAND2_X1 U507 ( .A1(n558), .A2(n654), .ZN(n560) );
  XNOR2_X2 U508 ( .A(n397), .B(KEYINPUT113), .ZN(n558) );
  NAND2_X1 U509 ( .A1(n402), .A2(n423), .ZN(n661) );
  NAND2_X1 U510 ( .A1(n402), .A2(n669), .ZN(n670) );
  AND2_X1 U511 ( .A1(n402), .A2(n385), .ZN(n709) );
  XNOR2_X2 U512 ( .A(n412), .B(n656), .ZN(n402) );
  XNOR2_X1 U513 ( .A(n403), .B(G128), .ZN(n519) );
  XNOR2_X2 U514 ( .A(G110), .B(KEYINPUT24), .ZN(n403) );
  XNOR2_X2 U515 ( .A(n404), .B(n525), .ZN(n591) );
  OR2_X2 U516 ( .A1(n701), .A2(G902), .ZN(n404) );
  XNOR2_X1 U517 ( .A(n406), .B(n405), .ZN(n701) );
  XNOR2_X1 U518 ( .A(n521), .B(n516), .ZN(n406) );
  NAND2_X1 U519 ( .A1(n407), .A2(n618), .ZN(n426) );
  AND2_X2 U520 ( .A1(n601), .A2(n600), .ZN(n407) );
  XNOR2_X2 U521 ( .A(n425), .B(n448), .ZN(n734) );
  XNOR2_X2 U522 ( .A(n408), .B(n443), .ZN(n587) );
  NAND2_X1 U523 ( .A1(n585), .A2(n584), .ZN(n408) );
  XNOR2_X1 U524 ( .A(n430), .B(KEYINPUT35), .ZN(n409) );
  XNOR2_X1 U525 ( .A(n430), .B(KEYINPUT35), .ZN(n722) );
  NAND2_X2 U526 ( .A1(n431), .A2(n383), .ZN(n430) );
  BUF_X1 U527 ( .A(n717), .Z(n411) );
  NAND2_X1 U528 ( .A1(n413), .A2(n384), .ZN(n412) );
  NAND2_X2 U529 ( .A1(n433), .A2(n456), .ZN(n419) );
  BUF_X1 U530 ( .A(n742), .Z(n415) );
  AND2_X2 U531 ( .A1(n418), .A2(n694), .ZN(n738) );
  BUF_X1 U532 ( .A(n433), .Z(n417) );
  NAND2_X1 U533 ( .A1(n692), .A2(n455), .ZN(n418) );
  NAND2_X1 U534 ( .A1(n649), .A2(n647), .ZN(n432) );
  XNOR2_X1 U535 ( .A(n427), .B(n378), .ZN(n464) );
  XNOR2_X1 U536 ( .A(n432), .B(n648), .ZN(n431) );
  INV_X1 U537 ( .A(n413), .ZN(n655) );
  XNOR2_X1 U538 ( .A(n485), .B(n484), .ZN(n500) );
  BUF_X2 U539 ( .A(n586), .Z(n607) );
  OR2_X2 U540 ( .A1(n696), .A2(G902), .ZN(n440) );
  XNOR2_X1 U541 ( .A(n425), .B(n540), .ZN(n696) );
  XNOR2_X2 U542 ( .A(n772), .B(G146), .ZN(n425) );
  XNOR2_X1 U543 ( .A(n427), .B(n449), .ZN(n448) );
  XNOR2_X2 U544 ( .A(n428), .B(n536), .ZN(n427) );
  XNOR2_X2 U545 ( .A(KEYINPUT66), .B(G101), .ZN(n536) );
  XNOR2_X2 U546 ( .A(n429), .B(KEYINPUT72), .ZN(n428) );
  XNOR2_X2 U547 ( .A(G110), .B(KEYINPUT73), .ZN(n429) );
  XNOR2_X2 U548 ( .A(n439), .B(KEYINPUT19), .ZN(n433) );
  XNOR2_X1 U549 ( .A(n434), .B(G110), .ZN(G12) );
  XNOR2_X1 U550 ( .A(n435), .B(KEYINPUT91), .ZN(n437) );
  NOR2_X2 U551 ( .A1(n659), .A2(n709), .ZN(n436) );
  NAND2_X1 U552 ( .A1(n672), .A2(KEYINPUT44), .ZN(n438) );
  XNOR2_X2 U553 ( .A(n440), .B(G472), .ZN(n579) );
  XNOR2_X2 U554 ( .A(n442), .B(n441), .ZN(n581) );
  NAND2_X1 U555 ( .A1(n591), .A2(n578), .ZN(n442) );
  NAND2_X1 U556 ( .A1(n444), .A2(n587), .ZN(n622) );
  INV_X1 U557 ( .A(n621), .ZN(n444) );
  INV_X1 U558 ( .A(n447), .ZN(n445) );
  XNOR2_X2 U559 ( .A(n508), .B(n507), .ZN(n772) );
  XNOR2_X2 U560 ( .A(n489), .B(n458), .ZN(n508) );
  NAND2_X1 U561 ( .A1(n451), .A2(n605), .ZN(n606) );
  XNOR2_X1 U562 ( .A(n451), .B(n721), .ZN(G45) );
  INV_X1 U563 ( .A(KEYINPUT90), .ZN(n454) );
  XNOR2_X1 U564 ( .A(n697), .B(n389), .ZN(n699) );
  NAND2_X1 U565 ( .A1(n640), .A2(n707), .ZN(n773) );
  XNOR2_X2 U566 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n458) );
  OR2_X1 U567 ( .A1(n691), .A2(n690), .ZN(n455) );
  OR2_X1 U568 ( .A1(n645), .A2(n644), .ZN(n456) );
  NOR2_X1 U569 ( .A1(n665), .A2(n546), .ZN(n457) );
  INV_X1 U570 ( .A(n410), .ZN(n580) );
  BUF_X1 U571 ( .A(n489), .Z(n491) );
  NAND2_X1 U572 ( .A1(n581), .A2(n579), .ZN(n583) );
  INV_X1 U573 ( .A(KEYINPUT22), .ZN(n656) );
  INV_X1 U574 ( .A(n745), .ZN(n698) );
  INV_X1 U575 ( .A(KEYINPUT127), .ZN(n704) );
  XNOR2_X1 U576 ( .A(n685), .B(n684), .ZN(G75) );
  XNOR2_X2 U577 ( .A(G128), .B(G143), .ZN(n489) );
  XNOR2_X1 U578 ( .A(n481), .B(n459), .ZN(n462) );
  NAND2_X1 U579 ( .A1(n774), .A2(G224), .ZN(n460) );
  XNOR2_X1 U580 ( .A(n460), .B(KEYINPUT94), .ZN(n461) );
  XNOR2_X1 U581 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U582 ( .A(n464), .B(n463), .ZN(n471) );
  XNOR2_X1 U583 ( .A(n465), .B(G119), .ZN(n533) );
  XNOR2_X1 U584 ( .A(n533), .B(n478), .ZN(n470) );
  XNOR2_X1 U585 ( .A(n466), .B(G107), .ZN(n490) );
  INV_X1 U586 ( .A(n490), .ZN(n468) );
  XNOR2_X1 U587 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U588 ( .A(n470), .B(n469), .ZN(n765) );
  XNOR2_X1 U589 ( .A(n471), .B(n765), .ZN(n742) );
  XNOR2_X2 U590 ( .A(KEYINPUT15), .B(G902), .ZN(n522) );
  INV_X1 U591 ( .A(n522), .ZN(n689) );
  NAND2_X1 U592 ( .A1(n496), .A2(n472), .ZN(n474) );
  NAND2_X1 U593 ( .A1(n474), .A2(G210), .ZN(n473) );
  AND2_X1 U594 ( .A1(n474), .A2(G214), .ZN(n597) );
  NAND2_X1 U595 ( .A1(n377), .A2(n597), .ZN(n499) );
  NAND2_X1 U596 ( .A1(n534), .A2(G214), .ZN(n476) );
  XNOR2_X1 U597 ( .A(n720), .B(KEYINPUT102), .ZN(n477) );
  XNOR2_X1 U598 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X2 U599 ( .A(G140), .B(G131), .ZN(n511) );
  XNOR2_X1 U600 ( .A(n514), .B(n511), .ZN(n771) );
  XNOR2_X1 U601 ( .A(n482), .B(n771), .ZN(n727) );
  NOR2_X1 U602 ( .A1(G902), .A2(n727), .ZN(n485) );
  XNOR2_X1 U603 ( .A(KEYINPUT8), .B(n486), .ZN(n515) );
  NAND2_X1 U604 ( .A1(G217), .A2(n515), .ZN(n487) );
  XNOR2_X1 U605 ( .A(n488), .B(n487), .ZN(n495) );
  XNOR2_X1 U606 ( .A(n491), .B(n490), .ZN(n493) );
  XOR2_X1 U607 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n492) );
  XNOR2_X1 U608 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U609 ( .A(n495), .B(n494), .ZN(n723) );
  NAND2_X1 U610 ( .A1(n723), .A2(n496), .ZN(n498) );
  INV_X1 U611 ( .A(G478), .ZN(n497) );
  XNOR2_X1 U612 ( .A(n498), .B(n497), .ZN(n501) );
  AND2_X1 U613 ( .A1(n500), .A2(n501), .ZN(n654) );
  NAND2_X1 U614 ( .A1(n499), .A2(n654), .ZN(n505) );
  INV_X1 U615 ( .A(n501), .ZN(n603) );
  NAND2_X1 U616 ( .A1(n500), .A2(n603), .ZN(n757) );
  XNOR2_X1 U617 ( .A(n757), .B(KEYINPUT104), .ZN(n638) );
  INV_X1 U618 ( .A(n500), .ZN(n604) );
  INV_X1 U619 ( .A(KEYINPUT105), .ZN(n502) );
  XNOR2_X2 U620 ( .A(n503), .B(n502), .ZN(n588) );
  NAND2_X1 U621 ( .A1(n558), .A2(n588), .ZN(n504) );
  NAND2_X1 U622 ( .A1(n505), .A2(n504), .ZN(n506) );
  XOR2_X1 U623 ( .A(KEYINPUT123), .B(n506), .Z(n544) );
  NAND2_X1 U624 ( .A1(n774), .A2(G227), .ZN(n509) );
  INV_X1 U625 ( .A(G469), .ZN(n512) );
  XNOR2_X2 U626 ( .A(n414), .B(KEYINPUT1), .ZN(n665) );
  INV_X1 U627 ( .A(n665), .ZN(n657) );
  NAND2_X1 U628 ( .A1(n515), .A2(G221), .ZN(n516) );
  XNOR2_X2 U629 ( .A(G137), .B(KEYINPUT23), .ZN(n517) );
  XNOR2_X1 U630 ( .A(n518), .B(n517), .ZN(n520) );
  XNOR2_X1 U631 ( .A(n520), .B(n519), .ZN(n521) );
  NAND2_X1 U632 ( .A1(n522), .A2(G234), .ZN(n523) );
  XNOR2_X1 U633 ( .A(n523), .B(KEYINPUT20), .ZN(n526) );
  NAND2_X1 U634 ( .A1(n526), .A2(G217), .ZN(n524) );
  XNOR2_X1 U635 ( .A(n524), .B(KEYINPUT25), .ZN(n525) );
  INV_X1 U636 ( .A(n526), .ZN(n528) );
  INV_X1 U637 ( .A(G221), .ZN(n527) );
  OR2_X1 U638 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U639 ( .A(n529), .B(KEYINPUT21), .ZN(n590) );
  OR2_X1 U640 ( .A1(n591), .A2(n590), .ZN(n546) );
  XNOR2_X1 U641 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U642 ( .A(n533), .B(n532), .ZN(n539) );
  NAND2_X1 U643 ( .A1(n534), .A2(G210), .ZN(n535) );
  XNOR2_X1 U644 ( .A(n535), .B(KEYINPUT99), .ZN(n537) );
  XNOR2_X1 U645 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U646 ( .A(n539), .B(n538), .ZN(n540) );
  NOR2_X1 U647 ( .A1(n546), .A2(n666), .ZN(n541) );
  NAND2_X1 U648 ( .A1(n657), .A2(n541), .ZN(n543) );
  XNOR2_X1 U649 ( .A(KEYINPUT74), .B(KEYINPUT33), .ZN(n542) );
  XNOR2_X1 U650 ( .A(n543), .B(n542), .ZN(n647) );
  BUF_X1 U651 ( .A(n647), .Z(n569) );
  NAND2_X1 U652 ( .A1(n544), .A2(n569), .ZN(n563) );
  NAND2_X1 U653 ( .A1(n457), .A2(n579), .ZN(n545) );
  INV_X1 U654 ( .A(n546), .ZN(n548) );
  NAND2_X1 U655 ( .A1(n423), .A2(n546), .ZN(n547) );
  NAND2_X1 U656 ( .A1(n547), .A2(KEYINPUT50), .ZN(n551) );
  NOR2_X1 U657 ( .A1(n548), .A2(KEYINPUT50), .ZN(n549) );
  NAND2_X1 U658 ( .A1(n423), .A2(n549), .ZN(n550) );
  NAND2_X1 U659 ( .A1(n551), .A2(n550), .ZN(n555) );
  INV_X1 U660 ( .A(n375), .ZN(n664) );
  NAND2_X1 U661 ( .A1(n375), .A2(n590), .ZN(n552) );
  XNOR2_X1 U662 ( .A(n552), .B(KEYINPUT49), .ZN(n553) );
  NOR2_X1 U663 ( .A1(n580), .A2(n553), .ZN(n554) );
  NAND2_X1 U664 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U665 ( .A1(n650), .A2(n556), .ZN(n557) );
  XOR2_X1 U666 ( .A(KEYINPUT51), .B(n557), .Z(n561) );
  INV_X1 U667 ( .A(KEYINPUT41), .ZN(n559) );
  NAND2_X1 U668 ( .A1(n561), .A2(n444), .ZN(n562) );
  NAND2_X1 U669 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U670 ( .A(n564), .B(KEYINPUT52), .ZN(n567) );
  XNOR2_X1 U671 ( .A(n565), .B(KEYINPUT14), .ZN(n574) );
  NAND2_X1 U672 ( .A1(G952), .A2(n574), .ZN(n566) );
  XOR2_X1 U673 ( .A(KEYINPUT96), .B(n566), .Z(n573) );
  NAND2_X1 U674 ( .A1(n567), .A2(n573), .ZN(n568) );
  XNOR2_X1 U675 ( .A(n568), .B(KEYINPUT124), .ZN(n571) );
  NAND2_X1 U676 ( .A1(n444), .A2(n569), .ZN(n570) );
  NAND2_X1 U677 ( .A1(n571), .A2(n570), .ZN(n682) );
  XNOR2_X1 U678 ( .A(n588), .B(KEYINPUT84), .ZN(n652) );
  INV_X1 U679 ( .A(KEYINPUT47), .ZN(n572) );
  AND2_X1 U680 ( .A1(n573), .A2(n774), .ZN(n645) );
  INV_X1 U681 ( .A(n645), .ZN(n577) );
  NAND2_X1 U682 ( .A1(G902), .A2(n574), .ZN(n641) );
  NOR2_X1 U683 ( .A1(G900), .A2(n641), .ZN(n575) );
  NAND2_X1 U684 ( .A1(n575), .A2(G953), .ZN(n576) );
  NAND2_X1 U685 ( .A1(n577), .A2(n576), .ZN(n594) );
  INV_X1 U686 ( .A(n590), .ZN(n653) );
  AND2_X1 U687 ( .A1(n594), .A2(n653), .ZN(n578) );
  INV_X1 U688 ( .A(KEYINPUT28), .ZN(n582) );
  XNOR2_X1 U689 ( .A(n583), .B(n582), .ZN(n585) );
  XNOR2_X1 U690 ( .A(n414), .B(KEYINPUT111), .ZN(n584) );
  INV_X1 U691 ( .A(n597), .ZN(n608) );
  NAND2_X1 U692 ( .A1(n400), .A2(n588), .ZN(n589) );
  NAND2_X1 U693 ( .A1(n589), .A2(KEYINPUT47), .ZN(n605) );
  NOR2_X1 U694 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U695 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U696 ( .A(n596), .B(KEYINPUT79), .ZN(n601) );
  OR2_X1 U697 ( .A1(n410), .A2(n597), .ZN(n599) );
  XNOR2_X1 U698 ( .A(KEYINPUT109), .B(KEYINPUT30), .ZN(n598) );
  XNOR2_X1 U699 ( .A(n599), .B(n598), .ZN(n600) );
  XNOR2_X1 U700 ( .A(n606), .B(KEYINPUT83), .ZN(n614) );
  INV_X1 U701 ( .A(n607), .ZN(n634) );
  AND2_X1 U702 ( .A1(n581), .A2(n608), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n609), .A2(n628), .ZN(n610) );
  NOR2_X1 U704 ( .A1(n610), .A2(n422), .ZN(n611) );
  XNOR2_X1 U705 ( .A(n611), .B(KEYINPUT36), .ZN(n612) );
  NAND2_X1 U706 ( .A1(n612), .A2(n657), .ZN(n613) );
  XNOR2_X1 U707 ( .A(n613), .B(KEYINPUT114), .ZN(n716) );
  AND2_X1 U708 ( .A1(n614), .A2(n716), .ZN(n615) );
  INV_X1 U709 ( .A(n377), .ZN(n618) );
  INV_X1 U710 ( .A(KEYINPUT39), .ZN(n619) );
  XNOR2_X1 U711 ( .A(n620), .B(KEYINPUT40), .ZN(n718) );
  XNOR2_X1 U712 ( .A(n622), .B(KEYINPUT42), .ZN(n717) );
  NAND2_X1 U713 ( .A1(n718), .A2(n717), .ZN(n623) );
  NAND2_X1 U714 ( .A1(n624), .A2(n625), .ZN(n627) );
  INV_X1 U715 ( .A(KEYINPUT48), .ZN(n626) );
  XNOR2_X1 U716 ( .A(n627), .B(n626), .ZN(n636) );
  INV_X1 U717 ( .A(n628), .ZN(n629) );
  NAND2_X1 U718 ( .A1(n630), .A2(n423), .ZN(n631) );
  OR2_X1 U719 ( .A1(n631), .A2(n422), .ZN(n633) );
  XOR2_X1 U720 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n632) );
  XNOR2_X1 U721 ( .A(n633), .B(n632), .ZN(n635) );
  NAND2_X1 U722 ( .A1(n635), .A2(n634), .ZN(n706) );
  NAND2_X1 U723 ( .A1(n636), .A2(n706), .ZN(n637) );
  XNOR2_X1 U724 ( .A(n637), .B(KEYINPUT89), .ZN(n640) );
  OR2_X1 U725 ( .A1(n639), .A2(n638), .ZN(n707) );
  INV_X1 U726 ( .A(n773), .ZN(n674) );
  INV_X1 U727 ( .A(n641), .ZN(n642) );
  NOR2_X1 U728 ( .A1(G898), .A2(n774), .ZN(n767) );
  NAND2_X1 U729 ( .A1(n642), .A2(n767), .ZN(n643) );
  XNOR2_X1 U730 ( .A(n643), .B(KEYINPUT97), .ZN(n644) );
  OR2_X1 U731 ( .A1(n655), .A2(n651), .ZN(n749) );
  NOR2_X1 U732 ( .A1(n657), .A2(n375), .ZN(n658) );
  INV_X1 U733 ( .A(KEYINPUT106), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n661), .B(n660), .ZN(n663) );
  AND2_X1 U735 ( .A1(n410), .A2(n375), .ZN(n662) );
  OR2_X1 U736 ( .A1(n423), .A2(n664), .ZN(n668) );
  INV_X1 U737 ( .A(n422), .ZN(n667) );
  NOR2_X1 U738 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U739 ( .A1(n409), .A2(KEYINPUT44), .ZN(n671) );
  BUF_X1 U740 ( .A(n686), .Z(n673) );
  NAND2_X1 U741 ( .A1(n674), .A2(n673), .ZN(n678) );
  INV_X1 U742 ( .A(KEYINPUT2), .ZN(n690) );
  XNOR2_X1 U743 ( .A(KEYINPUT82), .B(n690), .ZN(n675) );
  NAND2_X1 U744 ( .A1(n678), .A2(n675), .ZN(n677) );
  NOR2_X1 U745 ( .A1(n678), .A2(n690), .ZN(n693) );
  NAND2_X1 U746 ( .A1(n679), .A2(n694), .ZN(n680) );
  XNOR2_X1 U747 ( .A(n680), .B(KEYINPUT87), .ZN(n681) );
  NOR2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U749 ( .A1(n683), .A2(n774), .ZN(n685) );
  INV_X1 U750 ( .A(KEYINPUT53), .ZN(n684) );
  NOR2_X2 U751 ( .A1(n687), .A2(n773), .ZN(n688) );
  XNOR2_X1 U752 ( .A(n688), .B(KEYINPUT85), .ZN(n692) );
  XOR2_X1 U753 ( .A(KEYINPUT88), .B(n689), .Z(n691) );
  INV_X1 U754 ( .A(n693), .ZN(n694) );
  XOR2_X1 U755 ( .A(KEYINPUT115), .B(KEYINPUT62), .Z(n695) );
  NAND2_X1 U756 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U757 ( .A(n700), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U758 ( .A1(n738), .A2(G217), .ZN(n702) );
  XNOR2_X1 U759 ( .A(n702), .B(n376), .ZN(n703) );
  XNOR2_X1 U760 ( .A(n705), .B(n704), .ZN(G66) );
  XNOR2_X1 U761 ( .A(n706), .B(G140), .ZN(G42) );
  XNOR2_X1 U762 ( .A(n707), .B(G134), .ZN(G36) );
  XOR2_X1 U763 ( .A(G101), .B(KEYINPUT116), .Z(n708) );
  XNOR2_X1 U764 ( .A(n709), .B(n708), .ZN(G3) );
  XOR2_X1 U765 ( .A(G146), .B(n387), .Z(G48) );
  XOR2_X1 U766 ( .A(G116), .B(KEYINPUT121), .Z(n711) );
  NOR2_X1 U767 ( .A1(n757), .A2(n712), .ZN(n710) );
  XOR2_X1 U768 ( .A(n711), .B(n710), .Z(G18) );
  XOR2_X1 U769 ( .A(G113), .B(n713), .Z(G15) );
  XOR2_X1 U770 ( .A(KEYINPUT37), .B(KEYINPUT122), .Z(n714) );
  XNOR2_X1 U771 ( .A(n714), .B(G125), .ZN(n715) );
  XNOR2_X1 U772 ( .A(n716), .B(n715), .ZN(G27) );
  XNOR2_X1 U773 ( .A(n411), .B(G137), .ZN(G39) );
  XNOR2_X1 U774 ( .A(n718), .B(G131), .ZN(G33) );
  XNOR2_X1 U775 ( .A(n719), .B(G119), .ZN(G21) );
  XNOR2_X1 U776 ( .A(n720), .B(KEYINPUT120), .ZN(n721) );
  XOR2_X1 U777 ( .A(n409), .B(G122), .Z(G24) );
  NAND2_X1 U778 ( .A1(n416), .A2(G478), .ZN(n725) );
  XOR2_X1 U779 ( .A(KEYINPUT126), .B(n723), .Z(n724) );
  XNOR2_X1 U780 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X1 U781 ( .A1(n726), .A2(n745), .ZN(G63) );
  NAND2_X1 U782 ( .A1(n738), .A2(G475), .ZN(n729) );
  XNOR2_X1 U783 ( .A(n729), .B(n728), .ZN(n730) );
  XOR2_X1 U784 ( .A(KEYINPUT65), .B(KEYINPUT60), .Z(n731) );
  XNOR2_X1 U785 ( .A(n732), .B(n731), .ZN(G60) );
  NAND2_X1 U786 ( .A1(n416), .A2(G469), .ZN(n736) );
  XOR2_X1 U787 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n733) );
  XNOR2_X1 U788 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U789 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U790 ( .A1(n737), .A2(n745), .ZN(G54) );
  NAND2_X1 U791 ( .A1(n738), .A2(G210), .ZN(n744) );
  XNOR2_X1 U792 ( .A(KEYINPUT93), .B(KEYINPUT54), .ZN(n740) );
  XNOR2_X1 U793 ( .A(KEYINPUT55), .B(KEYINPUT92), .ZN(n739) );
  XNOR2_X1 U794 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U795 ( .A(n744), .B(n743), .ZN(n746) );
  XOR2_X1 U796 ( .A(KEYINPUT125), .B(KEYINPUT56), .Z(n747) );
  XNOR2_X1 U797 ( .A(n748), .B(n747), .ZN(G51) );
  INV_X1 U798 ( .A(n749), .ZN(n752) );
  NAND2_X1 U799 ( .A1(n752), .A2(n750), .ZN(n751) );
  XNOR2_X1 U800 ( .A(n751), .B(G104), .ZN(G6) );
  XOR2_X1 U801 ( .A(KEYINPUT26), .B(KEYINPUT117), .Z(n754) );
  NAND2_X1 U802 ( .A1(n752), .A2(n396), .ZN(n753) );
  XNOR2_X1 U803 ( .A(n754), .B(n753), .ZN(n756) );
  XOR2_X1 U804 ( .A(G107), .B(KEYINPUT27), .Z(n755) );
  XNOR2_X1 U805 ( .A(n756), .B(n755), .ZN(G9) );
  XOR2_X1 U806 ( .A(KEYINPUT29), .B(KEYINPUT119), .Z(n758) );
  XOR2_X1 U807 ( .A(n758), .B(n382), .Z(n760) );
  XOR2_X1 U808 ( .A(G128), .B(KEYINPUT118), .Z(n759) );
  XNOR2_X1 U809 ( .A(n760), .B(n759), .ZN(G30) );
  NAND2_X1 U810 ( .A1(n673), .A2(n774), .ZN(n764) );
  NAND2_X1 U811 ( .A1(G953), .A2(G224), .ZN(n761) );
  XNOR2_X1 U812 ( .A(KEYINPUT61), .B(n761), .ZN(n762) );
  NAND2_X1 U813 ( .A1(n762), .A2(G898), .ZN(n763) );
  NAND2_X1 U814 ( .A1(n764), .A2(n763), .ZN(n770) );
  XNOR2_X1 U815 ( .A(G110), .B(G101), .ZN(n766) );
  XOR2_X1 U816 ( .A(n766), .B(n765), .Z(n768) );
  NOR2_X1 U817 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U818 ( .A(n770), .B(n769), .ZN(G69) );
  XOR2_X1 U819 ( .A(n772), .B(n771), .Z(n776) );
  XNOR2_X1 U820 ( .A(n773), .B(n776), .ZN(n775) );
  NAND2_X1 U821 ( .A1(n775), .A2(n774), .ZN(n780) );
  XNOR2_X1 U822 ( .A(n776), .B(G227), .ZN(n777) );
  NAND2_X1 U823 ( .A1(n777), .A2(G900), .ZN(n778) );
  NAND2_X1 U824 ( .A1(n778), .A2(G953), .ZN(n779) );
  NAND2_X1 U825 ( .A1(n780), .A2(n779), .ZN(G72) );
endmodule

