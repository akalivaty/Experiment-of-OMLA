

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780;

  NAND2_X2 U368 ( .A1(n369), .A2(n368), .ZN(n489) );
  XNOR2_X1 U369 ( .A(n391), .B(KEYINPUT102), .ZN(n778) );
  NAND2_X1 U370 ( .A1(n559), .A2(n558), .ZN(n445) );
  XNOR2_X1 U371 ( .A(n548), .B(KEYINPUT100), .ZN(n485) );
  NAND2_X1 U372 ( .A1(n623), .A2(n553), .ZN(n548) );
  AND2_X1 U373 ( .A1(n701), .A2(n702), .ZN(n553) );
  OR2_X1 U374 ( .A1(n738), .A2(n431), .ZN(n430) );
  INV_X1 U375 ( .A(G146), .ZN(n447) );
  XNOR2_X1 U376 ( .A(n552), .B(n551), .ZN(n691) );
  NOR2_X1 U377 ( .A1(n442), .A2(n605), .ZN(n621) );
  XNOR2_X1 U378 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X2 U379 ( .A1(n395), .A2(n394), .ZN(n623) );
  INV_X1 U380 ( .A(n686), .ZN(n442) );
  NAND2_X1 U381 ( .A1(n428), .A2(KEYINPUT1), .ZN(n394) );
  NAND2_X1 U382 ( .A1(n432), .A2(n430), .ZN(n428) );
  AND2_X1 U383 ( .A1(n434), .A2(n433), .ZN(n432) );
  XNOR2_X1 U384 ( .A(n465), .B(n464), .ZN(n701) );
  XNOR2_X1 U385 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U386 ( .A(n491), .B(G137), .ZN(n466) );
  XNOR2_X2 U387 ( .A(n606), .B(KEYINPUT19), .ZN(n425) );
  XNOR2_X2 U388 ( .A(n346), .B(KEYINPUT81), .ZN(n606) );
  NAND2_X1 U389 ( .A1(n505), .A2(n714), .ZN(n346) );
  XNOR2_X2 U390 ( .A(n398), .B(n351), .ZN(n505) );
  AND2_X1 U391 ( .A1(n779), .A2(n545), .ZN(n374) );
  XNOR2_X1 U392 ( .A(n544), .B(n543), .ZN(n347) );
  XNOR2_X1 U393 ( .A(n544), .B(n543), .ZN(n378) );
  BUF_X1 U394 ( .A(n363), .Z(n348) );
  NAND2_X1 U395 ( .A1(n636), .A2(n635), .ZN(n349) );
  XNOR2_X1 U396 ( .A(n547), .B(KEYINPUT32), .ZN(n350) );
  NAND2_X1 U397 ( .A1(n636), .A2(n635), .ZN(n638) );
  XNOR2_X1 U398 ( .A(n547), .B(KEYINPUT32), .ZN(n779) );
  NAND2_X2 U399 ( .A1(n696), .A2(KEYINPUT2), .ZN(n635) );
  XNOR2_X2 U400 ( .A(n349), .B(n637), .ZN(n364) );
  XNOR2_X2 U401 ( .A(n638), .B(n637), .ZN(n363) );
  XNOR2_X1 U402 ( .A(n450), .B(KEYINPUT20), .ZN(n461) );
  NOR2_X1 U403 ( .A1(n717), .A2(n415), .ZN(n414) );
  INV_X1 U404 ( .A(n717), .ZN(n411) );
  XNOR2_X1 U405 ( .A(n526), .B(n525), .ZN(n649) );
  XNOR2_X1 U406 ( .A(n766), .B(n518), .ZN(n526) );
  XNOR2_X1 U407 ( .A(n524), .B(n523), .ZN(n525) );
  NOR2_X1 U408 ( .A1(n683), .A2(n444), .ZN(n614) );
  NAND2_X1 U409 ( .A1(n618), .A2(KEYINPUT67), .ZN(n387) );
  XNOR2_X1 U410 ( .A(n375), .B(KEYINPUT99), .ZN(n565) );
  NAND2_X1 U411 ( .A1(n376), .A2(n561), .ZN(n375) );
  OR2_X1 U412 ( .A1(n691), .A2(n676), .ZN(n376) );
  INV_X1 U413 ( .A(G131), .ZN(n473) );
  NAND2_X1 U414 ( .A1(n381), .A2(n380), .ZN(n408) );
  AND2_X1 U415 ( .A1(n778), .A2(n436), .ZN(n380) );
  NOR2_X1 U416 ( .A1(n437), .A2(n620), .ZN(n407) );
  XNOR2_X1 U417 ( .A(n463), .B(n462), .ZN(n464) );
  OR2_X1 U418 ( .A1(n639), .A2(G902), .ZN(n465) );
  XNOR2_X1 U419 ( .A(n493), .B(n446), .ZN(n515) );
  INV_X1 U420 ( .A(KEYINPUT10), .ZN(n446) );
  XNOR2_X1 U421 ( .A(n455), .B(n453), .ZN(n401) );
  XNOR2_X1 U422 ( .A(G110), .B(G140), .ZN(n455) );
  XNOR2_X1 U423 ( .A(G122), .B(KEYINPUT7), .ZN(n531) );
  XOR2_X1 U424 ( .A(KEYINPUT97), .B(KEYINPUT9), .Z(n532) );
  XNOR2_X1 U425 ( .A(n534), .B(n533), .ZN(n535) );
  INV_X1 U426 ( .A(KEYINPUT96), .ZN(n533) );
  XNOR2_X1 U427 ( .A(G107), .B(G116), .ZN(n534) );
  XNOR2_X1 U428 ( .A(KEYINPUT77), .B(KEYINPUT8), .ZN(n456) );
  NAND2_X1 U429 ( .A1(n410), .A2(n417), .ZN(n409) );
  AND2_X1 U430 ( .A1(n416), .A2(n413), .ZN(n412) );
  NOR2_X1 U431 ( .A1(n590), .A2(n589), .ZN(n613) );
  XNOR2_X1 U432 ( .A(n529), .B(n528), .ZN(n559) );
  BUF_X1 U433 ( .A(n768), .Z(n403) );
  NOR2_X1 U434 ( .A1(n355), .A2(n423), .ZN(n422) );
  NAND2_X1 U435 ( .A1(n443), .A2(n442), .ZN(n599) );
  NOR2_X1 U436 ( .A1(n690), .A2(n444), .ZN(n443) );
  NOR2_X1 U437 ( .A1(n383), .A2(n385), .ZN(n382) );
  NAND2_X1 U438 ( .A1(n387), .A2(n384), .ZN(n383) );
  INV_X1 U439 ( .A(n620), .ZN(n384) );
  XNOR2_X1 U440 ( .A(KEYINPUT48), .B(KEYINPUT79), .ZN(n620) );
  XNOR2_X1 U441 ( .A(G116), .B(G113), .ZN(n426) );
  NOR2_X1 U442 ( .A1(G237), .A2(G953), .ZN(n479) );
  XNOR2_X1 U443 ( .A(G140), .B(G131), .ZN(n468) );
  INV_X1 U444 ( .A(G237), .ZN(n502) );
  XNOR2_X1 U445 ( .A(n449), .B(n527), .ZN(n629) );
  XNOR2_X1 U446 ( .A(KEYINPUT85), .B(KEYINPUT15), .ZN(n449) );
  NOR2_X1 U447 ( .A1(n701), .A2(n440), .ZN(n603) );
  NAND2_X1 U448 ( .A1(n702), .A2(n441), .ZN(n440) );
  INV_X1 U449 ( .A(n585), .ZN(n441) );
  XNOR2_X1 U450 ( .A(n569), .B(n568), .ZN(n632) );
  XNOR2_X1 U451 ( .A(G113), .B(G122), .ZN(n516) );
  XNOR2_X1 U452 ( .A(G104), .B(G143), .ZN(n519) );
  XOR2_X1 U453 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n520) );
  XNOR2_X1 U454 ( .A(n515), .B(n468), .ZN(n766) );
  XOR2_X1 U455 ( .A(KEYINPUT18), .B(KEYINPUT73), .Z(n496) );
  XNOR2_X1 U456 ( .A(n581), .B(KEYINPUT38), .ZN(n715) );
  INV_X1 U457 ( .A(G902), .ZN(n527) );
  OR2_X1 U458 ( .A1(n353), .A2(G902), .ZN(n431) );
  NAND2_X1 U459 ( .A1(n353), .A2(G902), .ZN(n433) );
  NAND2_X1 U460 ( .A1(n461), .A2(G221), .ZN(n393) );
  INV_X1 U461 ( .A(n559), .ZN(n418) );
  XNOR2_X1 U462 ( .A(n483), .B(n482), .ZN(n664) );
  XNOR2_X1 U463 ( .A(n481), .B(KEYINPUT5), .ZN(n482) );
  NAND2_X1 U464 ( .A1(n406), .A2(n405), .ZN(n767) );
  NOR2_X1 U465 ( .A1(n408), .A2(n407), .ZN(n406) );
  NAND2_X1 U466 ( .A1(n386), .A2(n359), .ZN(n438) );
  XNOR2_X1 U467 ( .A(n397), .B(n396), .ZN(n758) );
  INV_X1 U468 ( .A(G107), .ZN(n396) );
  XNOR2_X1 U469 ( .A(G110), .B(G104), .ZN(n397) );
  XNOR2_X1 U470 ( .A(KEYINPUT16), .B(G122), .ZN(n488) );
  BUF_X1 U471 ( .A(n632), .Z(n750) );
  INV_X1 U472 ( .A(n562), .ZN(n423) );
  XNOR2_X1 U473 ( .A(n454), .B(n401), .ZN(n459) );
  XNOR2_X1 U474 ( .A(n404), .B(n356), .ZN(n538) );
  XNOR2_X1 U475 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U476 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U477 ( .A(n643), .B(n642), .ZN(n745) );
  XNOR2_X1 U478 ( .A(n421), .B(n419), .ZN(n776) );
  XNOR2_X1 U479 ( .A(n420), .B(KEYINPUT42), .ZN(n419) );
  INV_X1 U480 ( .A(KEYINPUT106), .ZN(n420) );
  INV_X1 U481 ( .A(KEYINPUT35), .ZN(n377) );
  AND2_X1 U482 ( .A1(n546), .A2(n562), .ZN(n424) );
  AND2_X1 U483 ( .A1(n613), .A2(n392), .ZN(n683) );
  INV_X1 U484 ( .A(n545), .ZN(n647) );
  XOR2_X1 U485 ( .A(n503), .B(KEYINPUT86), .Z(n351) );
  XNOR2_X1 U486 ( .A(n393), .B(n354), .ZN(n584) );
  INV_X1 U487 ( .A(n584), .ZN(n702) );
  AND2_X1 U488 ( .A1(n545), .A2(KEYINPUT44), .ZN(n352) );
  XNOR2_X1 U489 ( .A(KEYINPUT68), .B(G469), .ZN(n353) );
  XOR2_X1 U490 ( .A(KEYINPUT91), .B(KEYINPUT21), .Z(n354) );
  OR2_X1 U491 ( .A1(n623), .A2(n705), .ZN(n355) );
  XOR2_X1 U492 ( .A(n536), .B(n535), .Z(n356) );
  AND2_X1 U493 ( .A1(n350), .A2(n352), .ZN(n357) );
  AND2_X1 U494 ( .A1(n430), .A2(n429), .ZN(n358) );
  AND2_X1 U495 ( .A1(n388), .A2(n387), .ZN(n359) );
  NOR2_X1 U496 ( .A1(n690), .A2(n686), .ZN(n360) );
  INV_X1 U497 ( .A(KEYINPUT1), .ZN(n429) );
  XNOR2_X1 U498 ( .A(n379), .B(G122), .ZN(G24) );
  NAND2_X1 U499 ( .A1(n558), .A2(n418), .ZN(n717) );
  INV_X1 U500 ( .A(n558), .ZN(n541) );
  XNOR2_X1 U501 ( .A(n402), .B(G478), .ZN(n558) );
  INV_X1 U502 ( .A(n514), .ZN(n361) );
  XNOR2_X2 U503 ( .A(n487), .B(n486), .ZN(n730) );
  BUF_X1 U504 ( .A(n350), .Z(n362) );
  BUF_X1 U505 ( .A(n489), .Z(n365) );
  XNOR2_X1 U506 ( .A(n478), .B(G119), .ZN(n427) );
  NAND2_X1 U507 ( .A1(n427), .A2(n426), .ZN(n368) );
  NAND2_X1 U508 ( .A1(n366), .A2(n367), .ZN(n369) );
  INV_X1 U509 ( .A(n427), .ZN(n366) );
  INV_X1 U510 ( .A(n426), .ZN(n367) );
  BUF_X1 U511 ( .A(n425), .Z(n370) );
  NOR2_X1 U512 ( .A1(n565), .A2(n646), .ZN(n566) );
  NAND2_X1 U513 ( .A1(n371), .A2(n448), .ZN(n373) );
  NAND2_X1 U514 ( .A1(n374), .A2(n379), .ZN(n371) );
  NAND2_X1 U515 ( .A1(n373), .A2(n372), .ZN(n567) );
  NAND2_X1 U516 ( .A1(n379), .A2(n357), .ZN(n372) );
  XNOR2_X2 U517 ( .A(n540), .B(n377), .ZN(n379) );
  NAND2_X1 U518 ( .A1(n347), .A2(n422), .ZN(n545) );
  NAND2_X1 U519 ( .A1(n378), .A2(n424), .ZN(n547) );
  AND2_X1 U520 ( .A1(n347), .A2(n564), .ZN(n646) );
  NAND2_X1 U521 ( .A1(n382), .A2(n386), .ZN(n381) );
  NAND2_X1 U522 ( .A1(n390), .A2(n389), .ZN(n386) );
  INV_X1 U523 ( .A(n388), .ZN(n385) );
  NAND2_X1 U524 ( .A1(n619), .A2(KEYINPUT67), .ZN(n388) );
  NAND2_X1 U525 ( .A1(n626), .A2(n581), .ZN(n391) );
  INV_X1 U526 ( .A(n619), .ZN(n389) );
  NOR2_X1 U527 ( .A1(n618), .A2(KEYINPUT67), .ZN(n390) );
  INV_X1 U528 ( .A(n370), .ZN(n392) );
  INV_X1 U529 ( .A(n553), .ZN(n698) );
  NAND2_X1 U530 ( .A1(n358), .A2(n432), .ZN(n395) );
  INV_X1 U531 ( .A(n505), .ZN(n581) );
  NAND2_X1 U532 ( .A1(n655), .A2(n629), .ZN(n398) );
  XNOR2_X1 U533 ( .A(n501), .B(n500), .ZN(n655) );
  AND2_X2 U534 ( .A1(n634), .A2(n633), .ZN(n696) );
  NAND2_X1 U535 ( .A1(n399), .A2(n631), .ZN(n636) );
  NAND2_X1 U536 ( .A1(n628), .A2(n627), .ZN(n399) );
  XNOR2_X1 U537 ( .A(n400), .B(KEYINPUT34), .ZN(n539) );
  NOR2_X2 U538 ( .A1(n514), .A2(n730), .ZN(n400) );
  NOR2_X1 U539 ( .A1(n746), .A2(G902), .ZN(n402) );
  NAND2_X1 U540 ( .A1(n537), .A2(G217), .ZN(n404) );
  NAND2_X1 U541 ( .A1(n435), .A2(n438), .ZN(n405) );
  NAND2_X1 U542 ( .A1(n715), .A2(n714), .ZN(n719) );
  NAND2_X1 U543 ( .A1(n412), .A2(n409), .ZN(n729) );
  NAND2_X1 U544 ( .A1(n411), .A2(n714), .ZN(n410) );
  NAND2_X1 U545 ( .A1(n414), .A2(n715), .ZN(n413) );
  NAND2_X1 U546 ( .A1(n714), .A2(KEYINPUT41), .ZN(n415) );
  OR2_X1 U547 ( .A1(n715), .A2(KEYINPUT41), .ZN(n416) );
  INV_X1 U548 ( .A(KEYINPUT41), .ZN(n417) );
  NOR2_X1 U549 ( .A1(n780), .A2(n776), .ZN(n593) );
  NAND2_X1 U550 ( .A1(n712), .A2(n613), .ZN(n421) );
  NOR2_X2 U551 ( .A1(n425), .A2(n512), .ZN(n513) );
  NOR2_X2 U552 ( .A1(n585), .A2(n580), .ZN(n594) );
  XOR2_X2 U553 ( .A(KEYINPUT4), .B(KEYINPUT65), .Z(n491) );
  XNOR2_X2 U554 ( .A(n484), .B(G472), .ZN(n586) );
  NAND2_X1 U555 ( .A1(n432), .A2(n430), .ZN(n588) );
  NAND2_X1 U556 ( .A1(n738), .A2(n353), .ZN(n434) );
  AND2_X1 U557 ( .A1(n437), .A2(n620), .ZN(n435) );
  INV_X1 U558 ( .A(n695), .ZN(n436) );
  XNOR2_X1 U559 ( .A(n593), .B(KEYINPUT46), .ZN(n437) );
  XNOR2_X1 U560 ( .A(n439), .B(n587), .ZN(n590) );
  NAND2_X1 U561 ( .A1(n586), .A2(n603), .ZN(n439) );
  XNOR2_X2 U562 ( .A(n445), .B(n560), .ZN(n686) );
  INV_X1 U563 ( .A(KEYINPUT47), .ZN(n444) );
  XNOR2_X2 U564 ( .A(n447), .B(G125), .ZN(n493) );
  INV_X1 U565 ( .A(KEYINPUT44), .ZN(n448) );
  INV_X1 U566 ( .A(n639), .ZN(n640) );
  XNOR2_X1 U567 ( .A(KEYINPUT33), .B(KEYINPUT70), .ZN(n486) );
  XNOR2_X1 U568 ( .A(n471), .B(n490), .ZN(n472) );
  XNOR2_X1 U569 ( .A(n475), .B(n472), .ZN(n738) );
  BUF_X1 U570 ( .A(n757), .Z(n759) );
  BUF_X1 U571 ( .A(n655), .Z(n658) );
  NAND2_X1 U572 ( .A1(n629), .A2(G234), .ZN(n450) );
  XOR2_X1 U573 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n452) );
  XNOR2_X1 U574 ( .A(G128), .B(G137), .ZN(n451) );
  XNOR2_X1 U575 ( .A(n452), .B(n451), .ZN(n454) );
  INV_X1 U576 ( .A(G119), .ZN(n453) );
  XOR2_X2 U577 ( .A(KEYINPUT64), .B(G953), .Z(n768) );
  NAND2_X1 U578 ( .A1(n768), .A2(G234), .ZN(n457) );
  XNOR2_X1 U579 ( .A(n457), .B(n456), .ZN(n537) );
  NAND2_X1 U580 ( .A1(n537), .A2(G221), .ZN(n458) );
  XNOR2_X1 U581 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U582 ( .A(n515), .B(n460), .ZN(n639) );
  NAND2_X1 U583 ( .A1(G217), .A2(n461), .ZN(n463) );
  INV_X1 U584 ( .A(KEYINPUT25), .ZN(n462) );
  XNOR2_X2 U585 ( .A(G128), .B(G143), .ZN(n492) );
  XNOR2_X1 U586 ( .A(G134), .B(n492), .ZN(n530) );
  INV_X1 U587 ( .A(n530), .ZN(n467) );
  XNOR2_X2 U588 ( .A(n467), .B(n466), .ZN(n765) );
  XNOR2_X2 U589 ( .A(n765), .B(G146), .ZN(n475) );
  XNOR2_X1 U590 ( .A(G101), .B(n468), .ZN(n470) );
  NAND2_X1 U591 ( .A1(G227), .A2(n768), .ZN(n469) );
  XNOR2_X1 U592 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U593 ( .A(n758), .B(KEYINPUT69), .ZN(n490) );
  INV_X1 U594 ( .A(n475), .ZN(n474) );
  NAND2_X1 U595 ( .A1(n474), .A2(n473), .ZN(n477) );
  NAND2_X1 U596 ( .A1(n475), .A2(G131), .ZN(n476) );
  NAND2_X1 U597 ( .A1(n477), .A2(n476), .ZN(n483) );
  XNOR2_X2 U598 ( .A(G101), .B(KEYINPUT3), .ZN(n478) );
  XNOR2_X1 U599 ( .A(n479), .B(KEYINPUT72), .ZN(n522) );
  NAND2_X1 U600 ( .A1(G210), .A2(n522), .ZN(n480) );
  XNOR2_X1 U601 ( .A(n365), .B(n480), .ZN(n481) );
  NAND2_X1 U602 ( .A1(n664), .A2(n527), .ZN(n484) );
  XNOR2_X1 U603 ( .A(n586), .B(KEYINPUT6), .ZN(n602) );
  NOR2_X2 U604 ( .A1(n485), .A2(n602), .ZN(n487) );
  XNOR2_X2 U605 ( .A(n489), .B(n488), .ZN(n757) );
  XNOR2_X1 U606 ( .A(n757), .B(n490), .ZN(n501) );
  XOR2_X1 U607 ( .A(KEYINPUT17), .B(n491), .Z(n495) );
  XOR2_X1 U608 ( .A(n492), .B(n493), .Z(n494) );
  XNOR2_X1 U609 ( .A(n495), .B(n494), .ZN(n499) );
  NAND2_X1 U610 ( .A1(G224), .A2(n768), .ZN(n497) );
  XNOR2_X1 U611 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U612 ( .A(n499), .B(n498), .ZN(n500) );
  NAND2_X1 U613 ( .A1(n527), .A2(n502), .ZN(n504) );
  NAND2_X1 U614 ( .A1(n504), .A2(G210), .ZN(n503) );
  NAND2_X1 U615 ( .A1(n504), .A2(G214), .ZN(n714) );
  XOR2_X1 U616 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n507) );
  NAND2_X1 U617 ( .A1(G237), .A2(G234), .ZN(n506) );
  XNOR2_X1 U618 ( .A(n507), .B(n506), .ZN(n510) );
  NAND2_X1 U619 ( .A1(n510), .A2(G952), .ZN(n508) );
  XNOR2_X1 U620 ( .A(n508), .B(KEYINPUT88), .ZN(n728) );
  NOR2_X1 U621 ( .A1(n728), .A2(G953), .ZN(n574) );
  XNOR2_X1 U622 ( .A(KEYINPUT89), .B(G898), .ZN(n753) );
  NAND2_X1 U623 ( .A1(n753), .A2(G953), .ZN(n509) );
  XNOR2_X1 U624 ( .A(n509), .B(KEYINPUT90), .ZN(n760) );
  NAND2_X1 U625 ( .A1(G902), .A2(n510), .ZN(n571) );
  NOR2_X1 U626 ( .A1(n760), .A2(n571), .ZN(n511) );
  NOR2_X1 U627 ( .A1(n574), .A2(n511), .ZN(n512) );
  XNOR2_X2 U628 ( .A(n513), .B(KEYINPUT0), .ZN(n556) );
  INV_X1 U629 ( .A(n556), .ZN(n514) );
  XOR2_X1 U630 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n517) );
  XNOR2_X1 U631 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U632 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U633 ( .A(n521), .B(KEYINPUT95), .Z(n524) );
  AND2_X1 U634 ( .A1(n522), .A2(G214), .ZN(n523) );
  NAND2_X1 U635 ( .A1(n649), .A2(n527), .ZN(n529) );
  XOR2_X1 U636 ( .A(KEYINPUT13), .B(G475), .Z(n528) );
  XNOR2_X1 U637 ( .A(n532), .B(n531), .ZN(n536) );
  XNOR2_X1 U638 ( .A(n530), .B(n538), .ZN(n746) );
  AND2_X1 U639 ( .A1(n559), .A2(n541), .ZN(n596) );
  NAND2_X1 U640 ( .A1(n539), .A2(n596), .ZN(n540) );
  NOR2_X1 U641 ( .A1(n717), .A2(n584), .ZN(n542) );
  NAND2_X1 U642 ( .A1(n556), .A2(n542), .ZN(n544) );
  INV_X1 U643 ( .A(KEYINPUT22), .ZN(n543) );
  INV_X1 U644 ( .A(n701), .ZN(n562) );
  INV_X1 U645 ( .A(n586), .ZN(n549) );
  INV_X1 U646 ( .A(n549), .ZN(n705) );
  AND2_X1 U647 ( .A1(n602), .A2(n623), .ZN(n546) );
  NOR2_X1 U648 ( .A1(n548), .A2(n549), .ZN(n550) );
  XNOR2_X1 U649 ( .A(n550), .B(KEYINPUT92), .ZN(n709) );
  AND2_X1 U650 ( .A1(n556), .A2(n709), .ZN(n552) );
  INV_X1 U651 ( .A(KEYINPUT31), .ZN(n551) );
  AND2_X1 U652 ( .A1(n553), .A2(n588), .ZN(n578) );
  INV_X1 U653 ( .A(n578), .ZN(n554) );
  NOR2_X1 U654 ( .A1(n705), .A2(n554), .ZN(n555) );
  AND2_X1 U655 ( .A1(n361), .A2(n555), .ZN(n676) );
  OR2_X1 U656 ( .A1(n559), .A2(n558), .ZN(n557) );
  INV_X1 U657 ( .A(n557), .ZN(n690) );
  INV_X1 U658 ( .A(KEYINPUT98), .ZN(n560) );
  INV_X1 U659 ( .A(n360), .ZN(n561) );
  NOR2_X1 U660 ( .A1(n623), .A2(n562), .ZN(n563) );
  AND2_X1 U661 ( .A1(n602), .A2(n563), .ZN(n564) );
  NAND2_X1 U662 ( .A1(n567), .A2(n566), .ZN(n569) );
  INV_X1 U663 ( .A(KEYINPUT45), .ZN(n568) );
  NOR2_X2 U664 ( .A1(n632), .A2(n629), .ZN(n570) );
  XNOR2_X1 U665 ( .A(n570), .B(KEYINPUT78), .ZN(n628) );
  XOR2_X1 U666 ( .A(KEYINPUT80), .B(KEYINPUT39), .Z(n583) );
  OR2_X1 U667 ( .A1(n571), .A2(n403), .ZN(n572) );
  NOR2_X1 U668 ( .A1(G900), .A2(n572), .ZN(n573) );
  NOR2_X1 U669 ( .A1(n574), .A2(n573), .ZN(n585) );
  NAND2_X1 U670 ( .A1(n714), .A2(n586), .ZN(n577) );
  XNOR2_X1 U671 ( .A(KEYINPUT104), .B(KEYINPUT30), .ZN(n575) );
  XNOR2_X1 U672 ( .A(n575), .B(KEYINPUT103), .ZN(n576) );
  XNOR2_X1 U673 ( .A(n577), .B(n576), .ZN(n579) );
  NAND2_X1 U674 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U675 ( .A1(n594), .A2(n715), .ZN(n582) );
  XNOR2_X1 U676 ( .A(n583), .B(n582), .ZN(n591) );
  NOR2_X1 U677 ( .A1(n591), .A2(n557), .ZN(n695) );
  XOR2_X1 U678 ( .A(KEYINPUT105), .B(KEYINPUT28), .Z(n587) );
  INV_X1 U679 ( .A(n588), .ZN(n589) );
  INV_X1 U680 ( .A(n729), .ZN(n712) );
  NOR2_X1 U681 ( .A1(n591), .A2(n442), .ZN(n592) );
  XNOR2_X1 U682 ( .A(n592), .B(KEYINPUT40), .ZN(n780) );
  INV_X1 U683 ( .A(n594), .ZN(n598) );
  INV_X1 U684 ( .A(n581), .ZN(n595) );
  NAND2_X1 U685 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U686 ( .A1(n598), .A2(n597), .ZN(n682) );
  XOR2_X1 U687 ( .A(KEYINPUT76), .B(n599), .Z(n600) );
  NOR2_X1 U688 ( .A1(n682), .A2(n600), .ZN(n601) );
  XNOR2_X1 U689 ( .A(n601), .B(KEYINPUT74), .ZN(n612) );
  INV_X1 U690 ( .A(n602), .ZN(n604) );
  NAND2_X1 U691 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U692 ( .A(KEYINPUT107), .B(n621), .ZN(n609) );
  BUF_X1 U693 ( .A(n606), .Z(n607) );
  INV_X1 U694 ( .A(n607), .ZN(n608) );
  NOR2_X1 U695 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U696 ( .A(n610), .B(KEYINPUT36), .ZN(n611) );
  NAND2_X1 U697 ( .A1(n611), .A2(n623), .ZN(n693) );
  NAND2_X1 U698 ( .A1(n612), .A2(n693), .ZN(n619) );
  XNOR2_X1 U699 ( .A(n614), .B(KEYINPUT75), .ZN(n617) );
  NOR2_X1 U700 ( .A1(KEYINPUT47), .A2(n360), .ZN(n615) );
  NAND2_X1 U701 ( .A1(n683), .A2(n615), .ZN(n616) );
  NAND2_X1 U702 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U703 ( .A1(n621), .A2(n714), .ZN(n622) );
  XNOR2_X1 U704 ( .A(n622), .B(KEYINPUT101), .ZN(n624) );
  INV_X1 U705 ( .A(n623), .ZN(n697) );
  NAND2_X1 U706 ( .A1(n624), .A2(n697), .ZN(n625) );
  XNOR2_X1 U707 ( .A(KEYINPUT43), .B(n625), .ZN(n626) );
  XNOR2_X1 U708 ( .A(n767), .B(KEYINPUT71), .ZN(n627) );
  INV_X1 U709 ( .A(n629), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n630), .A2(KEYINPUT2), .ZN(n631) );
  INV_X1 U711 ( .A(n750), .ZN(n634) );
  INV_X1 U712 ( .A(n767), .ZN(n633) );
  INV_X1 U713 ( .A(KEYINPUT66), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n364), .A2(G217), .ZN(n641) );
  XNOR2_X1 U715 ( .A(n641), .B(n640), .ZN(n644) );
  NOR2_X1 U716 ( .A1(n403), .A2(G952), .ZN(n643) );
  INV_X1 U717 ( .A(KEYINPUT84), .ZN(n642) );
  NAND2_X1 U718 ( .A1(n644), .A2(n745), .ZN(n645) );
  XNOR2_X1 U719 ( .A(n645), .B(KEYINPUT123), .ZN(G66) );
  XOR2_X1 U720 ( .A(G101), .B(n646), .Z(G3) );
  XOR2_X1 U721 ( .A(G110), .B(n647), .Z(G12) );
  NAND2_X1 U722 ( .A1(n363), .A2(G475), .ZN(n651) );
  XOR2_X1 U723 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n648) );
  XNOR2_X1 U724 ( .A(n651), .B(n650), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n652), .A2(n745), .ZN(n654) );
  INV_X1 U726 ( .A(KEYINPUT60), .ZN(n653) );
  XNOR2_X1 U727 ( .A(n654), .B(n653), .ZN(G60) );
  NAND2_X1 U728 ( .A1(n364), .A2(G210), .ZN(n660) );
  XNOR2_X1 U729 ( .A(KEYINPUT82), .B(KEYINPUT54), .ZN(n656) );
  XOR2_X1 U730 ( .A(n656), .B(KEYINPUT55), .Z(n657) );
  XNOR2_X1 U731 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U732 ( .A1(n661), .A2(n745), .ZN(n663) );
  INV_X1 U733 ( .A(KEYINPUT56), .ZN(n662) );
  XNOR2_X1 U734 ( .A(n663), .B(n662), .ZN(G51) );
  NAND2_X1 U735 ( .A1(n364), .A2(G472), .ZN(n669) );
  BUF_X1 U736 ( .A(n664), .Z(n665) );
  XNOR2_X1 U737 ( .A(n665), .B(KEYINPUT108), .ZN(n667) );
  XOR2_X1 U738 ( .A(KEYINPUT62), .B(KEYINPUT83), .Z(n666) );
  XNOR2_X1 U739 ( .A(n669), .B(n668), .ZN(n670) );
  NAND2_X1 U740 ( .A1(n670), .A2(n745), .ZN(n671) );
  XNOR2_X1 U741 ( .A(n671), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U742 ( .A1(n686), .A2(n676), .ZN(n672) );
  XNOR2_X1 U743 ( .A(n672), .B(G104), .ZN(G6) );
  XOR2_X1 U744 ( .A(KEYINPUT27), .B(KEYINPUT110), .Z(n674) );
  XNOR2_X1 U745 ( .A(G107), .B(KEYINPUT26), .ZN(n673) );
  XNOR2_X1 U746 ( .A(n674), .B(n673), .ZN(n675) );
  XOR2_X1 U747 ( .A(KEYINPUT109), .B(n675), .Z(n678) );
  NAND2_X1 U748 ( .A1(n676), .A2(n690), .ZN(n677) );
  XNOR2_X1 U749 ( .A(n678), .B(n677), .ZN(G9) );
  XOR2_X1 U750 ( .A(KEYINPUT29), .B(KEYINPUT111), .Z(n680) );
  NAND2_X1 U751 ( .A1(n683), .A2(n690), .ZN(n679) );
  XNOR2_X1 U752 ( .A(n680), .B(n679), .ZN(n681) );
  XOR2_X1 U753 ( .A(G128), .B(n681), .Z(G30) );
  XOR2_X1 U754 ( .A(G143), .B(n682), .Z(G45) );
  NAND2_X1 U755 ( .A1(n683), .A2(n686), .ZN(n684) );
  XNOR2_X1 U756 ( .A(n684), .B(KEYINPUT112), .ZN(n685) );
  XNOR2_X1 U757 ( .A(G146), .B(n685), .ZN(G48) );
  XOR2_X1 U758 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n688) );
  NAND2_X1 U759 ( .A1(n691), .A2(n686), .ZN(n687) );
  XNOR2_X1 U760 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U761 ( .A(G113), .B(n689), .ZN(G15) );
  NAND2_X1 U762 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U763 ( .A(n692), .B(G116), .ZN(G18) );
  XOR2_X1 U764 ( .A(G125), .B(KEYINPUT37), .Z(n694) );
  XNOR2_X1 U765 ( .A(n693), .B(n694), .ZN(G27) );
  XOR2_X1 U766 ( .A(G134), .B(n695), .Z(G36) );
  XNOR2_X1 U767 ( .A(n696), .B(KEYINPUT2), .ZN(n734) );
  XOR2_X1 U768 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n700) );
  NAND2_X1 U769 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U770 ( .A(n700), .B(n699), .ZN(n708) );
  NOR2_X1 U771 ( .A1(n702), .A2(n423), .ZN(n703) );
  XOR2_X1 U772 ( .A(KEYINPUT49), .B(n703), .Z(n704) );
  NOR2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U774 ( .A(n706), .B(KEYINPUT115), .ZN(n707) );
  NOR2_X1 U775 ( .A1(n708), .A2(n707), .ZN(n710) );
  NOR2_X1 U776 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U777 ( .A(KEYINPUT51), .B(n711), .ZN(n713) );
  NAND2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n725) );
  NOR2_X1 U779 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U780 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U781 ( .A(KEYINPUT117), .B(n718), .Z(n721) );
  NOR2_X1 U782 ( .A1(n719), .A2(n360), .ZN(n720) );
  NOR2_X1 U783 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U784 ( .A1(n730), .A2(n722), .ZN(n723) );
  XOR2_X1 U785 ( .A(KEYINPUT118), .B(n723), .Z(n724) );
  NAND2_X1 U786 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U787 ( .A(KEYINPUT52), .B(n726), .Z(n727) );
  NOR2_X1 U788 ( .A1(n728), .A2(n727), .ZN(n732) );
  NOR2_X1 U789 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U790 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U791 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U792 ( .A1(G953), .A2(n735), .ZN(n736) );
  XOR2_X1 U793 ( .A(KEYINPUT53), .B(n736), .Z(n737) );
  XNOR2_X1 U794 ( .A(KEYINPUT119), .B(n737), .ZN(G75) );
  NAND2_X1 U795 ( .A1(n363), .A2(G469), .ZN(n742) );
  XOR2_X1 U796 ( .A(n738), .B(KEYINPUT120), .Z(n740) );
  XOR2_X1 U797 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n739) );
  XNOR2_X1 U798 ( .A(n742), .B(n741), .ZN(n743) );
  NAND2_X1 U799 ( .A1(n743), .A2(n745), .ZN(n744) );
  XNOR2_X1 U800 ( .A(n744), .B(KEYINPUT121), .ZN(G54) );
  INV_X1 U801 ( .A(n745), .ZN(n749) );
  NAND2_X1 U802 ( .A1(n348), .A2(G478), .ZN(n747) );
  XNOR2_X1 U803 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X1 U804 ( .A1(n749), .A2(n748), .ZN(G63) );
  NOR2_X1 U805 ( .A1(n750), .A2(G953), .ZN(n756) );
  NAND2_X1 U806 ( .A1(G953), .A2(G224), .ZN(n751) );
  XOR2_X1 U807 ( .A(KEYINPUT61), .B(n751), .Z(n752) );
  NOR2_X1 U808 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U809 ( .A(n754), .B(KEYINPUT124), .ZN(n755) );
  NOR2_X1 U810 ( .A1(n756), .A2(n755), .ZN(n764) );
  XNOR2_X1 U811 ( .A(n759), .B(n758), .ZN(n761) );
  NAND2_X1 U812 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U813 ( .A(n762), .B(KEYINPUT125), .ZN(n763) );
  XOR2_X1 U814 ( .A(n764), .B(n763), .Z(G69) );
  XNOR2_X1 U815 ( .A(n766), .B(n765), .ZN(n770) );
  XNOR2_X1 U816 ( .A(n767), .B(n770), .ZN(n769) );
  NAND2_X1 U817 ( .A1(n769), .A2(n403), .ZN(n774) );
  XNOR2_X1 U818 ( .A(G227), .B(n770), .ZN(n771) );
  NAND2_X1 U819 ( .A1(n771), .A2(G900), .ZN(n772) );
  NAND2_X1 U820 ( .A1(n772), .A2(G953), .ZN(n773) );
  NAND2_X1 U821 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U822 ( .A(KEYINPUT126), .B(n775), .ZN(G72) );
  XNOR2_X1 U823 ( .A(G137), .B(n776), .ZN(n777) );
  XNOR2_X1 U824 ( .A(n777), .B(KEYINPUT127), .ZN(G39) );
  XNOR2_X1 U825 ( .A(G140), .B(n778), .ZN(G42) );
  XNOR2_X1 U826 ( .A(n362), .B(G119), .ZN(G21) );
  XOR2_X1 U827 ( .A(G131), .B(n780), .Z(G33) );
endmodule

