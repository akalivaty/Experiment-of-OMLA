

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U554 ( .A(n689), .B(n688), .ZN(n787) );
  XNOR2_X1 U555 ( .A(G299), .B(G290), .ZN(n688) );
  NOR2_X1 U556 ( .A1(G299), .A2(n820), .ZN(n816) );
  XNOR2_X1 U557 ( .A(G166), .B(n685), .ZN(n686) );
  OR2_X1 U558 ( .A1(n891), .A2(n890), .ZN(n908) );
  XNOR2_X1 U559 ( .A(n711), .B(KEYINPUT115), .ZN(n712) );
  OR2_X1 U560 ( .A1(G301), .A2(n834), .ZN(n520) );
  XOR2_X1 U561 ( .A(KEYINPUT28), .B(n821), .Z(n521) );
  XNOR2_X1 U562 ( .A(KEYINPUT91), .B(n888), .ZN(n522) );
  INV_X1 U563 ( .A(n850), .ZN(n824) );
  AND2_X1 U564 ( .A1(n827), .A2(n520), .ZN(n840) );
  NOR2_X1 U565 ( .A1(n840), .A2(n839), .ZN(n841) );
  NAND2_X1 U566 ( .A1(n883), .A2(n799), .ZN(n850) );
  XNOR2_X1 U567 ( .A(G305), .B(n686), .ZN(n687) );
  NAND2_X1 U568 ( .A1(G160), .A2(G40), .ZN(n882) );
  NAND2_X1 U569 ( .A1(n522), .A2(n889), .ZN(n890) );
  XOR2_X1 U570 ( .A(KEYINPUT17), .B(n538), .Z(n644) );
  INV_X1 U571 ( .A(KEYINPUT117), .ZN(n758) );
  XNOR2_X1 U572 ( .A(KEYINPUT67), .B(n523), .ZN(n700) );
  NOR2_X1 U573 ( .A1(G651), .A2(n673), .ZN(n701) );
  XNOR2_X1 U574 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U575 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U576 ( .A1(G651), .A2(G543), .ZN(n704) );
  NAND2_X1 U577 ( .A1(G91), .A2(n704), .ZN(n525) );
  XOR2_X1 U578 ( .A(KEYINPUT0), .B(G543), .Z(n673) );
  XOR2_X1 U579 ( .A(G651), .B(KEYINPUT66), .Z(n527) );
  OR2_X1 U580 ( .A1(n673), .A2(n527), .ZN(n523) );
  NAND2_X1 U581 ( .A1(G78), .A2(n700), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U583 ( .A(KEYINPUT70), .B(n526), .Z(n532) );
  NOR2_X1 U584 ( .A1(G543), .A2(n527), .ZN(n528) );
  XOR2_X1 U585 ( .A(KEYINPUT1), .B(n528), .Z(n705) );
  NAND2_X1 U586 ( .A1(G65), .A2(n705), .ZN(n530) );
  NAND2_X1 U587 ( .A1(G53), .A2(n701), .ZN(n529) );
  AND2_X1 U588 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n532), .A2(n531), .ZN(G299) );
  INV_X1 U590 ( .A(G2104), .ZN(n533) );
  NOR2_X1 U591 ( .A1(n533), .A2(G2105), .ZN(n534) );
  XNOR2_X2 U592 ( .A(n534), .B(KEYINPUT64), .ZN(n645) );
  NAND2_X1 U593 ( .A1(n645), .A2(G101), .ZN(n535) );
  XOR2_X1 U594 ( .A(KEYINPUT23), .B(n535), .Z(n537) );
  AND2_X1 U595 ( .A1(n533), .A2(G2105), .ZN(n640) );
  NAND2_X1 U596 ( .A1(n640), .A2(G125), .ZN(n536) );
  NAND2_X1 U597 ( .A1(n537), .A2(n536), .ZN(n542) );
  NOR2_X1 U598 ( .A1(G2104), .A2(G2105), .ZN(n538) );
  NAND2_X1 U599 ( .A1(G137), .A2(n644), .ZN(n540) );
  AND2_X1 U600 ( .A1(G2104), .A2(G2105), .ZN(n638) );
  NAND2_X1 U601 ( .A1(G113), .A2(n638), .ZN(n539) );
  NAND2_X1 U602 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U603 ( .A1(n542), .A2(n541), .ZN(G160) );
  NAND2_X1 U604 ( .A1(G86), .A2(n704), .ZN(n544) );
  NAND2_X1 U605 ( .A1(G61), .A2(n705), .ZN(n543) );
  NAND2_X1 U606 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U607 ( .A(KEYINPUT76), .B(n545), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G73), .A2(n700), .ZN(n546) );
  XOR2_X1 U609 ( .A(KEYINPUT2), .B(n546), .Z(n547) );
  XNOR2_X1 U610 ( .A(n547), .B(KEYINPUT77), .ZN(n549) );
  NAND2_X1 U611 ( .A1(G48), .A2(n701), .ZN(n548) );
  NAND2_X1 U612 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U613 ( .A(KEYINPUT78), .B(n552), .Z(G305) );
  NAND2_X1 U614 ( .A1(G88), .A2(n704), .ZN(n554) );
  NAND2_X1 U615 ( .A1(G75), .A2(n700), .ZN(n553) );
  NAND2_X1 U616 ( .A1(n554), .A2(n553), .ZN(n557) );
  NAND2_X1 U617 ( .A1(G62), .A2(n705), .ZN(n555) );
  XNOR2_X1 U618 ( .A(KEYINPUT79), .B(n555), .ZN(n556) );
  NOR2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n701), .A2(G50), .ZN(n558) );
  NAND2_X1 U621 ( .A1(n559), .A2(n558), .ZN(G303) );
  INV_X1 U622 ( .A(G303), .ZN(G166) );
  NAND2_X1 U623 ( .A1(G60), .A2(n705), .ZN(n561) );
  NAND2_X1 U624 ( .A1(G47), .A2(n701), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U626 ( .A1(G85), .A2(n704), .ZN(n562) );
  XNOR2_X1 U627 ( .A(KEYINPUT65), .B(n562), .ZN(n563) );
  NOR2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U629 ( .A1(n700), .A2(G72), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(G290) );
  NAND2_X1 U631 ( .A1(G138), .A2(n644), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G102), .A2(n645), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n572) );
  NAND2_X1 U634 ( .A1(G126), .A2(n640), .ZN(n570) );
  NAND2_X1 U635 ( .A1(G114), .A2(n638), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U637 ( .A1(n572), .A2(n571), .ZN(G164) );
  NAND2_X1 U638 ( .A1(G124), .A2(n640), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(KEYINPUT44), .ZN(n576) );
  NAND2_X1 U640 ( .A1(G136), .A2(n644), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n574), .B(KEYINPUT108), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n638), .A2(G112), .ZN(n578) );
  NAND2_X1 U644 ( .A1(G100), .A2(n645), .ZN(n577) );
  NAND2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U646 ( .A1(n580), .A2(n579), .ZN(G162) );
  XOR2_X1 U647 ( .A(KEYINPUT73), .B(KEYINPUT18), .Z(n582) );
  NAND2_X1 U648 ( .A1(G123), .A2(n640), .ZN(n581) );
  XNOR2_X1 U649 ( .A(n582), .B(n581), .ZN(n589) );
  NAND2_X1 U650 ( .A1(G135), .A2(n644), .ZN(n584) );
  NAND2_X1 U651 ( .A1(G111), .A2(n638), .ZN(n583) );
  NAND2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U653 ( .A1(n645), .A2(G99), .ZN(n585) );
  XOR2_X1 U654 ( .A(KEYINPUT74), .B(n585), .Z(n586) );
  NOR2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n943) );
  NAND2_X1 U657 ( .A1(G127), .A2(n640), .ZN(n591) );
  NAND2_X1 U658 ( .A1(G115), .A2(n638), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U660 ( .A(KEYINPUT47), .B(n592), .ZN(n598) );
  NAND2_X1 U661 ( .A1(G139), .A2(n644), .ZN(n593) );
  XOR2_X1 U662 ( .A(KEYINPUT112), .B(n593), .Z(n596) );
  NAND2_X1 U663 ( .A1(G103), .A2(n645), .ZN(n594) );
  XNOR2_X1 U664 ( .A(KEYINPUT111), .B(n594), .ZN(n595) );
  NOR2_X1 U665 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U666 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U667 ( .A(KEYINPUT113), .B(n599), .ZN(n938) );
  XNOR2_X1 U668 ( .A(n943), .B(n938), .ZN(n609) );
  NAND2_X1 U669 ( .A1(G129), .A2(n640), .ZN(n601) );
  NAND2_X1 U670 ( .A1(G117), .A2(n638), .ZN(n600) );
  NAND2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U672 ( .A1(G105), .A2(n645), .ZN(n602) );
  XOR2_X1 U673 ( .A(KEYINPUT38), .B(n602), .Z(n603) );
  NOR2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U675 ( .A(KEYINPUT89), .B(n605), .Z(n607) );
  NAND2_X1 U676 ( .A1(n644), .A2(G141), .ZN(n606) );
  NAND2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n892) );
  XOR2_X1 U678 ( .A(G160), .B(n892), .Z(n608) );
  XNOR2_X1 U679 ( .A(n609), .B(n608), .ZN(n625) );
  XOR2_X1 U680 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n611) );
  XNOR2_X1 U681 ( .A(KEYINPUT114), .B(KEYINPUT110), .ZN(n610) );
  XNOR2_X1 U682 ( .A(n611), .B(n610), .ZN(n621) );
  NAND2_X1 U683 ( .A1(G130), .A2(n640), .ZN(n613) );
  NAND2_X1 U684 ( .A1(G118), .A2(n638), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n613), .A2(n612), .ZN(n619) );
  NAND2_X1 U686 ( .A1(G142), .A2(n644), .ZN(n615) );
  NAND2_X1 U687 ( .A1(G106), .A2(n645), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U689 ( .A(KEYINPUT45), .B(n616), .ZN(n617) );
  XNOR2_X1 U690 ( .A(KEYINPUT109), .B(n617), .ZN(n618) );
  NOR2_X1 U691 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U692 ( .A(n621), .B(n620), .Z(n623) );
  XNOR2_X1 U693 ( .A(G164), .B(G162), .ZN(n622) );
  XNOR2_X1 U694 ( .A(n623), .B(n622), .ZN(n624) );
  XOR2_X1 U695 ( .A(n625), .B(n624), .Z(n652) );
  NAND2_X1 U696 ( .A1(G104), .A2(n645), .ZN(n626) );
  XNOR2_X1 U697 ( .A(n626), .B(KEYINPUT82), .ZN(n628) );
  NAND2_X1 U698 ( .A1(G140), .A2(n644), .ZN(n627) );
  NAND2_X1 U699 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U700 ( .A(KEYINPUT34), .B(n629), .ZN(n635) );
  NAND2_X1 U701 ( .A1(n638), .A2(G116), .ZN(n630) );
  XOR2_X1 U702 ( .A(KEYINPUT83), .B(n630), .Z(n632) );
  NAND2_X1 U703 ( .A1(n640), .A2(G128), .ZN(n631) );
  NAND2_X1 U704 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U705 ( .A(n633), .B(KEYINPUT35), .Z(n634) );
  NOR2_X1 U706 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U707 ( .A(KEYINPUT36), .B(n636), .Z(n637) );
  XOR2_X1 U708 ( .A(KEYINPUT84), .B(n637), .Z(n903) );
  NAND2_X1 U709 ( .A1(G107), .A2(n638), .ZN(n639) );
  XNOR2_X1 U710 ( .A(n639), .B(KEYINPUT86), .ZN(n643) );
  NAND2_X1 U711 ( .A1(G119), .A2(n640), .ZN(n641) );
  XOR2_X1 U712 ( .A(KEYINPUT85), .B(n641), .Z(n642) );
  NAND2_X1 U713 ( .A1(n643), .A2(n642), .ZN(n650) );
  NAND2_X1 U714 ( .A1(G131), .A2(n644), .ZN(n647) );
  NAND2_X1 U715 ( .A1(G95), .A2(n645), .ZN(n646) );
  NAND2_X1 U716 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U717 ( .A(KEYINPUT87), .B(n648), .Z(n649) );
  NOR2_X1 U718 ( .A1(n650), .A2(n649), .ZN(n893) );
  XNOR2_X1 U719 ( .A(n903), .B(n893), .ZN(n651) );
  XNOR2_X1 U720 ( .A(n652), .B(n651), .ZN(n653) );
  NOR2_X1 U721 ( .A1(G37), .A2(n653), .ZN(G395) );
  NAND2_X1 U722 ( .A1(n704), .A2(G89), .ZN(n654) );
  XNOR2_X1 U723 ( .A(n654), .B(KEYINPUT4), .ZN(n656) );
  NAND2_X1 U724 ( .A1(G76), .A2(n700), .ZN(n655) );
  NAND2_X1 U725 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U726 ( .A(n657), .B(KEYINPUT5), .ZN(n662) );
  NAND2_X1 U727 ( .A1(G63), .A2(n705), .ZN(n659) );
  NAND2_X1 U728 ( .A1(G51), .A2(n701), .ZN(n658) );
  NAND2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U730 ( .A(KEYINPUT6), .B(n660), .Z(n661) );
  NAND2_X1 U731 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n663), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U733 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U734 ( .A1(G64), .A2(n705), .ZN(n665) );
  NAND2_X1 U735 ( .A1(G52), .A2(n701), .ZN(n664) );
  NAND2_X1 U736 ( .A1(n665), .A2(n664), .ZN(n672) );
  NAND2_X1 U737 ( .A1(n700), .A2(G77), .ZN(n666) );
  XNOR2_X1 U738 ( .A(n666), .B(KEYINPUT68), .ZN(n668) );
  NAND2_X1 U739 ( .A1(G90), .A2(n704), .ZN(n667) );
  NAND2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U741 ( .A(KEYINPUT69), .B(n669), .ZN(n670) );
  XNOR2_X1 U742 ( .A(KEYINPUT9), .B(n670), .ZN(n671) );
  NOR2_X1 U743 ( .A1(n672), .A2(n671), .ZN(G171) );
  NAND2_X1 U744 ( .A1(G87), .A2(n673), .ZN(n675) );
  NAND2_X1 U745 ( .A1(G74), .A2(G651), .ZN(n674) );
  NAND2_X1 U746 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U747 ( .A1(n705), .A2(n676), .ZN(n678) );
  NAND2_X1 U748 ( .A1(n701), .A2(G49), .ZN(n677) );
  NAND2_X1 U749 ( .A1(n678), .A2(n677), .ZN(G288) );
  XNOR2_X1 U750 ( .A(G286), .B(G171), .ZN(n690) );
  NAND2_X1 U751 ( .A1(G93), .A2(n704), .ZN(n680) );
  NAND2_X1 U752 ( .A1(G67), .A2(n705), .ZN(n679) );
  NAND2_X1 U753 ( .A1(n680), .A2(n679), .ZN(n684) );
  NAND2_X1 U754 ( .A1(G80), .A2(n700), .ZN(n682) );
  NAND2_X1 U755 ( .A1(G55), .A2(n701), .ZN(n681) );
  NAND2_X1 U756 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U757 ( .A1(n684), .A2(n683), .ZN(n789) );
  XNOR2_X1 U758 ( .A(G288), .B(KEYINPUT19), .ZN(n685) );
  XOR2_X1 U759 ( .A(n789), .B(n687), .Z(n689) );
  XNOR2_X1 U760 ( .A(n690), .B(n787), .ZN(n713) );
  NAND2_X1 U761 ( .A1(G56), .A2(n705), .ZN(n691) );
  XOR2_X1 U762 ( .A(KEYINPUT14), .B(n691), .Z(n697) );
  NAND2_X1 U763 ( .A1(n704), .A2(G81), .ZN(n692) );
  XNOR2_X1 U764 ( .A(n692), .B(KEYINPUT12), .ZN(n694) );
  NAND2_X1 U765 ( .A1(G68), .A2(n700), .ZN(n693) );
  NAND2_X1 U766 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U767 ( .A(KEYINPUT13), .B(n695), .Z(n696) );
  NOR2_X1 U768 ( .A1(n697), .A2(n696), .ZN(n699) );
  NAND2_X1 U769 ( .A1(n701), .A2(G43), .ZN(n698) );
  NAND2_X1 U770 ( .A1(n699), .A2(n698), .ZN(n1002) );
  NAND2_X1 U771 ( .A1(G79), .A2(n700), .ZN(n703) );
  NAND2_X1 U772 ( .A1(G54), .A2(n701), .ZN(n702) );
  NAND2_X1 U773 ( .A1(n703), .A2(n702), .ZN(n709) );
  NAND2_X1 U774 ( .A1(G92), .A2(n704), .ZN(n707) );
  NAND2_X1 U775 ( .A1(G66), .A2(n705), .ZN(n706) );
  NAND2_X1 U776 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U777 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U778 ( .A(n710), .B(KEYINPUT15), .ZN(n990) );
  INV_X1 U779 ( .A(n990), .ZN(n782) );
  XNOR2_X1 U780 ( .A(n1002), .B(n782), .ZN(n711) );
  NOR2_X1 U781 ( .A1(G37), .A2(n714), .ZN(G397) );
  XOR2_X1 U782 ( .A(G2451), .B(KEYINPUT102), .Z(n716) );
  XNOR2_X1 U783 ( .A(G2443), .B(G2446), .ZN(n715) );
  XNOR2_X1 U784 ( .A(n716), .B(n715), .ZN(n720) );
  XOR2_X1 U785 ( .A(G2435), .B(G2438), .Z(n718) );
  XNOR2_X1 U786 ( .A(G2454), .B(G2430), .ZN(n717) );
  XNOR2_X1 U787 ( .A(n718), .B(n717), .ZN(n719) );
  XOR2_X1 U788 ( .A(n720), .B(n719), .Z(n722) );
  XNOR2_X1 U789 ( .A(G2427), .B(KEYINPUT100), .ZN(n721) );
  XNOR2_X1 U790 ( .A(n722), .B(n721), .ZN(n725) );
  XOR2_X1 U791 ( .A(G1341), .B(G1348), .Z(n723) );
  XNOR2_X1 U792 ( .A(KEYINPUT101), .B(n723), .ZN(n724) );
  XOR2_X1 U793 ( .A(n725), .B(n724), .Z(n726) );
  AND2_X1 U794 ( .A1(G14), .A2(n726), .ZN(G401) );
  XNOR2_X1 U795 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 U796 ( .A(G132), .ZN(G219) );
  XNOR2_X1 U797 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  INV_X1 U798 ( .A(G57), .ZN(G237) );
  INV_X1 U799 ( .A(G120), .ZN(G236) );
  INV_X1 U800 ( .A(G108), .ZN(G238) );
  NOR2_X1 U801 ( .A1(G219), .A2(G220), .ZN(n727) );
  XOR2_X1 U802 ( .A(KEYINPUT80), .B(n727), .Z(n728) );
  XNOR2_X1 U803 ( .A(n728), .B(KEYINPUT22), .ZN(n729) );
  NOR2_X1 U804 ( .A1(G218), .A2(n729), .ZN(n730) );
  NAND2_X1 U805 ( .A1(G96), .A2(n730), .ZN(n914) );
  NAND2_X1 U806 ( .A1(G2106), .A2(n914), .ZN(n731) );
  XNOR2_X1 U807 ( .A(n731), .B(KEYINPUT81), .ZN(n735) );
  INV_X1 U808 ( .A(G567), .ZN(n768) );
  NOR2_X1 U809 ( .A1(G236), .A2(G238), .ZN(n732) );
  NAND2_X1 U810 ( .A1(G69), .A2(n732), .ZN(n733) );
  NOR2_X1 U811 ( .A1(G237), .A2(n733), .ZN(n916) );
  NOR2_X1 U812 ( .A1(n768), .A2(n916), .ZN(n734) );
  NOR2_X1 U813 ( .A1(n735), .A2(n734), .ZN(G319) );
  XOR2_X1 U814 ( .A(KEYINPUT42), .B(G2072), .Z(n737) );
  XNOR2_X1 U815 ( .A(G2067), .B(G2078), .ZN(n736) );
  XNOR2_X1 U816 ( .A(n737), .B(n736), .ZN(n738) );
  XOR2_X1 U817 ( .A(n738), .B(G2100), .Z(n740) );
  XNOR2_X1 U818 ( .A(G2090), .B(G2084), .ZN(n739) );
  XNOR2_X1 U819 ( .A(n740), .B(n739), .ZN(n744) );
  XOR2_X1 U820 ( .A(G2096), .B(KEYINPUT43), .Z(n742) );
  XNOR2_X1 U821 ( .A(KEYINPUT103), .B(G2678), .ZN(n741) );
  XNOR2_X1 U822 ( .A(n742), .B(n741), .ZN(n743) );
  XOR2_X1 U823 ( .A(n744), .B(n743), .Z(G227) );
  XOR2_X1 U824 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n746) );
  XNOR2_X1 U825 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n745) );
  XNOR2_X1 U826 ( .A(n746), .B(n745), .ZN(n747) );
  XOR2_X1 U827 ( .A(n747), .B(G2474), .Z(n749) );
  XNOR2_X1 U828 ( .A(G1996), .B(G1991), .ZN(n748) );
  XNOR2_X1 U829 ( .A(n749), .B(n748), .ZN(n757) );
  XOR2_X1 U830 ( .A(G1976), .B(G1966), .Z(n751) );
  XNOR2_X1 U831 ( .A(G1986), .B(G1971), .ZN(n750) );
  XNOR2_X1 U832 ( .A(n751), .B(n750), .ZN(n755) );
  XOR2_X1 U833 ( .A(KEYINPUT106), .B(G1981), .Z(n753) );
  XNOR2_X1 U834 ( .A(G1961), .B(G1956), .ZN(n752) );
  XNOR2_X1 U835 ( .A(n753), .B(n752), .ZN(n754) );
  XOR2_X1 U836 ( .A(n755), .B(n754), .Z(n756) );
  XNOR2_X1 U837 ( .A(n757), .B(n756), .ZN(G229) );
  NOR2_X1 U838 ( .A1(G395), .A2(G397), .ZN(n759) );
  XNOR2_X1 U839 ( .A(n759), .B(n758), .ZN(n765) );
  NOR2_X1 U840 ( .A1(G227), .A2(G229), .ZN(n760) );
  XOR2_X1 U841 ( .A(KEYINPUT49), .B(n760), .Z(n761) );
  NAND2_X1 U842 ( .A1(G319), .A2(n761), .ZN(n762) );
  NOR2_X1 U843 ( .A1(G401), .A2(n762), .ZN(n763) );
  XNOR2_X1 U844 ( .A(KEYINPUT116), .B(n763), .ZN(n764) );
  NAND2_X1 U845 ( .A1(n765), .A2(n764), .ZN(G225) );
  AND2_X1 U846 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U847 ( .A1(G7), .A2(G661), .ZN(n766) );
  XNOR2_X1 U848 ( .A(n766), .B(KEYINPUT10), .ZN(n767) );
  XNOR2_X1 U849 ( .A(KEYINPUT72), .B(n767), .ZN(G223) );
  NOR2_X1 U850 ( .A1(G223), .A2(n768), .ZN(n769) );
  XNOR2_X1 U851 ( .A(n769), .B(KEYINPUT11), .ZN(G234) );
  INV_X1 U852 ( .A(G860), .ZN(n784) );
  OR2_X1 U853 ( .A1(n1002), .A2(n784), .ZN(G153) );
  INV_X1 U854 ( .A(G171), .ZN(G301) );
  NAND2_X1 U855 ( .A1(G868), .A2(G301), .ZN(n771) );
  INV_X1 U856 ( .A(G868), .ZN(n790) );
  NAND2_X1 U857 ( .A1(n990), .A2(n790), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(G284) );
  NOR2_X1 U859 ( .A1(G868), .A2(G299), .ZN(n773) );
  NOR2_X1 U860 ( .A1(G286), .A2(n790), .ZN(n772) );
  NOR2_X1 U861 ( .A1(n773), .A2(n772), .ZN(G297) );
  NAND2_X1 U862 ( .A1(n784), .A2(G559), .ZN(n774) );
  NAND2_X1 U863 ( .A1(n774), .A2(n782), .ZN(n775) );
  XNOR2_X1 U864 ( .A(n775), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U865 ( .A1(G868), .A2(n1002), .ZN(n778) );
  NAND2_X1 U866 ( .A1(G868), .A2(n782), .ZN(n776) );
  NOR2_X1 U867 ( .A1(G559), .A2(n776), .ZN(n777) );
  NOR2_X1 U868 ( .A1(n778), .A2(n777), .ZN(G282) );
  XNOR2_X1 U869 ( .A(n943), .B(G2096), .ZN(n779) );
  XNOR2_X1 U870 ( .A(n779), .B(KEYINPUT75), .ZN(n781) );
  INV_X1 U871 ( .A(G2100), .ZN(n780) );
  NAND2_X1 U872 ( .A1(n781), .A2(n780), .ZN(G156) );
  NAND2_X1 U873 ( .A1(G559), .A2(n782), .ZN(n783) );
  XOR2_X1 U874 ( .A(n1002), .B(n783), .Z(n786) );
  NAND2_X1 U875 ( .A1(n784), .A2(n786), .ZN(n785) );
  XOR2_X1 U876 ( .A(n785), .B(n789), .Z(G145) );
  XOR2_X1 U877 ( .A(n787), .B(n786), .Z(n788) );
  NOR2_X1 U878 ( .A1(n790), .A2(n788), .ZN(n792) );
  AND2_X1 U879 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U880 ( .A1(n792), .A2(n791), .ZN(G295) );
  NAND2_X1 U881 ( .A1(G2078), .A2(G2084), .ZN(n793) );
  XOR2_X1 U882 ( .A(KEYINPUT20), .B(n793), .Z(n794) );
  NAND2_X1 U883 ( .A1(G2090), .A2(n794), .ZN(n795) );
  XNOR2_X1 U884 ( .A(KEYINPUT21), .B(n795), .ZN(n796) );
  NAND2_X1 U885 ( .A1(n796), .A2(G2072), .ZN(G158) );
  INV_X1 U886 ( .A(G319), .ZN(n798) );
  NAND2_X1 U887 ( .A1(G483), .A2(G661), .ZN(n797) );
  NOR2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n913) );
  NAND2_X1 U889 ( .A1(n913), .A2(G36), .ZN(G176) );
  NOR2_X1 U890 ( .A1(G164), .A2(G1384), .ZN(n883) );
  INV_X1 U891 ( .A(n882), .ZN(n799) );
  NAND2_X1 U892 ( .A1(G8), .A2(n850), .ZN(n876) );
  NOR2_X1 U893 ( .A1(G1981), .A2(G305), .ZN(n800) );
  XOR2_X1 U894 ( .A(n800), .B(KEYINPUT24), .Z(n801) );
  NOR2_X1 U895 ( .A1(n876), .A2(n801), .ZN(n881) );
  NAND2_X1 U896 ( .A1(G1348), .A2(n850), .ZN(n803) );
  NAND2_X1 U897 ( .A1(G2067), .A2(n824), .ZN(n802) );
  NAND2_X1 U898 ( .A1(n803), .A2(n802), .ZN(n810) );
  NOR2_X1 U899 ( .A1(n990), .A2(n810), .ZN(n809) );
  INV_X1 U900 ( .A(G1996), .ZN(n920) );
  NOR2_X1 U901 ( .A1(n850), .A2(n920), .ZN(n804) );
  XOR2_X1 U902 ( .A(n804), .B(KEYINPUT26), .Z(n806) );
  NAND2_X1 U903 ( .A1(n850), .A2(G1341), .ZN(n805) );
  NAND2_X1 U904 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U905 ( .A1(n807), .A2(n1002), .ZN(n808) );
  NOR2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n812) );
  AND2_X1 U907 ( .A1(n990), .A2(n810), .ZN(n811) );
  NOR2_X1 U908 ( .A1(n812), .A2(n811), .ZN(n819) );
  INV_X1 U909 ( .A(KEYINPUT93), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n824), .A2(G2072), .ZN(n813) );
  XOR2_X1 U911 ( .A(n813), .B(KEYINPUT27), .Z(n815) );
  NAND2_X1 U912 ( .A1(G1956), .A2(n850), .ZN(n814) );
  NAND2_X1 U913 ( .A1(n815), .A2(n814), .ZN(n820) );
  XNOR2_X1 U914 ( .A(n817), .B(n816), .ZN(n818) );
  NOR2_X1 U915 ( .A1(n819), .A2(n818), .ZN(n822) );
  NAND2_X1 U916 ( .A1(G299), .A2(n820), .ZN(n821) );
  NOR2_X1 U917 ( .A1(n822), .A2(n521), .ZN(n823) );
  XNOR2_X1 U918 ( .A(n823), .B(KEYINPUT29), .ZN(n827) );
  NAND2_X1 U919 ( .A1(G1961), .A2(n850), .ZN(n826) );
  XOR2_X1 U920 ( .A(KEYINPUT25), .B(G2078), .Z(n922) );
  NAND2_X1 U921 ( .A1(n824), .A2(n922), .ZN(n825) );
  NAND2_X1 U922 ( .A1(n826), .A2(n825), .ZN(n834) );
  NOR2_X1 U923 ( .A1(G2084), .A2(n850), .ZN(n843) );
  INV_X1 U924 ( .A(G8), .ZN(n828) );
  NOR2_X1 U925 ( .A1(n828), .A2(G1966), .ZN(n829) );
  AND2_X1 U926 ( .A1(n850), .A2(n829), .ZN(n830) );
  XOR2_X1 U927 ( .A(n830), .B(KEYINPUT92), .Z(n842) );
  NAND2_X1 U928 ( .A1(G8), .A2(n842), .ZN(n831) );
  NOR2_X1 U929 ( .A1(n843), .A2(n831), .ZN(n832) );
  XOR2_X1 U930 ( .A(n832), .B(KEYINPUT30), .Z(n833) );
  NOR2_X1 U931 ( .A1(G168), .A2(n833), .ZN(n837) );
  NAND2_X1 U932 ( .A1(G301), .A2(n834), .ZN(n835) );
  XOR2_X1 U933 ( .A(KEYINPUT94), .B(n835), .Z(n836) );
  NOR2_X1 U934 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n838), .B(KEYINPUT31), .ZN(n839) );
  XNOR2_X1 U936 ( .A(KEYINPUT95), .B(n841), .ZN(n848) );
  AND2_X1 U937 ( .A1(n848), .A2(n842), .ZN(n845) );
  NAND2_X1 U938 ( .A1(G8), .A2(n843), .ZN(n844) );
  NAND2_X1 U939 ( .A1(n845), .A2(n844), .ZN(n846) );
  XNOR2_X1 U940 ( .A(KEYINPUT96), .B(n846), .ZN(n859) );
  AND2_X1 U941 ( .A1(G286), .A2(G8), .ZN(n847) );
  NAND2_X1 U942 ( .A1(n848), .A2(n847), .ZN(n856) );
  NOR2_X1 U943 ( .A1(G1971), .A2(n876), .ZN(n849) );
  XNOR2_X1 U944 ( .A(KEYINPUT97), .B(n849), .ZN(n853) );
  NOR2_X1 U945 ( .A1(G2090), .A2(n850), .ZN(n851) );
  NOR2_X1 U946 ( .A1(G166), .A2(n851), .ZN(n852) );
  NAND2_X1 U947 ( .A1(n853), .A2(n852), .ZN(n854) );
  OR2_X1 U948 ( .A1(n828), .A2(n854), .ZN(n855) );
  AND2_X1 U949 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U950 ( .A(KEYINPUT32), .B(n857), .ZN(n858) );
  NAND2_X1 U951 ( .A1(n859), .A2(n858), .ZN(n875) );
  NOR2_X1 U952 ( .A1(G1976), .A2(G288), .ZN(n865) );
  NOR2_X1 U953 ( .A1(G1971), .A2(G303), .ZN(n860) );
  NOR2_X1 U954 ( .A1(n865), .A2(n860), .ZN(n997) );
  INV_X1 U955 ( .A(KEYINPUT33), .ZN(n861) );
  AND2_X1 U956 ( .A1(n997), .A2(n861), .ZN(n862) );
  NAND2_X1 U957 ( .A1(n875), .A2(n862), .ZN(n871) );
  INV_X1 U958 ( .A(n876), .ZN(n863) );
  NAND2_X1 U959 ( .A1(G1976), .A2(G288), .ZN(n993) );
  AND2_X1 U960 ( .A1(n863), .A2(n993), .ZN(n864) );
  NOR2_X1 U961 ( .A1(KEYINPUT33), .A2(n864), .ZN(n869) );
  NAND2_X1 U962 ( .A1(n865), .A2(KEYINPUT33), .ZN(n866) );
  OR2_X1 U963 ( .A1(n866), .A2(n876), .ZN(n867) );
  XOR2_X1 U964 ( .A(G1981), .B(G305), .Z(n1005) );
  NAND2_X1 U965 ( .A1(n867), .A2(n1005), .ZN(n868) );
  NOR2_X1 U966 ( .A1(n869), .A2(n868), .ZN(n870) );
  NAND2_X1 U967 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U968 ( .A(n872), .B(KEYINPUT98), .ZN(n879) );
  NOR2_X1 U969 ( .A1(G2090), .A2(G303), .ZN(n873) );
  NAND2_X1 U970 ( .A1(G8), .A2(n873), .ZN(n874) );
  NAND2_X1 U971 ( .A1(n875), .A2(n874), .ZN(n877) );
  NAND2_X1 U972 ( .A1(n877), .A2(n876), .ZN(n878) );
  NAND2_X1 U973 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U974 ( .A1(n881), .A2(n880), .ZN(n891) );
  NOR2_X1 U975 ( .A1(n883), .A2(n882), .ZN(n905) );
  XNOR2_X1 U976 ( .A(G2067), .B(KEYINPUT37), .ZN(n902) );
  NOR2_X1 U977 ( .A1(n903), .A2(n902), .ZN(n950) );
  NAND2_X1 U978 ( .A1(n905), .A2(n950), .ZN(n900) );
  XOR2_X1 U979 ( .A(KEYINPUT88), .B(G1991), .Z(n928) );
  NOR2_X1 U980 ( .A1(n928), .A2(n893), .ZN(n885) );
  AND2_X1 U981 ( .A1(n892), .A2(G1996), .ZN(n884) );
  NOR2_X1 U982 ( .A1(n885), .A2(n884), .ZN(n948) );
  XOR2_X1 U983 ( .A(n905), .B(KEYINPUT90), .Z(n886) );
  NOR2_X1 U984 ( .A1(n948), .A2(n886), .ZN(n897) );
  INV_X1 U985 ( .A(n897), .ZN(n887) );
  NAND2_X1 U986 ( .A1(n900), .A2(n887), .ZN(n888) );
  XNOR2_X1 U987 ( .A(G1986), .B(G290), .ZN(n999) );
  NAND2_X1 U988 ( .A1(n999), .A2(n905), .ZN(n889) );
  NOR2_X1 U989 ( .A1(G1996), .A2(n892), .ZN(n955) );
  AND2_X1 U990 ( .A1(n928), .A2(n893), .ZN(n946) );
  NOR2_X1 U991 ( .A1(G1986), .A2(G290), .ZN(n894) );
  XOR2_X1 U992 ( .A(n894), .B(KEYINPUT99), .Z(n895) );
  NOR2_X1 U993 ( .A1(n946), .A2(n895), .ZN(n896) );
  NOR2_X1 U994 ( .A1(n897), .A2(n896), .ZN(n898) );
  NOR2_X1 U995 ( .A1(n955), .A2(n898), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n899), .B(KEYINPUT39), .ZN(n901) );
  NAND2_X1 U997 ( .A1(n901), .A2(n900), .ZN(n904) );
  NAND2_X1 U998 ( .A1(n903), .A2(n902), .ZN(n952) );
  NAND2_X1 U999 ( .A1(n904), .A2(n952), .ZN(n906) );
  NAND2_X1 U1000 ( .A1(n906), .A2(n905), .ZN(n907) );
  NAND2_X1 U1001 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1002 ( .A(n909), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U1003 ( .A(G223), .ZN(n910) );
  NAND2_X1 U1004 ( .A1(G2106), .A2(n910), .ZN(G217) );
  AND2_X1 U1005 ( .A1(G15), .A2(G2), .ZN(n911) );
  NAND2_X1 U1006 ( .A1(G661), .A2(n911), .ZN(G259) );
  NAND2_X1 U1007 ( .A1(G3), .A2(G1), .ZN(n912) );
  NAND2_X1 U1008 ( .A1(n913), .A2(n912), .ZN(G188) );
  INV_X1 U1010 ( .A(n914), .ZN(n915) );
  NAND2_X1 U1011 ( .A1(n916), .A2(n915), .ZN(G261) );
  INV_X1 U1012 ( .A(G261), .ZN(G325) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G69), .ZN(G235) );
  INV_X1 U1015 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U1016 ( .A(G2084), .B(KEYINPUT54), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(n917), .B(G34), .ZN(n936) );
  XNOR2_X1 U1018 ( .A(G2090), .B(G35), .ZN(n933) );
  XNOR2_X1 U1019 ( .A(G2067), .B(G26), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(G33), .B(G2072), .ZN(n918) );
  NOR2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n927) );
  XNOR2_X1 U1022 ( .A(G32), .B(n920), .ZN(n921) );
  NAND2_X1 U1023 ( .A1(n921), .A2(G28), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(G27), .B(n922), .ZN(n923) );
  XNOR2_X1 U1025 ( .A(KEYINPUT122), .B(n923), .ZN(n924) );
  NOR2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n930) );
  XOR2_X1 U1028 ( .A(G25), .B(n928), .Z(n929) );
  NOR2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(KEYINPUT53), .B(n931), .ZN(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(n934), .B(KEYINPUT123), .ZN(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n1021) );
  NAND2_X1 U1034 ( .A1(KEYINPUT55), .A2(n1021), .ZN(n937) );
  NAND2_X1 U1035 ( .A1(G11), .A2(n937), .ZN(n1020) );
  XNOR2_X1 U1036 ( .A(G2072), .B(n938), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(n939), .B(KEYINPUT121), .ZN(n941) );
  XOR2_X1 U1038 ( .A(G2078), .B(G164), .Z(n940) );
  NOR2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1040 ( .A(KEYINPUT50), .B(n942), .Z(n962) );
  XNOR2_X1 U1041 ( .A(G160), .B(G2084), .ZN(n944) );
  NAND2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(n951), .B(KEYINPUT118), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n959) );
  XOR2_X1 U1048 ( .A(G2090), .B(G162), .Z(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1050 ( .A(KEYINPUT51), .B(n956), .Z(n957) );
  XNOR2_X1 U1051 ( .A(n957), .B(KEYINPUT119), .ZN(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1053 ( .A(KEYINPUT120), .B(n960), .Z(n961) );
  NOR2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(KEYINPUT52), .B(n963), .ZN(n965) );
  INV_X1 U1056 ( .A(KEYINPUT55), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1058 ( .A1(n966), .A2(G29), .ZN(n1018) );
  XOR2_X1 U1059 ( .A(G1986), .B(G24), .Z(n970) );
  XNOR2_X1 U1060 ( .A(G1971), .B(G22), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(G23), .B(G1976), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(n972), .B(n971), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(G1961), .B(G5), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(G21), .B(G1966), .ZN(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n986) );
  XOR2_X1 U1070 ( .A(G1348), .B(KEYINPUT59), .Z(n977) );
  XNOR2_X1 U1071 ( .A(G4), .B(n977), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(G20), .B(G1956), .ZN(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(G1341), .B(G19), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(G1981), .B(G6), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(KEYINPUT60), .B(n984), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1080 ( .A(n987), .B(KEYINPUT126), .Z(n988) );
  XNOR2_X1 U1081 ( .A(KEYINPUT61), .B(n988), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(G16), .A2(n989), .ZN(n1015) );
  XOR2_X1 U1083 ( .A(G16), .B(KEYINPUT56), .Z(n1013) );
  XNOR2_X1 U1084 ( .A(G171), .B(G1961), .ZN(n1001) );
  XNOR2_X1 U1085 ( .A(G1348), .B(KEYINPUT124), .ZN(n991) );
  XNOR2_X1 U1086 ( .A(n991), .B(n990), .ZN(n995) );
  NAND2_X1 U1087 ( .A1(G1971), .A2(G303), .ZN(n992) );
  NAND2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1011) );
  XNOR2_X1 U1093 ( .A(n1002), .B(G1341), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(G299), .B(G1956), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(G168), .B(G1966), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1098 ( .A(n1007), .B(KEYINPUT57), .ZN(n1008) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(KEYINPUT127), .B(n1016), .Z(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1025) );
  INV_X1 U1106 ( .A(n1021), .ZN(n1023) );
  NOR2_X1 U1107 ( .A1(G29), .A2(KEYINPUT55), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

