//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT32), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(G143), .B(G146), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT0), .B(G128), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT64), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT0), .A2(G128), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT0), .A2(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n197), .A2(G146), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n206), .B1(new_n195), .B2(G143), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n197), .A2(KEYINPUT65), .A3(G146), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n205), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n194), .A2(new_n204), .B1(new_n209), .B2(new_n200), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  INV_X1    g025(.A(G134), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(G137), .ZN(new_n213));
  INV_X1    g027(.A(G137), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT11), .A3(G134), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(G137), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G131), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n213), .A2(new_n215), .A3(new_n219), .A4(new_n216), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n210), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT1), .B1(new_n197), .B2(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G128), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n209), .A2(new_n225), .B1(new_n227), .B2(new_n199), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n212), .A2(G137), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n214), .A2(G134), .ZN(new_n230));
  OAI21_X1  g044(.A(G131), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n220), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n223), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n207), .A2(new_n208), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n196), .A3(new_n225), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n227), .A2(new_n199), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n220), .A2(new_n231), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n238), .A3(KEYINPUT66), .ZN(new_n239));
  INV_X1    g053(.A(G119), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G116), .ZN(new_n241));
  INV_X1    g055(.A(G116), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G119), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT2), .B(G113), .ZN(new_n245));
  XOR2_X1   g059(.A(new_n244), .B(new_n245), .Z(new_n246));
  NAND4_X1  g060(.A1(new_n222), .A2(new_n233), .A3(new_n239), .A4(new_n246), .ZN(new_n247));
  XOR2_X1   g061(.A(KEYINPUT67), .B(G237), .Z(new_n248));
  INV_X1    g062(.A(G953), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(G210), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT27), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT67), .B(G237), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G953), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT27), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(G210), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT26), .B(G101), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n251), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n256), .B1(new_n251), .B2(new_n255), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n247), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n237), .A2(new_n238), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n209), .A2(new_n200), .ZN(new_n262));
  NOR3_X1   g076(.A1(new_n192), .A2(new_n193), .A3(KEYINPUT64), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n203), .B1(new_n199), .B2(new_n202), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n218), .A2(new_n220), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n261), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n222), .A2(new_n233), .A3(new_n239), .A4(KEYINPUT30), .ZN(new_n270));
  INV_X1    g084(.A(new_n246), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n260), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT31), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT31), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n260), .A2(new_n272), .A3(new_n275), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n210), .A2(new_n221), .B1(new_n237), .B2(new_n238), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT28), .B1(new_n277), .B2(new_n246), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT68), .B1(new_n277), .B2(new_n246), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT68), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n267), .A2(new_n280), .A3(new_n271), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n281), .A3(new_n247), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n278), .B1(new_n282), .B2(KEYINPUT28), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n274), .B(new_n276), .C1(new_n283), .C2(new_n259), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n282), .A2(KEYINPUT28), .ZN(new_n287));
  INV_X1    g101(.A(new_n278), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n259), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n260), .A2(new_n272), .A3(new_n275), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n275), .B1(new_n260), .B2(new_n272), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT69), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n191), .B1(new_n286), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n272), .A2(new_n247), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT29), .B1(new_n297), .B2(new_n290), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n298), .B1(new_n289), .B2(new_n290), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n259), .A2(KEYINPUT29), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n222), .A2(new_n233), .A3(new_n239), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n271), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n247), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT70), .B1(new_n304), .B2(KEYINPUT28), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT28), .ZN(new_n307));
  AOI211_X1 g121(.A(new_n306), .B(new_n307), .C1(new_n303), .C2(new_n247), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n288), .B(new_n301), .C1(new_n305), .C2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n299), .A2(new_n300), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G472), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n296), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n284), .A2(new_n285), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n291), .A2(KEYINPUT69), .A3(new_n294), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT32), .B1(new_n315), .B2(new_n188), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n187), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n188), .B1(new_n286), .B2(new_n295), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n190), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n315), .A2(new_n191), .B1(G472), .B2(new_n310), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(KEYINPUT71), .ZN(new_n321));
  XNOR2_X1  g135(.A(G125), .B(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n195), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n325));
  INV_X1    g139(.A(G125), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(KEYINPUT74), .A2(G125), .A3(G140), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(KEYINPUT16), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT16), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n330), .B1(new_n326), .B2(G140), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n195), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n240), .A2(G128), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n224), .A2(G119), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n336), .B(KEYINPUT73), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT24), .B(G110), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n224), .A2(KEYINPUT23), .A3(G119), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n240), .A2(G128), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n334), .B(new_n341), .C1(new_n342), .C2(KEYINPUT23), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(G110), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n323), .B(new_n333), .C1(new_n340), .C2(new_n344), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n337), .A2(new_n339), .B1(G110), .B2(new_n343), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n329), .A2(new_n195), .A3(new_n331), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n346), .B1(new_n348), .B2(new_n332), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT22), .B(G137), .ZN(new_n351));
  INV_X1    g165(.A(G221), .ZN(new_n352));
  INV_X1    g166(.A(G234), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n352), .A2(new_n353), .A3(G953), .ZN(new_n354));
  XOR2_X1   g168(.A(new_n351), .B(new_n354), .Z(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n345), .A2(new_n349), .A3(new_n355), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT75), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT25), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(G902), .B1(new_n360), .B2(new_n361), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n359), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G217), .B1(new_n353), .B2(G902), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n366), .B(KEYINPUT72), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n357), .A2(new_n358), .A3(new_n364), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n362), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n365), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n367), .A2(G902), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n359), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n375));
  INV_X1    g189(.A(G107), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n375), .B1(new_n376), .B2(G104), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(G104), .ZN(new_n378));
  INV_X1    g192(.A(G104), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(KEYINPUT77), .A3(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G101), .ZN(new_n382));
  INV_X1    g196(.A(G101), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(G107), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n376), .A2(KEYINPUT3), .A3(G104), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT3), .B1(new_n376), .B2(G104), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n383), .B(new_n384), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n228), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT78), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n382), .A2(new_n387), .ZN(new_n391));
  INV_X1    g205(.A(new_n227), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n235), .B1(new_n209), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT78), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n388), .A2(new_n228), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n390), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n221), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT12), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT10), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n228), .A2(new_n400), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n394), .A2(new_n400), .B1(new_n401), .B2(new_n391), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT3), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n404), .B1(new_n379), .B2(G107), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n376), .A2(KEYINPUT3), .A3(G104), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n405), .A2(new_n406), .B1(new_n379), .B2(G107), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n403), .B1(new_n407), .B2(new_n383), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G101), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n407), .A2(new_n383), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT76), .B1(new_n412), .B2(new_n403), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT76), .ZN(new_n414));
  NOR4_X1   g228(.A1(new_n407), .A2(new_n414), .A3(KEYINPUT4), .A4(new_n383), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n411), .B(new_n210), .C1(new_n413), .C2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n402), .A2(new_n266), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G110), .B(G140), .ZN(new_n418));
  INV_X1    g232(.A(G227), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n419), .A2(G953), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n418), .B(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT12), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n397), .A2(new_n423), .A3(new_n221), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n399), .A2(new_n417), .A3(new_n422), .A4(new_n424), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n402), .A2(new_n266), .A3(new_n416), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n266), .B1(new_n402), .B2(new_n416), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n421), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G469), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n430), .A3(new_n300), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n399), .A2(new_n417), .A3(new_n424), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n421), .ZN(new_n433));
  OR3_X1    g247(.A1(new_n426), .A2(new_n427), .A3(new_n421), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(G469), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n430), .A2(new_n300), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n431), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT9), .B(G234), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n352), .B1(new_n440), .B2(new_n300), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AND4_X1   g258(.A1(new_n317), .A2(new_n321), .A3(new_n374), .A4(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G214), .B1(G237), .B2(G902), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G210), .B1(G237), .B2(G902), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n414), .B1(new_n410), .B2(KEYINPUT4), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n412), .A2(KEYINPUT76), .A3(new_n403), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n450), .A2(new_n451), .B1(new_n410), .B2(new_n408), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT80), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n241), .A2(new_n243), .A3(KEYINPUT5), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT5), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n240), .A3(G116), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G113), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT79), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n241), .A2(new_n243), .A3(KEYINPUT5), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT79), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n459), .A2(new_n460), .A3(G113), .A4(new_n456), .ZN(new_n461));
  OR2_X1    g275(.A1(new_n244), .A2(new_n245), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n458), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n453), .B1(new_n463), .B2(new_n388), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n244), .A2(new_n245), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n459), .A2(G113), .A3(new_n456), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n465), .B1(new_n466), .B2(KEYINPUT79), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n391), .A2(new_n467), .A3(KEYINPUT80), .A4(new_n461), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n452), .A2(new_n271), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(G110), .B(G122), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n469), .A2(KEYINPUT6), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n228), .A2(new_n326), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n472), .B1(new_n210), .B2(new_n326), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n249), .A2(G224), .ZN(new_n474));
  XOR2_X1   g288(.A(new_n473), .B(new_n474), .Z(new_n475));
  INV_X1    g289(.A(KEYINPUT81), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n469), .B2(new_n470), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n478), .B1(new_n469), .B2(new_n470), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n464), .A2(new_n468), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n271), .B(new_n411), .C1(new_n413), .C2(new_n415), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n470), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(KEYINPUT81), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n477), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT82), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n477), .A2(new_n479), .A3(KEYINPUT82), .A4(new_n484), .ZN(new_n488));
  AOI211_X1 g302(.A(new_n471), .B(new_n475), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT7), .ZN(new_n490));
  OR3_X1    g304(.A1(new_n473), .A2(new_n490), .A3(new_n474), .ZN(new_n491));
  INV_X1    g305(.A(new_n466), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n391), .B1(new_n492), .B2(new_n465), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n470), .B(KEYINPUT8), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n493), .B(new_n494), .C1(new_n391), .C2(new_n463), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n473), .B1(new_n490), .B2(new_n474), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n491), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n480), .A2(new_n470), .A3(new_n481), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n300), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n449), .B1(new_n489), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n471), .ZN(new_n502));
  INV_X1    g316(.A(new_n475), .ZN(new_n503));
  AOI211_X1 g317(.A(new_n476), .B(new_n470), .C1(new_n480), .C2(new_n481), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n498), .A2(KEYINPUT6), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT82), .B1(new_n506), .B2(new_n477), .ZN(new_n507));
  AND4_X1   g321(.A1(KEYINPUT82), .A2(new_n477), .A3(new_n479), .A4(new_n484), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n502), .B(new_n503), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n500), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(new_n448), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n447), .B1(new_n501), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n248), .A2(G214), .A3(new_n249), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(new_n197), .ZN(new_n514));
  AOI21_X1  g328(.A(G143), .B1(new_n253), .B2(G214), .ZN(new_n515));
  OAI211_X1 g329(.A(KEYINPUT18), .B(G131), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n327), .A2(G146), .A3(new_n328), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n323), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(new_n197), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n253), .A2(G143), .A3(G214), .ZN(new_n520));
  NAND2_X1  g334(.A1(KEYINPUT18), .A2(G131), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n516), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(G113), .B(G122), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT83), .B(G104), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n524), .B(new_n525), .Z(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(G131), .B1(new_n514), .B2(new_n515), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT17), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n519), .A2(new_n219), .A3(new_n520), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(KEYINPUT17), .B(G131), .C1(new_n514), .C2(new_n515), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT84), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n534), .B1(new_n348), .B2(new_n332), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n333), .A2(KEYINPUT84), .A3(new_n347), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n523), .B(new_n527), .C1(new_n532), .C2(new_n537), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n516), .A2(new_n518), .A3(new_n522), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT19), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n322), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n327), .A2(KEYINPUT19), .A3(new_n328), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n333), .B1(G146), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n528), .B2(new_n530), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n526), .B1(new_n539), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n538), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(G475), .A2(G902), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT20), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT20), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n547), .A2(new_n551), .A3(new_n548), .ZN(new_n552));
  INV_X1    g366(.A(new_n538), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n531), .A2(new_n535), .A3(new_n536), .A4(new_n533), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n527), .B1(new_n554), .B2(new_n523), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n300), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n550), .A2(new_n552), .B1(G475), .B2(new_n556), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n249), .A2(G952), .ZN(new_n558));
  NAND2_X1  g372(.A1(G234), .A2(G237), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n560), .B(KEYINPUT87), .Z(new_n561));
  AND3_X1   g375(.A1(new_n559), .A2(G902), .A3(G953), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT21), .B(G898), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G478), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n197), .A2(G128), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n224), .A2(G143), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT85), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n570), .B1(new_n568), .B2(new_n569), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n212), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(G116), .B(G122), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(new_n376), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT13), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n577), .B(G134), .C1(KEYINPUT13), .C2(new_n568), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n574), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n568), .A2(new_n569), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT85), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(G134), .A3(new_n571), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n574), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G122), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G116), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n376), .B1(new_n586), .B2(KEYINPUT14), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(new_n575), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n584), .A2(KEYINPUT86), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT86), .B1(new_n584), .B2(new_n588), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n580), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n440), .A2(G217), .A3(new_n249), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n572), .A2(new_n573), .A3(new_n212), .ZN(new_n594));
  AOI21_X1  g408(.A(G134), .B1(new_n582), .B2(new_n571), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n588), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT86), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n584), .A2(KEYINPUT86), .A3(new_n588), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n592), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n580), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n593), .A2(new_n602), .ZN(new_n603));
  AOI211_X1 g417(.A(KEYINPUT15), .B(new_n567), .C1(new_n603), .C2(new_n300), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n567), .A2(KEYINPUT15), .ZN(new_n605));
  AOI211_X1 g419(.A(G902), .B(new_n605), .C1(new_n593), .C2(new_n602), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n557), .A2(new_n566), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT88), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT88), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n557), .A2(new_n610), .A3(new_n566), .A4(new_n607), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n512), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n445), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  NAND2_X1  g430(.A1(new_n550), .A2(new_n552), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n556), .A2(G475), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT89), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(KEYINPUT89), .A2(KEYINPUT33), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n601), .B1(new_n600), .B2(new_n580), .ZN(new_n624));
  AOI211_X1 g438(.A(new_n579), .B(new_n592), .C1(new_n598), .C2(new_n599), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n593), .A2(new_n602), .A3(new_n620), .A4(new_n621), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT90), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n567), .A2(G902), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(G478), .B1(new_n603), .B2(new_n300), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n630), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n626), .B2(new_n627), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n629), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n634), .A2(KEYINPUT91), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT91), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n636), .A2(new_n629), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n632), .B1(new_n636), .B2(new_n629), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n566), .B(new_n619), .C1(new_n638), .C2(new_n642), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n509), .A2(new_n510), .A3(new_n448), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n448), .B1(new_n509), .B2(new_n510), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n446), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(G902), .B1(new_n313), .B2(new_n314), .ZN(new_n648));
  INV_X1    g462(.A(G472), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n318), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n650), .A2(new_n373), .A3(new_n443), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT34), .B(G104), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  OR2_X1    g468(.A1(new_n604), .A2(new_n606), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n557), .A3(new_n566), .ZN(new_n656));
  AOI211_X1 g470(.A(new_n447), .B(new_n656), .C1(new_n501), .C2(new_n511), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n651), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G107), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  NOR2_X1   g474(.A1(new_n350), .A2(KEYINPUT92), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n350), .A2(KEYINPUT92), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  OAI22_X1  g477(.A1(new_n661), .A2(new_n663), .B1(KEYINPUT36), .B2(new_n356), .ZN(new_n664));
  INV_X1    g478(.A(new_n661), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n356), .A2(KEYINPUT36), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n666), .A3(new_n662), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n664), .A2(new_n371), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n370), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT93), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT93), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n370), .A2(new_n671), .A3(new_n668), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n650), .A2(new_n443), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n512), .A3(new_n612), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT94), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n675), .B(new_n677), .ZN(G12));
  NOR2_X1   g492(.A1(new_n673), .A2(new_n443), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n317), .A2(new_n321), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n619), .A2(new_n607), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(G900), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n562), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n561), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n512), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n680), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(new_n224), .ZN(G30));
  NOR2_X1   g503(.A1(new_n644), .A2(new_n645), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT38), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT95), .B(KEYINPUT39), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n685), .B(new_n692), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n444), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT40), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n300), .B1(new_n304), .B2(new_n259), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n290), .B1(new_n272), .B2(new_n247), .ZN(new_n698));
  OAI21_X1  g512(.A(G472), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n319), .A2(new_n296), .A3(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n557), .A2(new_n607), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n702), .A2(new_n447), .A3(new_n669), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n696), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n694), .A2(new_n695), .ZN(new_n705));
  OR3_X1    g519(.A1(new_n691), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G143), .ZN(G45));
  AND3_X1   g521(.A1(new_n317), .A2(new_n321), .A3(new_n679), .ZN(new_n708));
  OAI21_X1  g522(.A(KEYINPUT91), .B1(new_n634), .B2(new_n637), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n640), .A2(new_n641), .A3(new_n639), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n685), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n619), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n646), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  NOR3_X1   g530(.A1(new_n312), .A2(new_n316), .A3(new_n187), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT71), .B1(new_n319), .B2(new_n320), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n429), .A2(new_n300), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(G469), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n442), .A3(new_n431), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT96), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n430), .B1(new_n429), .B2(new_n300), .ZN(new_n724));
  AOI211_X1 g538(.A(G469), .B(G902), .C1(new_n425), .C2(new_n428), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT96), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n442), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n723), .A2(new_n728), .A3(KEYINPUT97), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT97), .B1(new_n723), .B2(new_n728), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n719), .A2(new_n647), .A3(new_n731), .A4(new_n374), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT41), .B(G113), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G15));
  NAND4_X1  g548(.A1(new_n719), .A2(new_n731), .A3(new_n374), .A4(new_n657), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G116), .ZN(G18));
  INV_X1    g550(.A(KEYINPUT98), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n723), .A2(new_n728), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n737), .B1(new_n646), .B2(new_n738), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n723), .A2(new_n728), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n512), .A2(new_n740), .A3(KEYINPUT98), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n673), .ZN(new_n743));
  AND4_X1   g557(.A1(new_n612), .A2(new_n317), .A3(new_n321), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT99), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT99), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n742), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G119), .ZN(G21));
  OAI211_X1 g564(.A(new_n446), .B(new_n701), .C1(new_n644), .C2(new_n645), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n288), .B1(new_n305), .B2(new_n308), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n290), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n294), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n188), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n756), .B(new_n374), .C1(new_n648), .C2(new_n649), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n731), .A2(new_n752), .A3(new_n566), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G122), .ZN(G24));
  OAI211_X1 g574(.A(new_n756), .B(new_n669), .C1(new_n648), .C2(new_n649), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n557), .B1(new_n709), .B2(new_n710), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n763), .A3(new_n712), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n739), .B2(new_n741), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n326), .ZN(G27));
  INV_X1    g580(.A(new_n713), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n433), .A2(new_n434), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT100), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT100), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n433), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(G469), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n725), .A2(new_n436), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n441), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AND4_X1   g588(.A1(new_n446), .A2(new_n774), .A3(new_n501), .A4(new_n511), .ZN(new_n775));
  AOI211_X1 g589(.A(KEYINPUT101), .B(new_n373), .C1(new_n319), .C2(new_n320), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT101), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n189), .B1(new_n313), .B2(new_n314), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n296), .B(new_n311), .C1(new_n778), .C2(KEYINPUT32), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n777), .B1(new_n779), .B2(new_n374), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n767), .B(new_n775), .C1(new_n776), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT42), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n317), .A2(new_n321), .A3(new_n374), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n713), .A2(KEYINPUT42), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n775), .A3(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n782), .A2(KEYINPUT102), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT102), .B1(new_n782), .B2(new_n786), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G131), .ZN(G33));
  NAND3_X1  g604(.A1(new_n690), .A2(new_n446), .A3(new_n774), .ZN(new_n791));
  INV_X1    g605(.A(new_n686), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n783), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n212), .ZN(G36));
  NAND3_X1  g608(.A1(new_n769), .A2(KEYINPUT45), .A3(new_n771), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n430), .B1(new_n768), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT103), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n795), .A2(KEYINPUT103), .A3(new_n797), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n436), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(KEYINPUT46), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n431), .B1(new_n802), .B2(KEYINPUT46), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n441), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n806), .A2(new_n693), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n711), .A2(new_n557), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n808), .A2(KEYINPUT43), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(KEYINPUT43), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n650), .A3(new_n669), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT44), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n690), .A2(new_n446), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n811), .B2(new_n812), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n807), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G137), .ZN(G39));
  OAI22_X1  g631(.A1(new_n805), .A2(new_n441), .B1(KEYINPUT104), .B2(KEYINPUT47), .ZN(new_n818));
  XOR2_X1   g632(.A(KEYINPUT104), .B(KEYINPUT47), .Z(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n442), .B(new_n820), .C1(new_n803), .C2(new_n804), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n719), .A2(new_n814), .A3(new_n374), .A4(new_n713), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n818), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  XOR2_X1   g637(.A(KEYINPUT105), .B(G140), .Z(new_n824));
  XNOR2_X1  g638(.A(new_n823), .B(new_n824), .ZN(G42));
  INV_X1    g639(.A(KEYINPUT49), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n446), .B(new_n442), .C1(new_n726), .C2(new_n826), .ZN(new_n827));
  AOI211_X1 g641(.A(new_n827), .B(new_n808), .C1(new_n826), .C2(new_n726), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n700), .A2(new_n373), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n691), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n561), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n809), .A2(new_n831), .A3(new_n810), .ZN(new_n832));
  INV_X1    g646(.A(new_n814), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n740), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n776), .A2(new_n780), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g652(.A(new_n838), .B(KEYINPUT48), .Z(new_n839));
  NAND4_X1  g653(.A1(new_n809), .A2(new_n831), .A3(new_n758), .A4(new_n810), .ZN(new_n840));
  INV_X1    g654(.A(new_n742), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n829), .A2(new_n831), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n834), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n763), .ZN(new_n844));
  OAI221_X1 g658(.A(new_n558), .B1(new_n840), .B2(new_n841), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n691), .A2(new_n447), .A3(new_n740), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT50), .ZN(new_n848));
  OR3_X1    g662(.A1(new_n847), .A2(new_n840), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n847), .B2(new_n840), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR4_X1   g665(.A1(new_n834), .A2(new_n842), .A3(new_n619), .A4(new_n711), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(new_n835), .B2(new_n762), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n818), .A2(new_n821), .B1(new_n441), .B2(new_n726), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n840), .A2(new_n814), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n851), .B(new_n853), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(KEYINPUT112), .A3(KEYINPUT51), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT51), .B1(new_n856), .B2(KEYINPUT112), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n846), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT113), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(KEYINPUT113), .B(new_n846), .C1(new_n858), .C2(new_n859), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n669), .A2(new_n685), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n296), .A2(new_n699), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n774), .B(new_n866), .C1(new_n867), .C2(new_n316), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n751), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n708), .B2(new_n714), .ZN(new_n870));
  INV_X1    g684(.A(new_n764), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n646), .A2(new_n737), .A3(new_n738), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT98), .B1(new_n512), .B2(new_n740), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n680), .A2(new_n687), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n870), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT52), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n765), .A2(new_n688), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n879), .A2(KEYINPUT52), .A3(new_n870), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n445), .A2(new_n614), .B1(new_n647), .B2(new_n651), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT108), .ZN(new_n883));
  INV_X1    g697(.A(new_n656), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n884), .B(new_n446), .C1(new_n644), .C2(new_n645), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n651), .B1(new_n885), .B2(KEYINPUT107), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT107), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n512), .B2(new_n884), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n883), .B(new_n675), .C1(new_n886), .C2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n882), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n657), .A2(new_n887), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n885), .A2(KEYINPUT107), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(new_n651), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n883), .B1(new_n893), .B2(new_n675), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n784), .A2(new_n686), .A3(new_n775), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n619), .A2(new_n655), .A3(new_n685), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n690), .A2(new_n446), .A3(new_n897), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n680), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT109), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n871), .A2(new_n775), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n896), .A2(new_n899), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  OAI22_X1  g716(.A1(new_n680), .A2(new_n898), .B1(new_n764), .B2(new_n791), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT109), .B1(new_n903), .B2(new_n793), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n789), .A2(new_n881), .A3(new_n895), .A4(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT106), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n742), .A2(new_n747), .A3(new_n744), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n747), .B1(new_n742), .B2(new_n744), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n732), .A2(new_n735), .A3(new_n759), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n911), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n749), .A2(KEYINPUT106), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n865), .B1(new_n906), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n911), .B1(new_n748), .B2(new_n746), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n782), .A2(KEYINPUT53), .A3(new_n786), .ZN(new_n919));
  AND4_X1   g733(.A1(new_n918), .A2(new_n895), .A3(new_n905), .A4(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT111), .B1(new_n920), .B2(new_n881), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n918), .A2(new_n895), .A3(new_n905), .A4(new_n919), .ZN(new_n922));
  INV_X1    g736(.A(new_n881), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT111), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n916), .B(new_n917), .C1(new_n921), .C2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT110), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n910), .A2(new_n907), .A3(new_n911), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT106), .B1(new_n749), .B2(new_n913), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n788), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n782), .A2(KEYINPUT102), .A3(new_n786), .ZN(new_n932));
  AND4_X1   g746(.A1(new_n931), .A2(new_n895), .A3(new_n932), .A4(new_n905), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n930), .A2(new_n933), .A3(new_n865), .A4(new_n881), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT53), .B1(new_n906), .B2(new_n915), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT54), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n926), .A2(new_n927), .A3(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT110), .A4(KEYINPUT54), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n864), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(G952), .A2(G953), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT114), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n830), .B1(new_n939), .B2(new_n941), .ZN(G75));
  NOR2_X1   g756(.A1(new_n249), .A2(G952), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n930), .A2(new_n933), .A3(new_n881), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n920), .A2(KEYINPUT111), .A3(new_n881), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n924), .B1(new_n922), .B2(new_n923), .ZN(new_n946));
  AOI22_X1  g760(.A1(new_n865), .A2(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT116), .B1(new_n947), .B2(new_n300), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n945), .A2(new_n946), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n916), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT116), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n950), .A2(new_n951), .A3(G902), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n948), .A2(new_n449), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n502), .B1(new_n507), .B2(new_n508), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n475), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n509), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT55), .ZN(new_n957));
  XOR2_X1   g771(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n958));
  NOR2_X1   g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n943), .B1(new_n953), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n300), .B1(new_n949), .B2(new_n916), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT115), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(new_n962), .A3(G210), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT56), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n962), .B1(new_n961), .B2(G210), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n957), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n960), .A2(new_n967), .ZN(G51));
  INV_X1    g782(.A(new_n926), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n917), .B1(new_n949), .B2(new_n916), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n436), .B(KEYINPUT118), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT57), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n429), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n948), .A2(new_n952), .A3(new_n800), .A4(new_n801), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n943), .B1(new_n974), .B2(new_n975), .ZN(G54));
  AND2_X1   g790(.A1(KEYINPUT58), .A2(G475), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n948), .A2(new_n952), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n538), .A3(new_n546), .ZN(new_n979));
  INV_X1    g793(.A(new_n943), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n948), .A2(new_n952), .A3(new_n547), .A4(new_n977), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(G60));
  XOR2_X1   g796(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n983));
  NOR2_X1   g797(.A1(new_n567), .A2(new_n300), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n937), .A2(new_n938), .A3(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n628), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n628), .A2(new_n985), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n969), .B2(new_n970), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(KEYINPUT120), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT120), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n991), .B(new_n988), .C1(new_n969), .C2(new_n970), .ZN(new_n992));
  AOI221_X4 g806(.A(new_n943), .B1(new_n986), .B2(new_n987), .C1(new_n990), .C2(new_n992), .ZN(G63));
  INV_X1    g807(.A(KEYINPUT61), .ZN(new_n994));
  NAND2_X1  g808(.A1(G217), .A2(G902), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT60), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n947), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n664), .A2(new_n667), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT121), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n980), .B1(new_n997), .B2(new_n359), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n994), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OR2_X1    g817(.A1(new_n997), .A2(new_n359), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n1004), .A2(KEYINPUT61), .A3(new_n980), .A4(new_n1000), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1003), .A2(new_n1005), .ZN(G66));
  INV_X1    g820(.A(new_n563), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n249), .B1(new_n1007), .B2(G224), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n930), .A2(new_n895), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1008), .B1(new_n1009), .B2(new_n249), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n954), .B1(G898), .B2(new_n249), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1010), .B(new_n1011), .Z(G69));
  NAND2_X1  g826(.A1(new_n269), .A2(new_n270), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(new_n543), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1014), .B(KEYINPUT122), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n879), .A2(new_n715), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n706), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT62), .Z(new_n1018));
  NAND2_X1  g832(.A1(new_n844), .A2(new_n682), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT123), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n1020), .A2(new_n784), .A3(new_n694), .A4(new_n833), .ZN(new_n1021));
  AOI21_X1  g835(.A(KEYINPUT124), .B1(new_n816), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n816), .A2(KEYINPUT124), .A3(new_n1021), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  OAI211_X1 g838(.A(new_n1018), .B(new_n823), .C1(new_n1022), .C2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1015), .B1(new_n1025), .B2(new_n249), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1014), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n807), .A2(new_n752), .A3(new_n837), .ZN(new_n1028));
  NAND4_X1  g842(.A1(new_n816), .A2(new_n1028), .A3(new_n896), .A4(new_n1016), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n789), .A2(new_n823), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n249), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n683), .A2(G953), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1032), .B(KEYINPUT126), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1027), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n1026), .A2(new_n1034), .A3(KEYINPUT125), .ZN(new_n1035));
  OAI21_X1  g849(.A(G953), .B1(new_n419), .B2(new_n683), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1035), .B(new_n1036), .ZN(G72));
  NAND2_X1  g851(.A1(G472), .A2(G902), .ZN(new_n1038));
  XOR2_X1   g852(.A(new_n1038), .B(KEYINPUT63), .Z(new_n1039));
  OAI21_X1  g853(.A(new_n1039), .B1(new_n1025), .B2(new_n1009), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1040), .A2(new_n698), .ZN(new_n1041));
  OR2_X1    g855(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1039), .B1(new_n1042), .B2(new_n1009), .ZN(new_n1043));
  NOR2_X1   g857(.A1(new_n297), .A2(new_n259), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n943), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(new_n1039), .ZN(new_n1047));
  NOR3_X1   g861(.A1(new_n1044), .A2(new_n698), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n934), .A2(new_n935), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g863(.A(KEYINPUT127), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OR2_X1    g865(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1046), .B1(new_n1051), .B2(new_n1052), .ZN(G57));
endmodule


