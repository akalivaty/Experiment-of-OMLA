//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1184, new_n1185, new_n1186, new_n1187, new_n1189,
    new_n1190, new_n1191, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1247, new_n1248;
  OR3_X1    g0000(.A1(KEYINPUT64), .A2(G58), .A3(G68), .ZN(new_n201));
  OAI21_X1  g0001(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(G50), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G77), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT65), .Z(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT66), .ZN(new_n216));
  INV_X1    g0016(.A(G13), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n216), .B1(new_n209), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g0018(.A1(KEYINPUT66), .A2(G1), .A3(G13), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n210), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n203), .A2(new_n204), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(KEYINPUT67), .B(G238), .Z(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G58), .A2(G232), .ZN(new_n230));
  NAND4_X1  g0030(.A1(new_n227), .A2(new_n228), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n212), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n215), .B(new_n223), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  NAND2_X1  g0043(.A1(new_n204), .A2(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n225), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT68), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n218), .B(new_n219), .C1(new_n212), .C2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n256));
  OR2_X1    g0056(.A1(new_n256), .A2(KEYINPUT70), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(KEYINPUT70), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  AOI211_X1 g0060(.A(new_n255), .B(new_n260), .C1(new_n209), .C2(G20), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G77), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G20), .A2(G77), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT8), .B(G58), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n210), .A2(G33), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT15), .B(G87), .ZN(new_n268));
  OAI221_X1 g0068(.A(new_n263), .B1(new_n264), .B2(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n255), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n262), .B(new_n270), .C1(G77), .C2(new_n259), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n218), .A2(new_n219), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n272), .B1(new_n254), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G33), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G1698), .ZN(new_n280));
  INV_X1    g0080(.A(G107), .ZN(new_n281));
  OAI22_X1  g0081(.A1(new_n280), .A2(new_n224), .B1(new_n281), .B2(new_n279), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n276), .A2(new_n278), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n283), .A2(new_n236), .A3(G1698), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n275), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(G274), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(G1), .B(G13), .C1(new_n254), .C2(new_n273), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n289), .A2(new_n286), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n288), .B1(new_n290), .B2(G244), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n271), .B1(G200), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(new_n292), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n271), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n292), .A2(G179), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT71), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g0102(.A(new_n302), .B(KEYINPUT72), .Z(new_n303));
  NAND3_X1  g0103(.A1(new_n279), .A2(G232), .A3(G1698), .ZN(new_n304));
  INV_X1    g0104(.A(G1698), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n279), .A2(G226), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G33), .A2(G97), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT73), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n304), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n275), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n288), .B1(new_n290), .B2(G238), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT74), .B(KEYINPUT13), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n313), .A2(new_n314), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT14), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(new_n318), .A3(G169), .ZN(new_n319));
  OAI21_X1  g0119(.A(G169), .B1(new_n315), .B2(new_n316), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT14), .ZN(new_n321));
  INV_X1    g0121(.A(new_n313), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n315), .B1(KEYINPUT13), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G179), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n319), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n225), .A2(G20), .ZN(new_n326));
  INV_X1    g0126(.A(G77), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n326), .B1(new_n267), .B2(new_n327), .C1(new_n266), .C2(new_n204), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n255), .A2(new_n328), .ZN(new_n329));
  XOR2_X1   g0129(.A(new_n329), .B(KEYINPUT11), .Z(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(G68), .B2(new_n261), .ZN(new_n331));
  XOR2_X1   g0131(.A(KEYINPUT75), .B(KEYINPUT12), .Z(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n259), .B2(G68), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT76), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n217), .A2(G1), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT12), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n334), .B1(new_n326), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n331), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n325), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n323), .A2(G190), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n317), .A2(G200), .ZN(new_n342));
  INV_X1    g0142(.A(new_n339), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n279), .A2(G222), .A3(new_n305), .ZN(new_n346));
  INV_X1    g0146(.A(G223), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n346), .B1(new_n327), .B2(new_n279), .C1(new_n280), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n275), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n288), .B1(new_n290), .B2(G226), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(G179), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n296), .B2(new_n351), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n205), .A2(G20), .ZN(new_n354));
  INV_X1    g0154(.A(G150), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n264), .B(KEYINPUT69), .ZN(new_n356));
  OAI221_X1 g0156(.A(new_n354), .B1(new_n355), .B2(new_n266), .C1(new_n356), .C2(new_n267), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n255), .ZN(new_n358));
  INV_X1    g0158(.A(new_n256), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n255), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n204), .B1(new_n209), .B2(G20), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n360), .A2(new_n361), .B1(new_n204), .B2(new_n359), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n353), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n363), .B(KEYINPUT9), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n351), .A2(new_n294), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(G200), .B2(new_n351), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT10), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT10), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n365), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NOR4_X1   g0172(.A1(new_n303), .A2(new_n345), .A3(new_n364), .A4(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n356), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(G1), .B2(new_n210), .ZN(new_n375));
  INV_X1    g0175(.A(new_n360), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n375), .A2(new_n376), .B1(new_n256), .B2(new_n374), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT77), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(KEYINPUT3), .B2(new_n254), .ZN(new_n379));
  NOR3_X1   g0179(.A1(new_n277), .A2(KEYINPUT77), .A3(G33), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n278), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT7), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(new_n382), .A3(new_n210), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT77), .B1(new_n277), .B2(G33), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n378), .A2(new_n254), .A3(KEYINPUT3), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT7), .B1(new_n387), .B2(G20), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n383), .A2(new_n388), .A3(G68), .ZN(new_n389));
  INV_X1    g0189(.A(G58), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n201), .B(new_n202), .C1(new_n390), .C2(new_n225), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n391), .A2(G20), .B1(G159), .B2(new_n265), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n389), .A2(KEYINPUT16), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT78), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT79), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n276), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n254), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n399), .A3(new_n278), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n382), .B1(new_n400), .B2(new_n210), .ZN(new_n401));
  AOI211_X1 g0201(.A(KEYINPUT7), .B(G20), .C1(new_n276), .C2(new_n278), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n401), .A2(new_n225), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n392), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n396), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n389), .A2(KEYINPUT78), .A3(KEYINPUT16), .A4(new_n392), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n395), .A2(new_n255), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT80), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n272), .B1(G33), .B2(new_n211), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n393), .B2(new_n394), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT80), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n410), .A2(new_n411), .A3(new_n405), .A4(new_n406), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n377), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n290), .A2(G232), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n287), .B2(new_n286), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n347), .A2(new_n305), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n387), .B(new_n416), .C1(G226), .C2(new_n305), .ZN(new_n417));
  INV_X1    g0217(.A(G87), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n417), .B1(new_n254), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n415), .B1(new_n419), .B2(new_n275), .ZN(new_n420));
  INV_X1    g0220(.A(G200), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(G190), .B2(new_n420), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n413), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT82), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(KEYINPUT82), .A2(KEYINPUT17), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n426), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n413), .A2(new_n428), .A3(new_n423), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT18), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n420), .A2(new_n296), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(G179), .B2(new_n420), .ZN(new_n434));
  NOR4_X1   g0234(.A1(new_n413), .A2(KEYINPUT81), .A3(new_n432), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n408), .A2(new_n412), .ZN(new_n436));
  INV_X1    g0236(.A(new_n377), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n434), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT18), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n438), .A2(KEYINPUT18), .A3(new_n439), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT81), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n431), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n445), .A2(new_n287), .A3(G1), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT5), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(KEYINPUT84), .B2(G41), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT84), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(new_n273), .A3(KEYINPUT5), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n446), .A2(new_n289), .A3(new_n448), .A4(new_n450), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT85), .ZN(new_n452));
  INV_X1    g0252(.A(G244), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(G1698), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT4), .B1(new_n387), .B2(new_n454), .ZN(new_n455));
  AND2_X1   g0255(.A1(KEYINPUT4), .A2(G244), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n276), .A2(new_n278), .A3(new_n456), .A4(new_n305), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n276), .A2(new_n278), .A3(G250), .A4(G1698), .ZN(new_n458));
  INV_X1    g0258(.A(G283), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n457), .B(new_n458), .C1(new_n254), .C2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n275), .B1(new_n455), .B2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n450), .A2(new_n448), .A3(new_n209), .A4(G45), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n289), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G257), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n452), .A2(new_n461), .A3(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(KEYINPUT86), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT86), .ZN(new_n468));
  OR2_X1    g0268(.A1(new_n451), .A2(KEYINPUT85), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n451), .A2(KEYINPUT85), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n469), .A2(new_n470), .B1(G257), .B2(new_n464), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n468), .B1(new_n471), .B2(new_n461), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n296), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n466), .ZN(new_n474));
  INV_X1    g0274(.A(G179), .ZN(new_n475));
  NOR3_X1   g0275(.A1(new_n401), .A2(new_n281), .A3(new_n402), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n265), .A2(G77), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n477), .B(KEYINPUT83), .ZN(new_n478));
  XNOR2_X1  g0278(.A(G97), .B(G107), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT6), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n281), .A2(KEYINPUT6), .A3(G97), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n478), .B1(new_n484), .B2(new_n210), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n255), .B1(new_n476), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n256), .A2(G97), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n254), .A2(G1), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n255), .A2(new_n359), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n487), .B1(new_n489), .B2(G97), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n474), .A2(new_n475), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n473), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(G250), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(new_n209), .B2(G45), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n446), .B1(new_n289), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(G238), .A2(G1698), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n496), .B1(new_n453), .B2(G1698), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n387), .A2(new_n497), .B1(G33), .B2(G116), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n495), .B1(new_n498), .B2(new_n274), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(G179), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(new_n296), .B2(new_n499), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n387), .A2(new_n210), .A3(G68), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT19), .ZN(new_n503));
  INV_X1    g0303(.A(G97), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n503), .B1(new_n267), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(G20), .B1(new_n308), .B2(KEYINPUT19), .ZN(new_n506));
  NOR3_X1   g0306(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n502), .B(new_n505), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n255), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n260), .A2(new_n268), .ZN(new_n510));
  OR3_X1    g0310(.A1(new_n255), .A2(new_n359), .A3(new_n488), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n509), .B(new_n510), .C1(new_n268), .C2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n499), .A2(new_n294), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(G200), .B2(new_n499), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n489), .A2(G87), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n509), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n501), .A2(new_n512), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n466), .A2(KEYINPUT86), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n471), .A2(new_n468), .A3(new_n461), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(G190), .A3(new_n519), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n486), .A2(new_n490), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n466), .A2(G200), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n492), .A2(new_n517), .A3(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n387), .A2(KEYINPUT22), .A3(new_n210), .A4(G87), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT22), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n210), .A2(G87), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n526), .B1(new_n283), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G116), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n254), .A2(new_n529), .A3(G20), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT23), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(new_n210), .B2(G107), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n281), .A2(KEYINPUT23), .A3(G20), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n525), .A2(new_n528), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT24), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT24), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n525), .A2(new_n537), .A3(new_n528), .A4(new_n534), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n255), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT88), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n359), .B(new_n281), .C1(new_n541), .C2(KEYINPUT25), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(KEYINPUT25), .ZN(new_n543));
  OR2_X1    g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n543), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n511), .B2(new_n281), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT89), .ZN(new_n550));
  MUX2_X1   g0350(.A(G250), .B(G257), .S(G1698), .Z(new_n551));
  AOI22_X1  g0351(.A1(new_n387), .A2(new_n551), .B1(G33), .B2(G294), .ZN(new_n552));
  INV_X1    g0352(.A(G264), .ZN(new_n553));
  OAI22_X1  g0353(.A1(new_n552), .A2(new_n274), .B1(new_n553), .B2(new_n463), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT85), .ZN(new_n555));
  XNOR2_X1  g0355(.A(new_n451), .B(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n296), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  OR2_X1    g0357(.A1(new_n552), .A2(new_n274), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n464), .A2(G264), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n558), .A2(new_n452), .A3(new_n475), .A4(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n549), .A2(new_n550), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n547), .B1(new_n539), .B2(new_n255), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n557), .A2(new_n560), .ZN(new_n564));
  OAI21_X1  g0364(.A(KEYINPUT89), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n558), .A2(new_n452), .A3(new_n559), .ZN(new_n566));
  OR2_X1    g0366(.A1(new_n566), .A2(new_n294), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(G200), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n563), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n562), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n469), .A2(new_n470), .B1(G270), .B2(new_n464), .ZN(new_n571));
  NOR2_X1   g0371(.A1(G257), .A2(G1698), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n553), .B2(G1698), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n387), .A2(new_n573), .B1(G303), .B2(new_n283), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT87), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n274), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n574), .A2(new_n575), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n571), .B(G190), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(G20), .B1(G33), .B2(G283), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n254), .A2(G97), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n580), .A2(new_n581), .B1(G20), .B2(new_n529), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n255), .A2(KEYINPUT20), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT20), .B1(new_n255), .B2(new_n582), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n260), .A2(new_n529), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n488), .A2(new_n529), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n409), .A2(new_n259), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n470), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n451), .A2(KEYINPUT85), .ZN(new_n593));
  INV_X1    g0393(.A(G270), .ZN(new_n594));
  OAI22_X1  g0394(.A1(new_n592), .A2(new_n593), .B1(new_n594), .B2(new_n463), .ZN(new_n595));
  INV_X1    g0395(.A(new_n578), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(new_n576), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n579), .B(new_n591), .C1(new_n597), .C2(new_n421), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n571), .B(G179), .C1(new_n577), .C2(new_n578), .ZN(new_n599));
  OR2_X1    g0399(.A1(new_n599), .A2(new_n591), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT21), .ZN(new_n601));
  OAI21_X1  g0401(.A(G169), .B1(new_n586), .B2(new_n590), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n597), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n590), .ZN(new_n604));
  INV_X1    g0404(.A(new_n585), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n583), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n296), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n571), .B1(new_n577), .B2(new_n578), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(KEYINPUT21), .A3(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n598), .A2(new_n600), .A3(new_n603), .A4(new_n609), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n524), .A2(new_n570), .A3(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n373), .A2(new_n444), .A3(new_n611), .ZN(G372));
  AOI21_X1  g0412(.A(new_n434), .B1(new_n436), .B2(new_n437), .ZN(new_n613));
  XNOR2_X1  g0413(.A(new_n613), .B(new_n432), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n340), .A2(new_n301), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n344), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n615), .B1(new_n617), .B2(new_n431), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n369), .A2(KEYINPUT90), .A3(new_n371), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT90), .B1(new_n369), .B2(new_n371), .ZN(new_n620));
  OR2_X1    g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n364), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n373), .A2(new_n444), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n517), .A2(new_n473), .A3(new_n491), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n624), .A2(KEYINPUT26), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(KEYINPUT26), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n501), .A2(new_n512), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n492), .A2(new_n517), .A3(new_n523), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n600), .A2(new_n603), .A3(new_n609), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n549), .A2(new_n561), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n631), .B(new_n569), .C1(new_n632), .C2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n622), .B1(new_n623), .B2(new_n637), .ZN(G369));
  AND3_X1   g0438(.A1(new_n562), .A2(new_n565), .A3(new_n569), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n335), .A2(new_n210), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(new_n642), .A3(G213), .ZN(new_n643));
  INV_X1    g0443(.A(G343), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n639), .B1(new_n563), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n633), .B2(new_n646), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n632), .A2(new_n646), .ZN(new_n649));
  XNOR2_X1  g0449(.A(new_n649), .B(KEYINPUT91), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n634), .B2(new_n646), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n591), .A2(new_n646), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n632), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n610), .B2(new_n653), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G330), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n648), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n652), .A2(new_n659), .ZN(G399));
  INV_X1    g0460(.A(new_n213), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(G41), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n507), .A2(new_n529), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n663), .A2(G1), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n222), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n666), .B1(new_n667), .B2(new_n663), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT28), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n625), .A2(new_n626), .A3(KEYINPUT95), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT95), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n624), .A2(new_n671), .A3(KEYINPUT26), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n631), .A2(new_n569), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n562), .A2(new_n565), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(new_n632), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n628), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n646), .B1(new_n673), .B2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n678), .A2(KEYINPUT29), .ZN(new_n679));
  AOI211_X1 g0479(.A(KEYINPUT29), .B(new_n645), .C1(new_n630), .C2(new_n635), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n467), .A2(new_n472), .ZN(new_n682));
  INV_X1    g0482(.A(new_n599), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n554), .A2(new_n499), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n682), .A2(KEYINPUT93), .A3(new_n683), .A4(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT93), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n518), .A2(new_n519), .A3(new_n684), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n686), .B1(new_n687), .B2(new_n599), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT30), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n682), .A2(KEYINPUT30), .A3(new_n683), .A4(new_n684), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n499), .A2(new_n475), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n608), .A2(new_n566), .A3(new_n466), .A4(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n690), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g0494(.A(KEYINPUT92), .B(KEYINPUT31), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n694), .A2(new_n645), .A3(new_n696), .ZN(new_n697));
  AND4_X1   g0497(.A1(new_n603), .A2(new_n598), .A3(new_n600), .A4(new_n609), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n631), .A2(new_n639), .A3(new_n698), .A4(new_n646), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n691), .A2(new_n693), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT94), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n700), .B1(new_n690), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n685), .A2(new_n688), .A3(KEYINPUT94), .A4(new_n689), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n646), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n697), .B(new_n699), .C1(new_n704), .C2(KEYINPUT31), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n681), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT96), .Z(new_n708));
  OAI21_X1  g0508(.A(new_n669), .B1(new_n708), .B2(G1), .ZN(G364));
  NOR2_X1   g0509(.A1(new_n217), .A2(G20), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n209), .B1(new_n710), .B2(G45), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n662), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n658), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(G330), .B2(new_n655), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n220), .B1(G20), .B2(new_n296), .ZN(new_n716));
  NOR2_X1   g0516(.A1(G13), .A2(G33), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G20), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n661), .A2(new_n387), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n248), .B2(new_n445), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n722), .B1(new_n445), .B2(new_n222), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n213), .A2(new_n279), .ZN(new_n724));
  INV_X1    g0524(.A(G355), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n724), .A2(new_n725), .B1(G116), .B2(new_n213), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n720), .B1(new_n723), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n713), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n421), .A2(G179), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n210), .A2(G190), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n283), .B1(new_n731), .B2(new_n459), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n210), .A2(new_n475), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G200), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G190), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  XOR2_X1   g0536(.A(KEYINPUT33), .B(G317), .Z(new_n737));
  INV_X1    g0537(.A(G294), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n294), .A2(G179), .A3(G200), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n210), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n736), .A2(new_n737), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n734), .A2(new_n294), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n732), .B(new_n741), .C1(G326), .C2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n729), .A2(G20), .A3(G190), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n744), .A2(KEYINPUT101), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(KEYINPUT101), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G303), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n730), .A2(new_n475), .A3(new_n421), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT99), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G329), .ZN(new_n756));
  INV_X1    g0556(.A(new_n733), .ZN(new_n757));
  AOI21_X1  g0557(.A(G200), .B1(new_n757), .B2(KEYINPUT97), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(KEYINPUT97), .B2(new_n757), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G190), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n294), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G311), .A2(new_n760), .B1(new_n761), .B2(G322), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n743), .A2(new_n749), .A3(new_n756), .A4(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n740), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G97), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(new_n736), .B2(new_n225), .ZN(new_n766));
  INV_X1    g0566(.A(new_n742), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n279), .B1(new_n731), .B2(new_n281), .C1(new_n767), .C2(new_n204), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n766), .B(new_n768), .C1(G87), .C2(new_n748), .ZN(new_n769));
  INV_X1    g0569(.A(G159), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n754), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(KEYINPUT100), .B(KEYINPUT32), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n771), .B(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n760), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n769), .B(new_n773), .C1(new_n327), .C2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n761), .B(KEYINPUT98), .Z(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n390), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n763), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n728), .B1(new_n778), .B2(new_n716), .ZN(new_n779));
  INV_X1    g0579(.A(new_n719), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n655), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n715), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(G396));
  INV_X1    g0583(.A(new_n301), .ZN(new_n784));
  AND3_X1   g0584(.A1(new_n784), .A2(KEYINPUT104), .A3(new_n645), .ZN(new_n785));
  AOI21_X1  g0585(.A(KEYINPUT104), .B1(new_n784), .B2(new_n645), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n271), .A2(new_n645), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n785), .A2(new_n786), .B1(new_n302), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(new_n637), .B2(new_n645), .ZN(new_n791));
  INV_X1    g0591(.A(new_n635), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n789), .B(new_n646), .C1(new_n629), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n713), .B1(new_n794), .B2(new_n706), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n706), .B2(new_n794), .ZN(new_n796));
  INV_X1    g0596(.A(new_n713), .ZN(new_n797));
  INV_X1    g0597(.A(new_n716), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n718), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT102), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n797), .B1(new_n801), .B2(new_n327), .ZN(new_n802));
  INV_X1    g0602(.A(new_n761), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n529), .A2(new_n774), .B1(new_n803), .B2(new_n738), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G283), .A2(new_n735), .B1(new_n742), .B2(G303), .ZN(new_n805));
  INV_X1    g0605(.A(new_n731), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n279), .B1(new_n806), .B2(G87), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n805), .A2(new_n765), .A3(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G311), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n281), .A2(new_n747), .B1(new_n754), .B2(new_n809), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n804), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(G137), .A2(new_n742), .B1(new_n735), .B2(G150), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT103), .ZN(new_n813));
  INV_X1    g0613(.A(G143), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n813), .B1(new_n770), .B2(new_n774), .C1(new_n776), .C2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT34), .ZN(new_n816));
  INV_X1    g0616(.A(G132), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n204), .A2(new_n747), .B1(new_n754), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n806), .A2(G68), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n819), .B(new_n387), .C1(new_n390), .C2(new_n740), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n811), .B1(new_n816), .B2(new_n821), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n802), .B1(new_n798), .B2(new_n822), .C1(new_n789), .C2(new_n718), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n796), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G384));
  NOR2_X1   g0625(.A1(new_n710), .A2(new_n209), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n410), .A2(new_n406), .ZN(new_n827));
  AOI21_X1  g0627(.A(KEYINPUT16), .B1(new_n389), .B2(new_n392), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n437), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n643), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT81), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n613), .A2(new_n832), .A3(KEYINPUT18), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n438), .A2(new_n439), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n432), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n443), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n427), .A2(new_n430), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n831), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT38), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n438), .A2(new_n830), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT37), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n834), .A2(new_n840), .A3(new_n841), .A4(new_n424), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n829), .B1(new_n439), .B2(new_n830), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n424), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT37), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n838), .A2(new_n839), .A3(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n831), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n832), .B1(new_n613), .B2(KEYINPUT18), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n850), .A2(new_n435), .A3(new_n440), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n849), .B1(new_n851), .B2(new_n431), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT38), .B1(new_n852), .B2(new_n846), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT39), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n840), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n614), .B2(new_n431), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n834), .A2(new_n840), .A3(new_n424), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT37), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n842), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g0660(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT39), .ZN(new_n863));
  OAI211_X1 g0663(.A(KEYINPUT38), .B(new_n846), .C1(new_n444), .C2(new_n831), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n854), .A2(KEYINPUT105), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n340), .A2(new_n645), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n839), .B1(new_n838), .B2(new_n847), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n864), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT105), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n869), .A2(new_n870), .A3(KEYINPUT39), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n866), .A2(new_n867), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n343), .A2(new_n646), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n325), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n345), .B2(new_n873), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n784), .A2(new_n646), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n876), .B1(new_n793), .B2(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n878), .A2(new_n869), .B1(new_n614), .B2(new_n643), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n872), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n444), .B(new_n373), .C1(new_n679), .C2(new_n680), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n622), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n880), .B(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n869), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n699), .A2(new_n696), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n704), .A2(new_n885), .ZN(new_n886));
  AOI211_X1 g0686(.A(KEYINPUT31), .B(new_n646), .C1(new_n702), .C2(new_n703), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT40), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(new_n789), .A4(new_n875), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n695), .B1(new_n611), .B2(new_n646), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n702), .A2(new_n703), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n891), .B1(new_n892), .B2(new_n646), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT31), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n704), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n893), .A2(new_n875), .A3(new_n789), .A4(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n862), .B2(new_n864), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n884), .A2(new_n890), .B1(new_n897), .B2(new_n889), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n623), .A2(new_n887), .A3(new_n886), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n657), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n899), .B2(new_n898), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n826), .B1(new_n883), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n883), .B2(new_n901), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n483), .A2(KEYINPUT35), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n483), .A2(KEYINPUT35), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n904), .A2(G116), .A3(new_n221), .A4(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT36), .ZN(new_n907));
  OAI21_X1  g0707(.A(G77), .B1(new_n390), .B2(new_n225), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n244), .B1(new_n667), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(G1), .A3(new_n217), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n903), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT107), .Z(G367));
  OAI21_X1  g0712(.A(new_n517), .B1(new_n516), .B2(new_n646), .ZN(new_n913));
  OR3_X1    g0713(.A1(new_n628), .A2(new_n516), .A3(new_n646), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n915), .A2(KEYINPUT108), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(KEYINPUT108), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT43), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(KEYINPUT43), .B2(new_n915), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n492), .B(new_n523), .C1(new_n521), .C2(new_n646), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n492), .B2(new_n646), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT109), .Z(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n651), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT110), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT42), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n922), .A2(new_n675), .ZN(new_n928));
  INV_X1    g0728(.A(new_n492), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n646), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n926), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  MUX2_X1   g0731(.A(new_n918), .B(new_n919), .S(new_n931), .Z(new_n932));
  AND3_X1   g0732(.A1(new_n922), .A2(new_n658), .A3(new_n648), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n652), .A2(new_n922), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT45), .Z(new_n936));
  NOR2_X1   g0736(.A1(new_n652), .A2(new_n922), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT44), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n659), .A2(KEYINPUT111), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n658), .B(new_n648), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(new_n650), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n708), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n708), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n662), .B(KEYINPUT41), .Z(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n934), .B1(new_n948), .B2(new_n712), .ZN(new_n949));
  INV_X1    g0749(.A(new_n721), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n720), .B1(new_n213), .B2(new_n268), .C1(new_n950), .C2(new_n242), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n951), .A2(KEYINPUT112), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(KEYINPUT112), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n952), .A2(new_n953), .A3(new_n797), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n767), .A2(new_n809), .B1(new_n281), .B2(new_n740), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(G294), .B2(new_n735), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n387), .B1(G97), .B2(new_n806), .ZN(new_n957));
  INV_X1    g0757(.A(G317), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n956), .B(new_n957), .C1(new_n958), .C2(new_n754), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(G283), .B2(new_n760), .ZN(new_n960));
  OAI21_X1  g0760(.A(KEYINPUT113), .B1(new_n747), .B2(new_n529), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT46), .Z(new_n962));
  INV_X1    g0762(.A(G303), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n960), .B(new_n962), .C1(new_n963), .C2(new_n776), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n806), .A2(G77), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n279), .B(new_n965), .C1(new_n736), .C2(new_n770), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n767), .A2(new_n814), .B1(new_n225), .B2(new_n740), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n755), .A2(G137), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n968), .B(new_n969), .C1(new_n390), .C2(new_n747), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n204), .A2(new_n774), .B1(new_n803), .B2(new_n355), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n964), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT47), .Z(new_n973));
  OAI221_X1 g0773(.A(new_n954), .B1(new_n780), .B2(new_n915), .C1(new_n973), .C2(new_n798), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n949), .A2(new_n974), .ZN(G387));
  OR2_X1    g0775(.A1(new_n648), .A2(new_n780), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n724), .A2(new_n665), .B1(G107), .B2(new_n213), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n239), .A2(new_n445), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n264), .A2(G50), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT50), .ZN(new_n980));
  AOI211_X1 g0780(.A(G45), .B(new_n664), .C1(G68), .C2(G77), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n950), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n977), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n720), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n713), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n747), .A2(new_n327), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n381), .B1(G97), .B2(new_n806), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(new_n355), .C2(new_n754), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT114), .ZN(new_n990));
  INV_X1    g0790(.A(new_n268), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n764), .A2(new_n991), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(new_n767), .B2(new_n770), .C1(new_n356), .C2(new_n736), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G50), .B2(new_n761), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n990), .B(new_n994), .C1(new_n225), .C2(new_n774), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G311), .A2(new_n735), .B1(new_n742), .B2(G322), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n963), .B2(new_n774), .C1(new_n776), .C2(new_n958), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(KEYINPUT48), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(KEYINPUT48), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n748), .A2(G294), .B1(G283), .B2(new_n764), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n381), .B1(new_n529), .B2(new_n731), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n755), .B2(G326), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT116), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n995), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n985), .B1(new_n1010), .B2(new_n716), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n943), .A2(new_n712), .B1(new_n976), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n944), .A2(new_n662), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n708), .A2(new_n943), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(G393));
  NAND3_X1  g0815(.A1(new_n939), .A2(new_n658), .A3(new_n648), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n936), .A2(new_n659), .A3(new_n938), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1018), .A2(new_n711), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n984), .B1(G97), .B2(new_n661), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n721), .A2(new_n252), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n797), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n761), .A2(G159), .B1(G150), .B2(new_n742), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT51), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n764), .A2(G77), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n204), .B2(new_n736), .C1(new_n774), .C2(new_n264), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n381), .B1(G87), .B2(new_n806), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n747), .B2(new_n225), .C1(new_n814), .C2(new_n754), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT117), .Z(new_n1030));
  AOI22_X1  g0830(.A1(new_n761), .A2(G311), .B1(G317), .B2(new_n742), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT52), .Z(new_n1032));
  AOI21_X1  g0832(.A(new_n279), .B1(new_n806), .B2(G107), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n529), .B2(new_n740), .C1(new_n736), .C2(new_n963), .ZN(new_n1034));
  INV_X1    g0834(.A(G322), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n459), .A2(new_n747), .B1(new_n754), .B2(new_n1035), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1034), .B(new_n1036), .C1(G294), .C2(new_n760), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1027), .A2(new_n1030), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1022), .B1(new_n798), .B2(new_n1038), .C1(new_n922), .C2(new_n780), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1019), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT118), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n944), .A2(new_n1018), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1044), .B(new_n662), .C1(new_n944), .C2(new_n941), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1045), .ZN(G390));
  NAND3_X1  g0846(.A1(new_n888), .A2(G330), .A3(new_n789), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1047), .A2(new_n876), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n878), .A2(new_n867), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n866), .B2(new_n871), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n789), .B(new_n646), .C1(new_n673), .C2(new_n677), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n877), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n867), .B1(new_n1052), .B2(new_n875), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n862), .A2(new_n864), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1048), .B1(new_n1050), .B2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n705), .A2(G330), .A3(new_n875), .A4(new_n789), .ZN(new_n1058));
  AOI211_X1 g0858(.A(KEYINPUT105), .B(new_n863), .C1(new_n868), .C2(new_n864), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n870), .B1(new_n869), .B2(KEYINPUT39), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1059), .B1(new_n1060), .B2(new_n865), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1058), .B(new_n1055), .C1(new_n1061), .C2(new_n1049), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1057), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n373), .A2(new_n888), .A3(G330), .A4(new_n444), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n881), .A2(new_n622), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n893), .A2(new_n789), .A3(new_n895), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n876), .B1(new_n1066), .B2(new_n657), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1067), .A2(new_n877), .A3(new_n1058), .A4(new_n1051), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n876), .B1(new_n706), .B2(new_n790), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n876), .B2(new_n1047), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n793), .A2(new_n877), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(KEYINPUT119), .A2(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1068), .A2(KEYINPUT119), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1065), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1063), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1057), .A2(new_n1062), .A3(new_n1074), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(new_n662), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1057), .A2(new_n712), .A3(new_n1062), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n504), .A2(new_n774), .B1(new_n803), .B2(new_n529), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G107), .A2(new_n735), .B1(new_n742), .B2(G283), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1081), .A2(new_n283), .A3(new_n819), .A4(new_n1025), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n418), .A2(new_n747), .B1(new_n754), .B2(new_n738), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n1080), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n735), .A2(G137), .ZN(new_n1085));
  INV_X1    g0885(.A(G128), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1085), .B1(new_n767), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G159), .B2(new_n764), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(KEYINPUT54), .B(G143), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1088), .B1(new_n774), .B2(new_n1089), .C1(new_n817), .C2(new_n803), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT53), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n747), .B2(new_n355), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n748), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1090), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n279), .B1(new_n731), .B2(new_n204), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n755), .B2(G125), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT120), .Z(new_n1097));
  AOI21_X1  g0897(.A(new_n1084), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n713), .B1(new_n374), .B2(new_n800), .C1(new_n1098), .C2(new_n798), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT121), .Z(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n1061), .B2(new_n718), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1078), .A2(new_n1079), .A3(new_n1101), .ZN(G378));
  INV_X1    g0902(.A(new_n364), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n619), .B2(new_n620), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n363), .A2(new_n830), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1103), .B(new_n1105), .C1(new_n619), .C2(new_n620), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1109), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n838), .A2(new_n847), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1113), .A2(KEYINPUT38), .B1(new_n860), .B2(new_n861), .ZN(new_n1114));
  OAI21_X1  g0914(.A(KEYINPUT40), .B1(new_n1114), .B2(new_n896), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n896), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n869), .A2(new_n889), .A3(new_n1116), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n657), .B(new_n1112), .C1(new_n1115), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1112), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n898), .B2(G330), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n880), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n889), .B1(new_n1054), .B2(new_n1116), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n890), .B1(new_n864), .B2(new_n868), .ZN(new_n1123));
  OAI21_X1  g0923(.A(G330), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n1112), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n898), .A2(G330), .A3(new_n1119), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1125), .A2(new_n872), .A3(new_n1126), .A4(new_n879), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1121), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n712), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n797), .B1(new_n801), .B2(new_n204), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n803), .A2(new_n1086), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G150), .A2(new_n764), .B1(new_n742), .B2(G125), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1132), .B1(new_n817), .B2(new_n736), .C1(new_n747), .C2(new_n1089), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(G137), .C2(new_n760), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1135), .A2(KEYINPUT59), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(KEYINPUT59), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n755), .A2(G124), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n254), .A2(new_n273), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n806), .B2(G159), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n740), .A2(new_n225), .B1(new_n731), .B2(new_n390), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n736), .A2(new_n504), .B1(new_n767), .B2(new_n529), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1142), .B(new_n1143), .C1(new_n991), .C2(new_n760), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n281), .B2(new_n803), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n986), .A2(G41), .A3(new_n387), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n459), .B2(new_n754), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n1148), .A2(KEYINPUT58), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(KEYINPUT58), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n204), .B(new_n1139), .C1(new_n387), .C2(G41), .ZN(new_n1151));
  AND4_X1   g0951(.A1(new_n1141), .A2(new_n1149), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1130), .B1(new_n798), .B2(new_n1152), .C1(new_n1119), .C2(new_n718), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1129), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1065), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1077), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n1128), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT57), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1158), .B1(new_n1121), .B2(new_n1127), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n663), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1154), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(G375));
  NAND3_X1  g0963(.A1(new_n1072), .A2(new_n1073), .A3(new_n1065), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1075), .A2(new_n947), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n381), .B1(G58), .B2(new_n806), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(new_n747), .B2(new_n770), .C1(new_n1086), .C2(new_n754), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1089), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G132), .A2(new_n742), .B1(new_n735), .B2(new_n1168), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n204), .B2(new_n740), .C1(new_n774), .C2(new_n355), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n776), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1167), .B(new_n1170), .C1(new_n1171), .C2(G137), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n281), .A2(new_n774), .B1(new_n803), .B2(new_n459), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G116), .A2(new_n735), .B1(new_n742), .B2(G294), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1174), .A2(new_n283), .A3(new_n965), .A4(new_n992), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n504), .A2(new_n747), .B1(new_n754), .B2(new_n963), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n1173), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n716), .B1(new_n1172), .B2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1178), .B(new_n713), .C1(G68), .C2(new_n800), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n876), .B2(new_n717), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1180), .B1(new_n1181), .B2(new_n712), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1165), .A2(new_n1182), .ZN(G381));
  NOR3_X1   g0983(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT122), .Z(new_n1185));
  NOR4_X1   g0985(.A1(new_n1185), .A2(G387), .A3(G390), .A4(G381), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(G375), .A2(G378), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(G407));
  NAND2_X1  g0988(.A1(new_n644), .A2(G213), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(G407), .A2(G213), .A3(new_n1191), .ZN(G409));
  AND2_X1   g0992(.A1(new_n949), .A2(new_n974), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(G390), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(G387), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT125), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n1193), .B2(G390), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(G393), .B(new_n782), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1196), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1194), .A2(new_n1197), .A3(new_n1195), .A4(new_n1199), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1203), .A2(KEYINPUT61), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1077), .A2(new_n1155), .B1(new_n1127), .B2(new_n1121), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1154), .B1(new_n947), .B2(new_n1205), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(G378), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT123), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1162), .B2(G378), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1156), .A2(new_n1160), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1210), .B(new_n662), .C1(KEYINPUT57), .C2(new_n1205), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1154), .ZN(new_n1212));
  AND4_X1   g1012(.A1(new_n1208), .A2(new_n1211), .A3(G378), .A4(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1207), .B1(new_n1209), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n1189), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1075), .A2(KEYINPUT60), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1216), .A2(new_n1164), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n662), .B1(new_n1216), .B2(new_n1164), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1182), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1219), .A2(new_n824), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n824), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT63), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1214), .A2(KEYINPUT124), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT124), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1226), .B(new_n1207), .C1(new_n1209), .C2(new_n1213), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1225), .A2(new_n1189), .A3(new_n1223), .A4(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT63), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1225), .A2(new_n1189), .A3(new_n1227), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1190), .A2(G2897), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1222), .B(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1230), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1204), .B1(new_n1215), .B2(new_n1224), .C1(new_n1229), .C2(new_n1234), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1233), .A2(new_n1215), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1236), .A2(KEYINPUT61), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT62), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1215), .A2(new_n1238), .A3(new_n1222), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1228), .A2(new_n1238), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1239), .B1(new_n1240), .B2(KEYINPUT126), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT126), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1228), .A2(new_n1242), .A3(new_n1238), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1237), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1203), .B(KEYINPUT127), .Z(new_n1245));
  OAI21_X1  g1045(.A(new_n1235), .B1(new_n1244), .B2(new_n1245), .ZN(G405));
  OAI22_X1  g1046(.A1(new_n1209), .A2(new_n1213), .B1(G378), .B2(new_n1162), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(new_n1223), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1203), .B(new_n1248), .ZN(G402));
endmodule


