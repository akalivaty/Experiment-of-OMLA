

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587;

  NOR2_X1 U325 ( .A1(n370), .A2(n369), .ZN(n371) );
  XNOR2_X1 U326 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U327 ( .A(KEYINPUT65), .B(n455), .Z(n293) );
  XOR2_X1 U328 ( .A(n409), .B(n408), .Z(n294) );
  XOR2_X1 U329 ( .A(G204GAT), .B(G92GAT), .Z(n295) );
  AND2_X1 U330 ( .A1(n511), .A2(n530), .ZN(n359) );
  XNOR2_X1 U331 ( .A(KEYINPUT25), .B(KEYINPUT90), .ZN(n361) );
  XNOR2_X1 U332 ( .A(n362), .B(n361), .ZN(n367) );
  INV_X1 U333 ( .A(KEYINPUT31), .ZN(n412) );
  NOR2_X1 U334 ( .A1(n367), .A2(n366), .ZN(n368) );
  XNOR2_X1 U335 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U336 ( .A(n464), .B(KEYINPUT54), .ZN(n465) );
  XNOR2_X1 U337 ( .A(KEYINPUT110), .B(KEYINPUT47), .ZN(n453) );
  XNOR2_X1 U338 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n319) );
  XNOR2_X1 U339 ( .A(n415), .B(n414), .ZN(n419) );
  XNOR2_X1 U340 ( .A(n454), .B(n453), .ZN(n461) );
  XNOR2_X1 U341 ( .A(n411), .B(n295), .ZN(n325) );
  NOR2_X1 U342 ( .A1(n506), .A2(n467), .ZN(n570) );
  XNOR2_X1 U343 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U344 ( .A(n388), .B(n387), .ZN(n452) );
  NOR2_X1 U345 ( .A1(n476), .A2(n505), .ZN(n442) );
  XNOR2_X1 U346 ( .A(n471), .B(KEYINPUT117), .ZN(n566) );
  XNOR2_X1 U347 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U348 ( .A(n446), .B(KEYINPUT108), .ZN(n447) );
  XNOR2_X1 U349 ( .A(n475), .B(n474), .ZN(G1349GAT) );
  XNOR2_X1 U350 ( .A(n448), .B(n447), .ZN(G1337GAT) );
  XOR2_X1 U351 ( .A(G85GAT), .B(G148GAT), .Z(n297) );
  XNOR2_X1 U352 ( .A(G134GAT), .B(G120GAT), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U354 ( .A(KEYINPUT86), .B(KEYINPUT6), .Z(n299) );
  XNOR2_X1 U355 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U357 ( .A(n301), .B(n300), .Z(n309) );
  XOR2_X1 U358 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n303) );
  XNOR2_X1 U359 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U361 ( .A(G141GAT), .B(n304), .Z(n334) );
  XOR2_X1 U362 ( .A(G57GAT), .B(KEYINPUT5), .Z(n306) );
  XNOR2_X1 U363 ( .A(KEYINPUT85), .B(KEYINPUT4), .ZN(n305) );
  XNOR2_X1 U364 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U365 ( .A(n334), .B(n307), .ZN(n308) );
  XNOR2_X1 U366 ( .A(n309), .B(n308), .ZN(n316) );
  XOR2_X1 U367 ( .A(G127GAT), .B(KEYINPUT0), .Z(n311) );
  XNOR2_X1 U368 ( .A(G113GAT), .B(KEYINPUT78), .ZN(n310) );
  XNOR2_X1 U369 ( .A(n311), .B(n310), .ZN(n353) );
  XOR2_X1 U370 ( .A(G162GAT), .B(n353), .Z(n313) );
  NAND2_X1 U371 ( .A1(G225GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U372 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U373 ( .A(G29GAT), .B(n314), .Z(n315) );
  XOR2_X1 U374 ( .A(n316), .B(n315), .Z(n443) );
  XOR2_X1 U375 ( .A(G36GAT), .B(G218GAT), .Z(n382) );
  XOR2_X1 U376 ( .A(G211GAT), .B(KEYINPUT21), .Z(n318) );
  XNOR2_X1 U377 ( .A(G197GAT), .B(KEYINPUT83), .ZN(n317) );
  XNOR2_X1 U378 ( .A(n318), .B(n317), .ZN(n340) );
  XOR2_X1 U379 ( .A(KEYINPUT87), .B(n340), .Z(n324) );
  XNOR2_X1 U380 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n320) );
  XNOR2_X1 U381 ( .A(n320), .B(n319), .ZN(n322) );
  XOR2_X1 U382 ( .A(G169GAT), .B(G190GAT), .Z(n321) );
  XNOR2_X1 U383 ( .A(n322), .B(n321), .ZN(n348) );
  XNOR2_X1 U384 ( .A(G8GAT), .B(n348), .ZN(n323) );
  XNOR2_X1 U385 ( .A(n324), .B(n323), .ZN(n326) );
  XOR2_X1 U386 ( .A(G176GAT), .B(G64GAT), .Z(n411) );
  XNOR2_X1 U387 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U388 ( .A(n382), .B(n327), .Z(n329) );
  NAND2_X1 U389 ( .A1(G226GAT), .A2(G233GAT), .ZN(n328) );
  XOR2_X2 U390 ( .A(n329), .B(n328), .Z(n511) );
  XOR2_X1 U391 ( .A(n511), .B(KEYINPUT88), .Z(n330) );
  XNOR2_X1 U392 ( .A(n330), .B(KEYINPUT27), .ZN(n364) );
  NOR2_X1 U393 ( .A1(n443), .A2(n364), .ZN(n544) );
  XOR2_X1 U394 ( .A(KEYINPUT82), .B(KEYINPUT23), .Z(n332) );
  XNOR2_X1 U395 ( .A(G22GAT), .B(G218GAT), .ZN(n331) );
  XNOR2_X1 U396 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U397 ( .A(n334), .B(n333), .ZN(n344) );
  XOR2_X1 U398 ( .A(G78GAT), .B(G148GAT), .Z(n336) );
  XNOR2_X1 U399 ( .A(G106GAT), .B(G204GAT), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n336), .B(n335), .ZN(n420) );
  XOR2_X1 U401 ( .A(G50GAT), .B(G162GAT), .Z(n381) );
  XOR2_X1 U402 ( .A(n420), .B(n381), .Z(n338) );
  NAND2_X1 U403 ( .A1(G228GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U404 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U405 ( .A(n339), .B(KEYINPUT22), .Z(n342) );
  XNOR2_X1 U406 ( .A(n340), .B(KEYINPUT24), .ZN(n341) );
  XNOR2_X1 U407 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n468) );
  XOR2_X1 U409 ( .A(n468), .B(KEYINPUT28), .Z(n517) );
  INV_X1 U410 ( .A(n517), .ZN(n524) );
  NAND2_X1 U411 ( .A1(n544), .A2(n524), .ZN(n529) );
  XOR2_X1 U412 ( .A(KEYINPUT64), .B(KEYINPUT79), .Z(n346) );
  XNOR2_X1 U413 ( .A(KEYINPUT80), .B(KEYINPUT20), .ZN(n345) );
  XNOR2_X1 U414 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U415 ( .A(n348), .B(n347), .ZN(n357) );
  XNOR2_X1 U416 ( .A(G43GAT), .B(G134GAT), .ZN(n385) );
  XNOR2_X1 U417 ( .A(G99GAT), .B(G71GAT), .ZN(n349) );
  XNOR2_X1 U418 ( .A(n349), .B(G120GAT), .ZN(n421) );
  XNOR2_X1 U419 ( .A(n385), .B(n421), .ZN(n351) );
  NAND2_X1 U420 ( .A1(G227GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U421 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U422 ( .A(n352), .B(G176GAT), .Z(n355) );
  XNOR2_X1 U423 ( .A(G15GAT), .B(n353), .ZN(n354) );
  XNOR2_X1 U424 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U425 ( .A(n357), .B(n356), .Z(n522) );
  XNOR2_X1 U426 ( .A(n522), .B(KEYINPUT81), .ZN(n358) );
  NOR2_X1 U427 ( .A1(n529), .A2(n358), .ZN(n370) );
  INV_X1 U428 ( .A(n522), .ZN(n530) );
  XNOR2_X1 U429 ( .A(n359), .B(KEYINPUT89), .ZN(n360) );
  NAND2_X1 U430 ( .A1(n360), .A2(n468), .ZN(n362) );
  NOR2_X1 U431 ( .A1(n530), .A2(n468), .ZN(n363) );
  XNOR2_X1 U432 ( .A(KEYINPUT26), .B(n363), .ZN(n569) );
  INV_X1 U433 ( .A(n569), .ZN(n365) );
  NOR2_X1 U434 ( .A1(n365), .A2(n364), .ZN(n366) );
  INV_X1 U435 ( .A(n443), .ZN(n506) );
  NOR2_X1 U436 ( .A1(n368), .A2(n506), .ZN(n369) );
  XNOR2_X1 U437 ( .A(n371), .B(KEYINPUT91), .ZN(n483) );
  INV_X1 U438 ( .A(n483), .ZN(n389) );
  XOR2_X1 U439 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n373) );
  XNOR2_X1 U440 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U442 ( .A(n374), .B(G99GAT), .Z(n377) );
  XNOR2_X1 U443 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n375) );
  XNOR2_X1 U444 ( .A(n375), .B(KEYINPUT7), .ZN(n433) );
  XNOR2_X1 U445 ( .A(n433), .B(G190GAT), .ZN(n376) );
  XNOR2_X1 U446 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U447 ( .A(G85GAT), .B(G92GAT), .Z(n408) );
  XNOR2_X1 U448 ( .A(n378), .B(n408), .ZN(n380) );
  XOR2_X1 U449 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n379) );
  XNOR2_X1 U450 ( .A(n380), .B(n379), .ZN(n388) );
  XOR2_X1 U451 ( .A(n382), .B(n381), .Z(n384) );
  NAND2_X1 U452 ( .A1(G232GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U453 ( .A(n384), .B(n383), .ZN(n386) );
  INV_X1 U454 ( .A(n452), .ZN(n565) );
  XOR2_X1 U455 ( .A(KEYINPUT36), .B(n565), .Z(n584) );
  NOR2_X1 U456 ( .A1(n389), .A2(n584), .ZN(n406) );
  XOR2_X1 U457 ( .A(G8GAT), .B(G1GAT), .Z(n391) );
  XNOR2_X1 U458 ( .A(G15GAT), .B(G22GAT), .ZN(n390) );
  XNOR2_X1 U459 ( .A(n391), .B(n390), .ZN(n432) );
  XNOR2_X1 U460 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n392) );
  XNOR2_X1 U461 ( .A(KEYINPUT72), .B(n392), .ZN(n409) );
  XOR2_X1 U462 ( .A(n432), .B(n409), .Z(n405) );
  XOR2_X1 U463 ( .A(KEYINPUT15), .B(KEYINPUT77), .Z(n394) );
  NAND2_X1 U464 ( .A1(G231GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U465 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U466 ( .A(n395), .B(KEYINPUT12), .Z(n403) );
  XOR2_X1 U467 ( .A(G211GAT), .B(G71GAT), .Z(n397) );
  XNOR2_X1 U468 ( .A(G183GAT), .B(G127GAT), .ZN(n396) );
  XNOR2_X1 U469 ( .A(n397), .B(n396), .ZN(n401) );
  XOR2_X1 U470 ( .A(KEYINPUT14), .B(G64GAT), .Z(n399) );
  XNOR2_X1 U471 ( .A(G155GAT), .B(G78GAT), .ZN(n398) );
  XNOR2_X1 U472 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U473 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U474 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U475 ( .A(n405), .B(n404), .Z(n579) );
  NAND2_X1 U476 ( .A1(n406), .A2(n579), .ZN(n407) );
  XOR2_X1 U477 ( .A(n407), .B(KEYINPUT37), .Z(n476) );
  NAND2_X1 U478 ( .A1(G230GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U479 ( .A(n294), .B(n410), .ZN(n415) );
  XNOR2_X1 U480 ( .A(n411), .B(KEYINPUT74), .ZN(n413) );
  XOR2_X1 U481 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n417) );
  XNOR2_X1 U482 ( .A(KEYINPUT73), .B(KEYINPUT75), .ZN(n416) );
  XNOR2_X1 U483 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U484 ( .A(n419), .B(n418), .Z(n423) );
  XNOR2_X1 U485 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n575) );
  XOR2_X1 U487 ( .A(n575), .B(KEYINPUT41), .Z(n549) );
  XOR2_X1 U488 ( .A(n549), .B(KEYINPUT100), .Z(n534) );
  XOR2_X1 U489 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n425) );
  XNOR2_X1 U490 ( .A(G141GAT), .B(KEYINPUT68), .ZN(n424) );
  XNOR2_X1 U491 ( .A(n425), .B(n424), .ZN(n441) );
  XOR2_X1 U492 ( .A(G197GAT), .B(G113GAT), .Z(n427) );
  XNOR2_X1 U493 ( .A(G169GAT), .B(G36GAT), .ZN(n426) );
  XNOR2_X1 U494 ( .A(n427), .B(n426), .ZN(n429) );
  XOR2_X1 U495 ( .A(G50GAT), .B(G43GAT), .Z(n428) );
  XNOR2_X1 U496 ( .A(n429), .B(n428), .ZN(n437) );
  XNOR2_X1 U497 ( .A(KEYINPUT71), .B(KEYINPUT69), .ZN(n430) );
  XNOR2_X1 U498 ( .A(n430), .B(KEYINPUT67), .ZN(n431) );
  XOR2_X1 U499 ( .A(n431), .B(KEYINPUT70), .Z(n435) );
  XNOR2_X1 U500 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U501 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U502 ( .A(n437), .B(n436), .ZN(n439) );
  NAND2_X1 U503 ( .A1(G229GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U504 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U505 ( .A(n441), .B(n440), .ZN(n571) );
  NAND2_X1 U506 ( .A1(n534), .A2(n571), .ZN(n505) );
  XOR2_X1 U507 ( .A(KEYINPUT106), .B(n442), .Z(n525) );
  NOR2_X1 U508 ( .A1(n443), .A2(n525), .ZN(n445) );
  XNOR2_X1 U509 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n444) );
  XNOR2_X1 U510 ( .A(n445), .B(n444), .ZN(G1336GAT) );
  INV_X1 U511 ( .A(n511), .ZN(n463) );
  NOR2_X1 U512 ( .A1(n525), .A2(n463), .ZN(n448) );
  INV_X1 U513 ( .A(G92GAT), .ZN(n446) );
  INV_X1 U514 ( .A(n579), .ZN(n560) );
  NOR2_X1 U515 ( .A1(n549), .A2(n571), .ZN(n449) );
  XNOR2_X1 U516 ( .A(n449), .B(KEYINPUT46), .ZN(n450) );
  NOR2_X1 U517 ( .A1(n560), .A2(n450), .ZN(n451) );
  NAND2_X1 U518 ( .A1(n452), .A2(n451), .ZN(n454) );
  INV_X1 U519 ( .A(n571), .ZN(n556) );
  NOR2_X1 U520 ( .A1(n579), .A2(n584), .ZN(n456) );
  XOR2_X1 U521 ( .A(KEYINPUT111), .B(KEYINPUT45), .Z(n455) );
  XNOR2_X1 U522 ( .A(n456), .B(n293), .ZN(n457) );
  NAND2_X1 U523 ( .A1(n457), .A2(n575), .ZN(n458) );
  NOR2_X1 U524 ( .A1(n556), .A2(n458), .ZN(n459) );
  XNOR2_X1 U525 ( .A(KEYINPUT112), .B(n459), .ZN(n460) );
  NOR2_X1 U526 ( .A1(n461), .A2(n460), .ZN(n462) );
  XNOR2_X1 U527 ( .A(KEYINPUT48), .B(n462), .ZN(n546) );
  NOR2_X1 U528 ( .A1(n463), .A2(n546), .ZN(n466) );
  INV_X1 U529 ( .A(KEYINPUT116), .ZN(n464) );
  NAND2_X1 U530 ( .A1(n468), .A2(n570), .ZN(n469) );
  XNOR2_X1 U531 ( .A(KEYINPUT55), .B(n469), .ZN(n470) );
  NAND2_X1 U532 ( .A1(n470), .A2(n530), .ZN(n471) );
  NAND2_X1 U533 ( .A1(n566), .A2(n534), .ZN(n475) );
  XOR2_X1 U534 ( .A(G176GAT), .B(KEYINPUT56), .Z(n473) );
  XNOR2_X1 U535 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n472) );
  XOR2_X1 U536 ( .A(KEYINPUT95), .B(KEYINPUT39), .Z(n479) );
  NAND2_X1 U537 ( .A1(n556), .A2(n575), .ZN(n485) );
  NOR2_X1 U538 ( .A1(n476), .A2(n485), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n477), .B(KEYINPUT38), .ZN(n502) );
  NAND2_X1 U540 ( .A1(n502), .A2(n506), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n479), .B(n478), .ZN(n481) );
  INV_X1 U542 ( .A(G29GAT), .ZN(n480) );
  XNOR2_X1 U543 ( .A(n481), .B(n480), .ZN(G1328GAT) );
  NOR2_X1 U544 ( .A1(n565), .A2(n579), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n482), .B(KEYINPUT16), .ZN(n484) );
  NAND2_X1 U546 ( .A1(n484), .A2(n483), .ZN(n504) );
  NOR2_X1 U547 ( .A1(n485), .A2(n504), .ZN(n493) );
  NAND2_X1 U548 ( .A1(n506), .A2(n493), .ZN(n488) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n486), .B(KEYINPUT92), .ZN(n487) );
  XNOR2_X1 U551 ( .A(n488), .B(n487), .ZN(G1324GAT) );
  XOR2_X1 U552 ( .A(G8GAT), .B(KEYINPUT93), .Z(n490) );
  NAND2_X1 U553 ( .A1(n493), .A2(n511), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n490), .B(n489), .ZN(G1325GAT) );
  XOR2_X1 U555 ( .A(G15GAT), .B(KEYINPUT35), .Z(n492) );
  NAND2_X1 U556 ( .A1(n493), .A2(n530), .ZN(n491) );
  XNOR2_X1 U557 ( .A(n492), .B(n491), .ZN(G1326GAT) );
  NAND2_X1 U558 ( .A1(n493), .A2(n517), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n494), .B(KEYINPUT94), .ZN(n495) );
  XNOR2_X1 U560 ( .A(G22GAT), .B(n495), .ZN(G1327GAT) );
  NAND2_X1 U561 ( .A1(n511), .A2(n502), .ZN(n496) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(n496), .ZN(G1329GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT40), .B(KEYINPUT98), .Z(n498) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(KEYINPUT97), .ZN(n497) );
  XNOR2_X1 U565 ( .A(n498), .B(n497), .ZN(n501) );
  NAND2_X1 U566 ( .A1(n502), .A2(n530), .ZN(n499) );
  XNOR2_X1 U567 ( .A(n499), .B(KEYINPUT96), .ZN(n500) );
  XNOR2_X1 U568 ( .A(n501), .B(n500), .ZN(G1330GAT) );
  NAND2_X1 U569 ( .A1(n502), .A2(n517), .ZN(n503) );
  XNOR2_X1 U570 ( .A(n503), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U571 ( .A(G57GAT), .B(KEYINPUT99), .Z(n508) );
  NOR2_X1 U572 ( .A1(n505), .A2(n504), .ZN(n518) );
  NAND2_X1 U573 ( .A1(n518), .A2(n506), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(n510) );
  XOR2_X1 U575 ( .A(KEYINPUT42), .B(KEYINPUT101), .Z(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1332GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n513) );
  NAND2_X1 U578 ( .A1(n518), .A2(n511), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G64GAT), .B(n514), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n518), .A2(n530), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n515), .B(KEYINPUT104), .ZN(n516) );
  XNOR2_X1 U583 ( .A(G71GAT), .B(n516), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n520) );
  NAND2_X1 U585 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U587 ( .A(G78GAT), .B(n521), .Z(G1335GAT) );
  NOR2_X1 U588 ( .A1(n525), .A2(n522), .ZN(n523) );
  XOR2_X1 U589 ( .A(G99GAT), .B(n523), .Z(G1338GAT) );
  NOR2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n527) );
  XNOR2_X1 U591 ( .A(KEYINPUT109), .B(KEYINPUT44), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NOR2_X1 U594 ( .A1(n546), .A2(n529), .ZN(n531) );
  NAND2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n532), .B(KEYINPUT113), .ZN(n540) );
  NAND2_X1 U597 ( .A1(n540), .A2(n556), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n533), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U600 ( .A1(n540), .A2(n534), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U602 ( .A(G120GAT), .B(n537), .ZN(G1341GAT) );
  NAND2_X1 U603 ( .A1(n560), .A2(n540), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n538), .B(KEYINPUT50), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U607 ( .A1(n540), .A2(n565), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U609 ( .A(G134GAT), .B(n543), .Z(G1343GAT) );
  NAND2_X1 U610 ( .A1(n544), .A2(n569), .ZN(n545) );
  NOR2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n554), .A2(n556), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n547), .B(G141GAT), .ZN(G1344GAT) );
  INV_X1 U614 ( .A(n554), .ZN(n548) );
  NOR2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n551) );
  XNOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(n552), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n560), .A2(n554), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n554), .A2(n565), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U623 ( .A1(n566), .A2(n556), .ZN(n559) );
  XOR2_X1 U624 ( .A(G169GAT), .B(KEYINPUT118), .Z(n557) );
  XNOR2_X1 U625 ( .A(KEYINPUT119), .B(n557), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1348GAT) );
  XOR2_X1 U627 ( .A(G183GAT), .B(KEYINPUT121), .Z(n562) );
  NAND2_X1 U628 ( .A1(n566), .A2(n560), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1350GAT) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n563), .B(KEYINPUT122), .ZN(n564) );
  XOR2_X1 U632 ( .A(KEYINPUT123), .B(n564), .Z(n568) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1351GAT) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n583) );
  NOR2_X1 U636 ( .A1(n571), .A2(n583), .ZN(n573) );
  XNOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(n574), .ZN(G1352GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n583), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT124), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n578), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n583), .ZN(n581) );
  XNOR2_X1 U645 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(n582), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

