

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591;

  XNOR2_X1 U323 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U324 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n514) );
  XNOR2_X1 U325 ( .A(n374), .B(n342), .ZN(n345) );
  XNOR2_X1 U326 ( .A(n515), .B(n514), .ZN(n547) );
  NOR2_X1 U327 ( .A1(n557), .A2(n556), .ZN(n567) );
  XOR2_X1 U328 ( .A(KEYINPUT94), .B(KEYINPUT34), .Z(n292) );
  XNOR2_X1 U329 ( .A(G1GAT), .B(KEYINPUT95), .ZN(n291) );
  XNOR2_X1 U330 ( .A(n292), .B(n291), .ZN(n452) );
  XOR2_X1 U331 ( .A(G120GAT), .B(G148GAT), .Z(n341) );
  XOR2_X1 U332 ( .A(G57GAT), .B(G85GAT), .Z(n294) );
  XNOR2_X1 U333 ( .A(G29GAT), .B(G141GAT), .ZN(n293) );
  XNOR2_X1 U334 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U335 ( .A(n341), .B(n295), .Z(n297) );
  NAND2_X1 U336 ( .A1(G225GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U337 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U338 ( .A(n298), .B(KEYINPUT87), .Z(n302) );
  XOR2_X1 U339 ( .A(KEYINPUT0), .B(KEYINPUT82), .Z(n300) );
  XNOR2_X1 U340 ( .A(G113GAT), .B(G134GAT), .ZN(n299) );
  XNOR2_X1 U341 ( .A(n300), .B(n299), .ZN(n355) );
  XNOR2_X1 U342 ( .A(n355), .B(KEYINPUT1), .ZN(n301) );
  XNOR2_X1 U343 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U344 ( .A(KEYINPUT88), .B(KEYINPUT4), .Z(n304) );
  XNOR2_X1 U345 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n303) );
  XNOR2_X1 U346 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U347 ( .A(n306), .B(n305), .Z(n310) );
  XNOR2_X1 U348 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n307) );
  XNOR2_X1 U349 ( .A(n307), .B(KEYINPUT3), .ZN(n392) );
  XNOR2_X1 U350 ( .A(G1GAT), .B(G127GAT), .ZN(n308) );
  XNOR2_X1 U351 ( .A(n308), .B(G155GAT), .ZN(n446) );
  XNOR2_X1 U352 ( .A(n392), .B(n446), .ZN(n309) );
  XNOR2_X1 U353 ( .A(n310), .B(n309), .ZN(n411) );
  XNOR2_X1 U354 ( .A(KEYINPUT89), .B(n411), .ZN(n491) );
  XOR2_X1 U355 ( .A(KEYINPUT72), .B(KEYINPUT68), .Z(n312) );
  XNOR2_X1 U356 ( .A(KEYINPUT69), .B(KEYINPUT30), .ZN(n311) );
  XNOR2_X1 U357 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U358 ( .A(G197GAT), .B(G113GAT), .Z(n314) );
  XOR2_X1 U359 ( .A(G50GAT), .B(G141GAT), .Z(n396) );
  XOR2_X1 U360 ( .A(G169GAT), .B(G36GAT), .Z(n378) );
  XNOR2_X1 U361 ( .A(n396), .B(n378), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U363 ( .A(n316), .B(n315), .Z(n318) );
  NAND2_X1 U364 ( .A1(G229GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U366 ( .A(KEYINPUT71), .B(KEYINPUT29), .Z(n320) );
  XNOR2_X1 U367 ( .A(G1GAT), .B(G8GAT), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U369 ( .A(n322), .B(n321), .Z(n331) );
  INV_X1 U370 ( .A(G43GAT), .ZN(n323) );
  NAND2_X1 U371 ( .A1(G29GAT), .A2(n323), .ZN(n326) );
  INV_X1 U372 ( .A(G29GAT), .ZN(n324) );
  NAND2_X1 U373 ( .A1(n324), .A2(G43GAT), .ZN(n325) );
  NAND2_X1 U374 ( .A1(n326), .A2(n325), .ZN(n328) );
  XNOR2_X1 U375 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n327) );
  XNOR2_X1 U376 ( .A(n328), .B(n327), .ZN(n414) );
  XNOR2_X1 U377 ( .A(G15GAT), .B(G22GAT), .ZN(n329) );
  XNOR2_X1 U378 ( .A(n329), .B(KEYINPUT70), .ZN(n438) );
  XNOR2_X1 U379 ( .A(n414), .B(n438), .ZN(n330) );
  XNOR2_X1 U380 ( .A(n331), .B(n330), .ZN(n576) );
  XNOR2_X1 U381 ( .A(KEYINPUT73), .B(n576), .ZN(n558) );
  INV_X1 U382 ( .A(n558), .ZN(n510) );
  INV_X1 U383 ( .A(G204GAT), .ZN(n339) );
  INV_X1 U384 ( .A(KEYINPUT76), .ZN(n332) );
  NAND2_X1 U385 ( .A1(n332), .A2(G92GAT), .ZN(n335) );
  INV_X1 U386 ( .A(G92GAT), .ZN(n333) );
  NAND2_X1 U387 ( .A1(n333), .A2(KEYINPUT76), .ZN(n334) );
  NAND2_X1 U388 ( .A1(n335), .A2(n334), .ZN(n337) );
  XNOR2_X1 U389 ( .A(G176GAT), .B(G64GAT), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n339), .B(n338), .ZN(n374) );
  XOR2_X1 U392 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n340) );
  XOR2_X1 U393 ( .A(KEYINPUT13), .B(KEYINPUT74), .Z(n344) );
  XNOR2_X1 U394 ( .A(G71GAT), .B(G57GAT), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n344), .B(n343), .ZN(n437) );
  XOR2_X1 U396 ( .A(n345), .B(n437), .Z(n347) );
  XOR2_X1 U397 ( .A(G106GAT), .B(G78GAT), .Z(n390) );
  XOR2_X1 U398 ( .A(G99GAT), .B(G85GAT), .Z(n419) );
  XNOR2_X1 U399 ( .A(n390), .B(n419), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n347), .B(n346), .ZN(n352) );
  XOR2_X1 U401 ( .A(KEYINPUT77), .B(KEYINPUT31), .Z(n349) );
  NAND2_X1 U402 ( .A1(G230GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U404 ( .A(KEYINPUT75), .B(n350), .Z(n351) );
  XNOR2_X1 U405 ( .A(n352), .B(n351), .ZN(n579) );
  NOR2_X1 U406 ( .A1(n510), .A2(n579), .ZN(n463) );
  XOR2_X1 U407 ( .A(G190GAT), .B(G99GAT), .Z(n354) );
  NAND2_X1 U408 ( .A1(G227GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n356) );
  XOR2_X1 U410 ( .A(n356), .B(n355), .Z(n364) );
  XOR2_X1 U411 ( .A(G183GAT), .B(KEYINPUT83), .Z(n358) );
  XNOR2_X1 U412 ( .A(G43GAT), .B(KEYINPUT20), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U414 ( .A(G71GAT), .B(G176GAT), .Z(n360) );
  XNOR2_X1 U415 ( .A(G169GAT), .B(G15GAT), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U417 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U418 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U419 ( .A(n365), .B(G120GAT), .Z(n369) );
  XOR2_X1 U420 ( .A(KEYINPUT17), .B(KEYINPUT84), .Z(n367) );
  XNOR2_X1 U421 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n367), .B(n366), .ZN(n370) );
  XNOR2_X1 U423 ( .A(n370), .B(G127GAT), .ZN(n368) );
  XOR2_X1 U424 ( .A(n369), .B(n368), .Z(n470) );
  XOR2_X1 U425 ( .A(KEYINPUT90), .B(n370), .Z(n372) );
  NAND2_X1 U426 ( .A1(G226GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U428 ( .A(n374), .B(n373), .ZN(n382) );
  XNOR2_X1 U429 ( .A(G8GAT), .B(G183GAT), .ZN(n375) );
  XNOR2_X1 U430 ( .A(n375), .B(G211GAT), .ZN(n445) );
  XOR2_X1 U431 ( .A(G190GAT), .B(KEYINPUT79), .Z(n418) );
  XOR2_X1 U432 ( .A(n445), .B(n418), .Z(n380) );
  XOR2_X1 U433 ( .A(KEYINPUT85), .B(KEYINPUT21), .Z(n377) );
  XNOR2_X1 U434 ( .A(G197GAT), .B(G218GAT), .ZN(n376) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n391) );
  XNOR2_X1 U436 ( .A(n378), .B(n391), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U438 ( .A(n382), .B(n381), .Z(n493) );
  XOR2_X1 U439 ( .A(n493), .B(KEYINPUT91), .Z(n383) );
  XNOR2_X1 U440 ( .A(n383), .B(KEYINPUT27), .ZN(n406) );
  NOR2_X1 U441 ( .A1(n406), .A2(n491), .ZN(n516) );
  XOR2_X1 U442 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n385) );
  XNOR2_X1 U443 ( .A(KEYINPUT86), .B(KEYINPUT24), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U445 ( .A(G148GAT), .B(G155GAT), .Z(n387) );
  XNOR2_X1 U446 ( .A(G211GAT), .B(G204GAT), .ZN(n386) );
  XNOR2_X1 U447 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n400) );
  XOR2_X1 U449 ( .A(n391), .B(n390), .Z(n398) );
  XOR2_X1 U450 ( .A(G22GAT), .B(n392), .Z(n394) );
  NAND2_X1 U451 ( .A1(G228GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U453 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n400), .B(n399), .ZN(n554) );
  XNOR2_X1 U456 ( .A(n554), .B(KEYINPUT28), .ZN(n474) );
  INV_X1 U457 ( .A(n474), .ZN(n519) );
  NAND2_X1 U458 ( .A1(n516), .A2(n519), .ZN(n401) );
  NOR2_X1 U459 ( .A1(n470), .A2(n401), .ZN(n402) );
  XNOR2_X1 U460 ( .A(KEYINPUT92), .B(n402), .ZN(n413) );
  INV_X1 U461 ( .A(n470), .ZN(n557) );
  NOR2_X1 U462 ( .A1(n557), .A2(n493), .ZN(n403) );
  NOR2_X1 U463 ( .A1(n554), .A2(n403), .ZN(n404) );
  XOR2_X1 U464 ( .A(KEYINPUT25), .B(n404), .Z(n409) );
  NAND2_X1 U465 ( .A1(n554), .A2(n557), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n405), .B(KEYINPUT26), .ZN(n574) );
  NOR2_X1 U467 ( .A1(n574), .A2(n406), .ZN(n407) );
  XOR2_X1 U468 ( .A(KEYINPUT93), .B(n407), .Z(n408) );
  NOR2_X1 U469 ( .A1(n409), .A2(n408), .ZN(n410) );
  NOR2_X1 U470 ( .A1(n411), .A2(n410), .ZN(n412) );
  NOR2_X1 U471 ( .A1(n413), .A2(n412), .ZN(n460) );
  INV_X1 U472 ( .A(G50GAT), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n417) );
  NAND2_X1 U474 ( .A1(G232GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n417), .B(n416), .ZN(n423) );
  XOR2_X1 U476 ( .A(KEYINPUT11), .B(n418), .Z(n421) );
  XNOR2_X1 U477 ( .A(G92GAT), .B(n419), .ZN(n420) );
  XOR2_X1 U478 ( .A(n421), .B(n420), .Z(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n425) );
  XNOR2_X1 U480 ( .A(G36GAT), .B(G218GAT), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n433) );
  XOR2_X1 U482 ( .A(KEYINPUT9), .B(G106GAT), .Z(n427) );
  XNOR2_X1 U483 ( .A(G134GAT), .B(G162GAT), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U485 ( .A(KEYINPUT67), .B(KEYINPUT78), .Z(n429) );
  XNOR2_X1 U486 ( .A(KEYINPUT10), .B(KEYINPUT66), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U488 ( .A(n431), .B(n430), .Z(n432) );
  XOR2_X1 U489 ( .A(n433), .B(n432), .Z(n568) );
  XOR2_X1 U490 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n435) );
  NAND2_X1 U491 ( .A1(G231GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U493 ( .A(n436), .B(KEYINPUT12), .Z(n440) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U496 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n442) );
  XNOR2_X1 U497 ( .A(G78GAT), .B(G64GAT), .ZN(n441) );
  XNOR2_X1 U498 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U499 ( .A(n444), .B(n443), .Z(n448) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n448), .B(n447), .ZN(n583) );
  NOR2_X1 U502 ( .A1(n568), .A2(n583), .ZN(n449) );
  XOR2_X1 U503 ( .A(KEYINPUT16), .B(n449), .Z(n450) );
  NOR2_X1 U504 ( .A1(n460), .A2(n450), .ZN(n479) );
  NAND2_X1 U505 ( .A1(n463), .A2(n479), .ZN(n457) );
  NOR2_X1 U506 ( .A1(n491), .A2(n457), .ZN(n451) );
  XOR2_X1 U507 ( .A(n452), .B(n451), .Z(G1324GAT) );
  NOR2_X1 U508 ( .A1(n493), .A2(n457), .ZN(n453) );
  XOR2_X1 U509 ( .A(G8GAT), .B(n453), .Z(G1325GAT) );
  NOR2_X1 U510 ( .A1(n557), .A2(n457), .ZN(n455) );
  XNOR2_X1 U511 ( .A(KEYINPUT35), .B(KEYINPUT96), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U513 ( .A(G15GAT), .B(n456), .ZN(G1326GAT) );
  NOR2_X1 U514 ( .A1(n519), .A2(n457), .ZN(n459) );
  XNOR2_X1 U515 ( .A(G22GAT), .B(KEYINPUT97), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n459), .B(n458), .ZN(G1327GAT) );
  XOR2_X1 U517 ( .A(KEYINPUT99), .B(KEYINPUT39), .Z(n467) );
  XOR2_X1 U518 ( .A(KEYINPUT38), .B(KEYINPUT98), .Z(n465) );
  XOR2_X1 U519 ( .A(KEYINPUT36), .B(n568), .Z(n588) );
  NOR2_X1 U520 ( .A1(n588), .A2(n460), .ZN(n461) );
  NAND2_X1 U521 ( .A1(n583), .A2(n461), .ZN(n462) );
  XNOR2_X1 U522 ( .A(KEYINPUT37), .B(n462), .ZN(n490) );
  NAND2_X1 U523 ( .A1(n463), .A2(n490), .ZN(n464) );
  XNOR2_X1 U524 ( .A(n465), .B(n464), .ZN(n475) );
  INV_X1 U525 ( .A(n491), .ZN(n551) );
  NAND2_X1 U526 ( .A1(n475), .A2(n551), .ZN(n466) );
  XNOR2_X1 U527 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U528 ( .A(G29GAT), .B(n468), .Z(G1328GAT) );
  INV_X1 U529 ( .A(n493), .ZN(n548) );
  NAND2_X1 U530 ( .A1(n475), .A2(n548), .ZN(n469) );
  XNOR2_X1 U531 ( .A(n469), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U532 ( .A(KEYINPUT40), .B(KEYINPUT100), .Z(n472) );
  NAND2_X1 U533 ( .A1(n475), .A2(n470), .ZN(n471) );
  XNOR2_X1 U534 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U535 ( .A(G43GAT), .B(n473), .Z(G1330GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n477) );
  NAND2_X1 U537 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U539 ( .A(G50GAT), .B(n478), .ZN(G1331GAT) );
  XNOR2_X1 U540 ( .A(KEYINPUT41), .B(n579), .ZN(n538) );
  XNOR2_X1 U541 ( .A(n538), .B(KEYINPUT103), .ZN(n560) );
  AND2_X1 U542 ( .A1(n576), .A2(n560), .ZN(n489) );
  NAND2_X1 U543 ( .A1(n489), .A2(n479), .ZN(n485) );
  NOR2_X1 U544 ( .A1(n491), .A2(n485), .ZN(n481) );
  XNOR2_X1 U545 ( .A(KEYINPUT42), .B(KEYINPUT104), .ZN(n480) );
  XNOR2_X1 U546 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U547 ( .A(G57GAT), .B(n482), .Z(G1332GAT) );
  NOR2_X1 U548 ( .A1(n493), .A2(n485), .ZN(n483) );
  XOR2_X1 U549 ( .A(G64GAT), .B(n483), .Z(G1333GAT) );
  NOR2_X1 U550 ( .A1(n557), .A2(n485), .ZN(n484) );
  XOR2_X1 U551 ( .A(G71GAT), .B(n484), .Z(G1334GAT) );
  NOR2_X1 U552 ( .A1(n519), .A2(n485), .ZN(n487) );
  XNOR2_X1 U553 ( .A(KEYINPUT43), .B(KEYINPUT105), .ZN(n486) );
  XNOR2_X1 U554 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U555 ( .A(G78GAT), .B(n488), .Z(G1335GAT) );
  NAND2_X1 U556 ( .A1(n490), .A2(n489), .ZN(n497) );
  NOR2_X1 U557 ( .A1(n491), .A2(n497), .ZN(n492) );
  XOR2_X1 U558 ( .A(G85GAT), .B(n492), .Z(G1336GAT) );
  NOR2_X1 U559 ( .A1(n493), .A2(n497), .ZN(n494) );
  XOR2_X1 U560 ( .A(KEYINPUT106), .B(n494), .Z(n495) );
  XNOR2_X1 U561 ( .A(G92GAT), .B(n495), .ZN(G1337GAT) );
  NOR2_X1 U562 ( .A1(n557), .A2(n497), .ZN(n496) );
  XOR2_X1 U563 ( .A(G99GAT), .B(n496), .Z(G1338GAT) );
  NOR2_X1 U564 ( .A1(n519), .A2(n497), .ZN(n499) );
  XNOR2_X1 U565 ( .A(KEYINPUT107), .B(KEYINPUT44), .ZN(n498) );
  XNOR2_X1 U566 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U567 ( .A(G106GAT), .B(n500), .ZN(G1339GAT) );
  XNOR2_X1 U568 ( .A(G113GAT), .B(KEYINPUT113), .ZN(n522) );
  NOR2_X1 U569 ( .A1(n576), .A2(n538), .ZN(n502) );
  XNOR2_X1 U570 ( .A(KEYINPUT109), .B(KEYINPUT46), .ZN(n501) );
  XNOR2_X1 U571 ( .A(n502), .B(n501), .ZN(n505) );
  INV_X1 U572 ( .A(n568), .ZN(n544) );
  XOR2_X1 U573 ( .A(n583), .B(KEYINPUT108), .Z(n564) );
  INV_X1 U574 ( .A(n564), .ZN(n503) );
  AND2_X1 U575 ( .A1(n544), .A2(n503), .ZN(n504) );
  NAND2_X1 U576 ( .A1(n505), .A2(n504), .ZN(n507) );
  XOR2_X1 U577 ( .A(KEYINPUT47), .B(KEYINPUT110), .Z(n506) );
  XNOR2_X1 U578 ( .A(n507), .B(n506), .ZN(n513) );
  OR2_X1 U579 ( .A1(n588), .A2(n583), .ZN(n508) );
  XNOR2_X1 U580 ( .A(KEYINPUT45), .B(n508), .ZN(n509) );
  NOR2_X1 U581 ( .A1(n579), .A2(n509), .ZN(n511) );
  NAND2_X1 U582 ( .A1(n511), .A2(n510), .ZN(n512) );
  NAND2_X1 U583 ( .A1(n513), .A2(n512), .ZN(n515) );
  NAND2_X1 U584 ( .A1(n547), .A2(n516), .ZN(n517) );
  XOR2_X1 U585 ( .A(KEYINPUT111), .B(n517), .Z(n534) );
  NOR2_X1 U586 ( .A1(n534), .A2(n557), .ZN(n518) );
  NAND2_X1 U587 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U588 ( .A(KEYINPUT112), .B(n520), .Z(n530) );
  AND2_X1 U589 ( .A1(n558), .A2(n530), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n522), .B(n521), .ZN(G1340GAT) );
  XOR2_X1 U591 ( .A(G120GAT), .B(KEYINPUT114), .Z(n524) );
  NAND2_X1 U592 ( .A1(n530), .A2(n560), .ZN(n523) );
  XNOR2_X1 U593 ( .A(n524), .B(n523), .ZN(n526) );
  XOR2_X1 U594 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n525) );
  XNOR2_X1 U595 ( .A(n526), .B(n525), .ZN(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n528) );
  NAND2_X1 U597 ( .A1(n564), .A2(n530), .ZN(n527) );
  XNOR2_X1 U598 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U599 ( .A(G127GAT), .B(n529), .Z(G1342GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n532) );
  NAND2_X1 U601 ( .A1(n568), .A2(n530), .ZN(n531) );
  XNOR2_X1 U602 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U603 ( .A(G134GAT), .B(n533), .Z(G1343GAT) );
  OR2_X1 U604 ( .A1(n574), .A2(n534), .ZN(n543) );
  NOR2_X1 U605 ( .A1(n576), .A2(n543), .ZN(n535) );
  XOR2_X1 U606 ( .A(G141GAT), .B(n535), .Z(G1344GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n537) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n536) );
  XNOR2_X1 U609 ( .A(n537), .B(n536), .ZN(n540) );
  NOR2_X1 U610 ( .A1(n538), .A2(n543), .ZN(n539) );
  XOR2_X1 U611 ( .A(n540), .B(n539), .Z(G1345GAT) );
  NOR2_X1 U612 ( .A1(n583), .A2(n543), .ZN(n542) );
  XNOR2_X1 U613 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n541) );
  XNOR2_X1 U614 ( .A(n542), .B(n541), .ZN(G1346GAT) );
  NOR2_X1 U615 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U616 ( .A(KEYINPUT120), .B(n545), .Z(n546) );
  XNOR2_X1 U617 ( .A(G162GAT), .B(n546), .ZN(G1347GAT) );
  NAND2_X1 U618 ( .A1(n548), .A2(n547), .ZN(n550) );
  XOR2_X1 U619 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n549) );
  XNOR2_X1 U620 ( .A(n550), .B(n549), .ZN(n552) );
  NOR2_X1 U621 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n553), .B(KEYINPUT65), .ZN(n573) );
  NOR2_X1 U623 ( .A1(n554), .A2(n573), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n555), .B(KEYINPUT55), .ZN(n556) );
  NAND2_X1 U625 ( .A1(n567), .A2(n558), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(n559), .ZN(G1348GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n562) );
  NAND2_X1 U628 ( .A1(n567), .A2(n560), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G176GAT), .ZN(G1349GAT) );
  NAND2_X1 U631 ( .A1(n567), .A2(n564), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(KEYINPUT122), .ZN(n566) );
  XNOR2_X1 U633 ( .A(G183GAT), .B(n566), .ZN(G1350GAT) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1351GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n572) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n578) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U641 ( .A(KEYINPUT123), .B(n575), .Z(n580) );
  INV_X1 U642 ( .A(n580), .ZN(n587) );
  NOR2_X1 U643 ( .A1(n576), .A2(n587), .ZN(n577) );
  XOR2_X1 U644 ( .A(n578), .B(n577), .Z(G1352GAT) );
  XOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .Z(n582) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n587), .ZN(n585) );
  XNOR2_X1 U649 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(G211GAT), .B(n586), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U653 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

