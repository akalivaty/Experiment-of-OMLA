//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n202));
  NAND2_X1  g001(.A1(G229gat), .A2(G233gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n203), .B(KEYINPUT13), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G8gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(G15gat), .B(G22gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(G1gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT89), .ZN(new_n209));
  INV_X1    g008(.A(G1gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT16), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n209), .B1(new_n207), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n207), .A2(new_n209), .A3(new_n211), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n207), .A2(new_n211), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT88), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n215), .B(new_n216), .C1(G1gat), .C2(new_n207), .ZN(new_n217));
  INV_X1    g016(.A(G22gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G15gat), .ZN(new_n219));
  INV_X1    g018(.A(G15gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G22gat), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n219), .A2(new_n221), .A3(new_n211), .A4(KEYINPUT88), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n222), .A2(G8gat), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n213), .A2(new_n214), .B1(new_n217), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT15), .ZN(new_n225));
  AND2_X1   g024(.A1(G43gat), .A2(G50gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(G43gat), .A2(G50gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n225), .B1(new_n228), .B2(KEYINPUT86), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G36gat), .ZN(new_n231));
  INV_X1    g030(.A(G29gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT84), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT84), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G29gat), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n231), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n232), .A2(new_n231), .A3(KEYINPUT14), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT14), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(G29gat), .B2(G36gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n236), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n228), .A2(KEYINPUT86), .A3(new_n225), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n230), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  OR2_X1    g042(.A1(G43gat), .A2(G50gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(G43gat), .A2(G50gat), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n225), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(new_n236), .B2(new_n240), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT85), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI211_X1 g048(.A(KEYINPUT85), .B(new_n246), .C1(new_n236), .C2(new_n240), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n224), .A2(KEYINPUT93), .A3(new_n243), .A4(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT84), .B(G29gat), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n239), .B(new_n237), .C1(new_n253), .C2(new_n231), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT85), .B1(new_n254), .B2(new_n246), .ZN(new_n255));
  INV_X1    g054(.A(new_n250), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n243), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n212), .ZN(new_n258));
  OR2_X1    g057(.A1(new_n207), .A2(G1gat), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n258), .A2(new_n259), .A3(new_n206), .A4(new_n214), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n217), .A2(new_n223), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n252), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT93), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n265), .B1(new_n257), .B2(new_n262), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n205), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT92), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n243), .B(KEYINPUT17), .C1(new_n255), .C2(new_n256), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n224), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT87), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n254), .A2(new_n229), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n249), .A2(new_n250), .B1(new_n272), .B2(new_n242), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n273), .B2(KEYINPUT17), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT17), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n257), .A2(KEYINPUT87), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n270), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n263), .A2(KEYINPUT18), .A3(new_n203), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n268), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n262), .B1(new_n273), .B2(KEYINPUT17), .ZN(new_n280));
  AOI211_X1 g079(.A(new_n271), .B(KEYINPUT17), .C1(new_n251), .C2(new_n243), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT87), .B1(new_n257), .B2(new_n275), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n263), .A2(KEYINPUT18), .A3(new_n203), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(KEYINPUT92), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n267), .B1(new_n279), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT90), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n263), .A2(new_n203), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n287), .B1(new_n277), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n288), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n283), .A2(KEYINPUT90), .A3(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n289), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n286), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G113gat), .B(G141gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(G169gat), .B(G197gat), .Z(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(KEYINPUT12), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT83), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n202), .B1(new_n294), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n302), .B1(new_n286), .B2(new_n293), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT94), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n286), .A2(new_n293), .A3(new_n300), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G1gat), .B(G29gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(KEYINPUT0), .ZN(new_n310));
  XOR2_X1   g109(.A(G57gat), .B(G85gat), .Z(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT5), .ZN(new_n313));
  XOR2_X1   g112(.A(G127gat), .B(G134gat), .Z(new_n314));
  XNOR2_X1  g113(.A(G113gat), .B(G120gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n314), .B1(KEYINPUT1), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT71), .ZN(new_n317));
  INV_X1    g116(.A(G113gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G120gat), .ZN(new_n319));
  XOR2_X1   g118(.A(KEYINPUT72), .B(G120gat), .Z(new_n320));
  OAI21_X1  g119(.A(new_n319), .B1(new_n320), .B2(new_n318), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n314), .A2(KEYINPUT1), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G155gat), .B(G162gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G141gat), .B(G148gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n327), .B1(KEYINPUT2), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n328), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n326), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT2), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT75), .B(G162gat), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n332), .B1(new_n333), .B2(G155gat), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n329), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n325), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n329), .B(KEYINPUT76), .C1(new_n334), .C2(new_n331), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n324), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G225gat), .A2(G233gat), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n313), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n337), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n324), .A2(new_n335), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT4), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n339), .A2(KEYINPUT3), .A3(new_n340), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n351), .A2(new_n324), .A3(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n348), .A2(new_n344), .A3(new_n350), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n346), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n349), .B(new_n347), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n357), .A2(new_n313), .A3(new_n344), .A4(new_n354), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n312), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n348), .A2(new_n350), .ZN(new_n360));
  INV_X1    g159(.A(new_n354), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n345), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n362), .B(KEYINPUT39), .C1(new_n345), .C2(new_n343), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT39), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n364), .B(new_n345), .C1(new_n360), .C2(new_n361), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n365), .A2(KEYINPUT81), .A3(new_n312), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT81), .B1(new_n365), .B2(new_n312), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT40), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n359), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G226gat), .A2(G233gat), .ZN(new_n371));
  XOR2_X1   g170(.A(KEYINPUT68), .B(G190gat), .Z(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT27), .B(G183gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT28), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT27), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(G183gat), .ZN(new_n377));
  INV_X1    g176(.A(G183gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(KEYINPUT69), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT69), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT27), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n378), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  OR2_X1    g181(.A1(new_n382), .A2(KEYINPUT70), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(KEYINPUT70), .ZN(new_n384));
  AOI211_X1 g183(.A(new_n372), .B(new_n377), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n375), .B1(new_n385), .B2(KEYINPUT28), .ZN(new_n386));
  INV_X1    g185(.A(G190gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n378), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(G169gat), .A2(G176gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n390), .A2(KEYINPUT26), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n391), .B1(G169gat), .B2(G176gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(KEYINPUT26), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n388), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n386), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G169gat), .ZN(new_n396));
  INV_X1    g195(.A(G176gat), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT65), .ZN(new_n398));
  OAI22_X1  g197(.A1(new_n396), .A2(new_n397), .B1(new_n398), .B2(KEYINPUT23), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n398), .A2(KEYINPUT23), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n390), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n389), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n389), .A2(KEYINPUT23), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT64), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n401), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT66), .ZN(new_n407));
  NAND3_X1  g206(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(new_n378), .B2(new_n387), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n406), .A2(new_n407), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n407), .B2(new_n406), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT25), .ZN(new_n413));
  XOR2_X1   g212(.A(KEYINPUT67), .B(KEYINPUT24), .Z(new_n414));
  OAI221_X1 g213(.A(new_n408), .B1(new_n414), .B2(new_n388), .C1(G183gat), .C2(new_n372), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n401), .A2(KEYINPUT25), .A3(new_n403), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n412), .A2(new_n413), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n395), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n371), .B1(new_n418), .B2(KEYINPUT29), .ZN(new_n419));
  XNOR2_X1  g218(.A(G197gat), .B(G204gat), .ZN(new_n420));
  INV_X1    g219(.A(G211gat), .ZN(new_n421));
  INV_X1    g220(.A(G218gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n420), .B1(KEYINPUT22), .B2(new_n423), .ZN(new_n424));
  XOR2_X1   g223(.A(G211gat), .B(G218gat), .Z(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  OR2_X1    g225(.A1(new_n426), .A2(KEYINPUT73), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(KEYINPUT73), .A3(new_n425), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n413), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n386), .A2(new_n394), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n371), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n430), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G8gat), .B(G36gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(G64gat), .B(G92gat), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n438), .B(new_n439), .Z(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n441), .B1(new_n395), .B2(new_n417), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n435), .B1(new_n442), .B2(new_n371), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n437), .B(new_n440), .C1(new_n430), .C2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT30), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n440), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n419), .A2(new_n430), .A3(new_n436), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n443), .A2(new_n430), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OR2_X1    g249(.A1(new_n443), .A2(new_n430), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n451), .A2(KEYINPUT30), .A3(new_n437), .A4(new_n440), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n446), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n363), .B(KEYINPUT40), .C1(new_n366), .C2(new_n367), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n370), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT79), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n353), .A2(new_n441), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n456), .B1(new_n429), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G228gat), .A2(G233gat), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT3), .B1(new_n426), .B2(new_n441), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n459), .B1(new_n460), .B2(new_n336), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n429), .A2(new_n457), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n462), .B1(KEYINPUT79), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n352), .B1(new_n429), .B2(KEYINPUT29), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n465), .A2(new_n341), .B1(new_n429), .B2(new_n457), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n464), .B(G22gat), .C1(new_n459), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n341), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n459), .B1(new_n468), .B2(new_n463), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n463), .A2(KEYINPUT79), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n470), .A2(new_n458), .A3(new_n461), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n218), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  XOR2_X1   g271(.A(G78gat), .B(G106gat), .Z(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT31), .B(G50gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(KEYINPUT80), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n467), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n475), .A2(KEYINPUT80), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n478), .B1(new_n467), .B2(new_n472), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n455), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n359), .A2(KEYINPUT6), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n356), .A2(new_n358), .A3(new_n312), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT6), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n444), .B(new_n483), .C1(new_n486), .C2(new_n359), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n419), .A2(new_n429), .A3(new_n436), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n488), .B(KEYINPUT37), .C1(new_n429), .C2(new_n443), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n451), .A2(new_n437), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n447), .B(new_n489), .C1(new_n490), .C2(KEYINPUT37), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT38), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT37), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n450), .B1(new_n494), .B2(new_n440), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n492), .B1(new_n490), .B2(KEYINPUT37), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n487), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  XOR2_X1   g297(.A(G15gat), .B(G43gat), .Z(new_n499));
  XNOR2_X1  g298(.A(G71gat), .B(G99gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n325), .B1(new_n395), .B2(new_n417), .ZN(new_n503));
  AND2_X1   g302(.A1(G227gat), .A2(G233gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n433), .A2(new_n324), .A3(new_n434), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT33), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n504), .B1(new_n503), .B2(new_n505), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT34), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI211_X1 g310(.A(KEYINPUT34), .B(new_n504), .C1(new_n503), .C2(new_n505), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n508), .A2(new_n511), .A3(new_n512), .ZN(new_n515));
  INV_X1    g314(.A(new_n506), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT32), .ZN(new_n517));
  OAI22_X1  g316(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n511), .A2(new_n512), .ZN(new_n519));
  INV_X1    g318(.A(new_n508), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n516), .A2(new_n517), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n522), .A3(new_n513), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n518), .A2(KEYINPUT36), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT36), .B1(new_n518), .B2(new_n523), .ZN(new_n525));
  OAI22_X1  g324(.A1(new_n482), .A2(new_n498), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT77), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n486), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n359), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n484), .A2(KEYINPUT77), .A3(new_n485), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT78), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT78), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n528), .A2(new_n529), .A3(new_n533), .A4(new_n530), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n534), .A3(new_n483), .ZN(new_n535));
  INV_X1    g334(.A(new_n453), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n481), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n526), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT35), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n483), .B1(new_n486), .B2(new_n359), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n481), .A2(new_n518), .A3(new_n523), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n521), .A2(new_n522), .A3(new_n513), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n522), .B1(new_n521), .B2(new_n513), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n535), .A2(new_n536), .A3(new_n481), .A4(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n543), .B1(new_n547), .B2(KEYINPUT35), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n308), .B1(new_n538), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n551));
  OR2_X1    g350(.A1(G71gat), .A2(G78gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(G71gat), .A2(G78gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT97), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n552), .A2(KEYINPUT97), .A3(new_n553), .ZN(new_n557));
  OR2_X1    g356(.A1(G57gat), .A2(G64gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT96), .ZN(new_n559));
  NAND2_X1  g358(.A1(G57gat), .A2(G64gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n560), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT96), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n556), .A2(new_n557), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n554), .A2(KEYINPUT95), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT95), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n552), .A2(new_n566), .A3(new_n553), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n565), .B(new_n567), .C1(new_n551), .C2(new_n562), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(KEYINPUT21), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G183gat), .B(G211gat), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n573), .B(new_n574), .Z(new_n575));
  AOI21_X1  g374(.A(new_n262), .B1(KEYINPUT21), .B2(new_n570), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(KEYINPUT100), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(KEYINPUT100), .ZN(new_n580));
  XOR2_X1   g379(.A(G127gat), .B(G155gat), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT99), .ZN(new_n582));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n583), .B(KEYINPUT98), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n582), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n579), .A2(new_n580), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n586), .B1(new_n579), .B2(new_n580), .ZN(new_n588));
  OR3_X1    g387(.A1(new_n575), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n575), .B1(new_n587), .B2(new_n588), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n592), .B(KEYINPUT101), .Z(new_n593));
  INV_X1    g392(.A(KEYINPUT41), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G134gat), .B(G162gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n599), .B(KEYINPUT104), .Z(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n274), .A2(new_n276), .ZN(new_n602));
  NAND2_X1  g401(.A1(G85gat), .A2(G92gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT7), .ZN(new_n604));
  OR2_X1    g403(.A1(G99gat), .A2(G106gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(KEYINPUT102), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(G85gat), .ZN(new_n608));
  INV_X1    g407(.A(G92gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n604), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT102), .B1(new_n605), .B2(new_n606), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n615), .B1(new_n273), .B2(KEYINPUT17), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n602), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT103), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n602), .A2(KEYINPUT103), .A3(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n615), .ZN(new_n622));
  OAI22_X1  g421(.A1(new_n622), .A2(new_n273), .B1(new_n594), .B2(new_n593), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n601), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  AOI211_X1 g424(.A(new_n600), .B(new_n623), .C1(new_n619), .C2(new_n620), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n598), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n620), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT103), .B1(new_n602), .B2(new_n616), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n624), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n600), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n621), .A2(new_n601), .A3(new_n624), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n631), .A2(new_n597), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n611), .A2(new_n612), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n611), .A2(new_n612), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n564), .B(new_n568), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n569), .A2(new_n613), .A3(new_n614), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT10), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n615), .A2(new_n570), .A3(KEYINPUT10), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n636), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n639), .A2(new_n640), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n644), .B1(new_n645), .B2(new_n636), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  OR2_X1    g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n642), .A2(new_n643), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n635), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n645), .A2(new_n636), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n652), .A2(new_n653), .A3(new_n649), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n591), .A2(new_n634), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n550), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(new_n535), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(new_n210), .ZN(G1324gat));
  NOR2_X1   g460(.A1(new_n659), .A2(new_n536), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n206), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT105), .B(KEYINPUT16), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(new_n206), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n663), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n668), .B1(new_n664), .B2(new_n667), .ZN(G1325gat));
  OR2_X1    g468(.A1(new_n524), .A2(new_n525), .ZN(new_n670));
  OAI21_X1  g469(.A(G15gat), .B1(new_n659), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n546), .A2(new_n220), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n671), .B1(new_n659), .B2(new_n672), .ZN(G1326gat));
  NOR2_X1   g472(.A1(new_n659), .A2(new_n481), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT43), .B(G22gat), .Z(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  INV_X1    g475(.A(new_n253), .ZN(new_n677));
  INV_X1    g476(.A(new_n634), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n526), .A2(new_n537), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(new_n548), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g481(.A(KEYINPUT44), .B(new_n678), .C1(new_n679), .C2(new_n548), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n591), .A2(new_n655), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n685), .A2(new_n307), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n677), .B1(new_n687), .B2(new_n535), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT45), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n685), .A2(new_n678), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT106), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n550), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n535), .A2(new_n677), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n689), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n550), .A2(KEYINPUT45), .A3(new_n691), .A4(new_n693), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n688), .A2(new_n695), .A3(new_n696), .ZN(G1328gat));
  OAI21_X1  g496(.A(G36gat), .B1(new_n687), .B2(new_n536), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n536), .A2(G36gat), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT46), .B1(new_n692), .B2(new_n700), .ZN(new_n701));
  OR3_X1    g500(.A1(new_n692), .A2(KEYINPUT46), .A3(new_n700), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n698), .A2(new_n701), .A3(new_n702), .ZN(G1329gat));
  INV_X1    g502(.A(new_n670), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n684), .A2(G43gat), .A3(new_n704), .A4(new_n686), .ZN(new_n705));
  OR2_X1    g504(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n550), .A2(new_n546), .A3(new_n691), .ZN(new_n707));
  INV_X1    g506(.A(G43gat), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n707), .A2(new_n708), .B1(KEYINPUT107), .B2(KEYINPUT47), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n705), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n706), .B1(new_n705), .B2(new_n709), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(G1330gat));
  NOR2_X1   g511(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT109), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n682), .A2(new_n480), .A3(new_n683), .A4(new_n686), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(G50gat), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n481), .A2(G50gat), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n550), .A2(new_n691), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n714), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n720), .ZN(new_n722));
  INV_X1    g521(.A(new_n714), .ZN(new_n723));
  AOI211_X1 g522(.A(new_n722), .B(new_n723), .C1(new_n716), .C2(new_n718), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n721), .A2(new_n724), .ZN(G1331gat));
  NAND4_X1  g524(.A1(new_n308), .A2(new_n591), .A3(new_n634), .A4(new_n655), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n726), .B1(new_n538), .B2(new_n549), .ZN(new_n727));
  INV_X1    g526(.A(new_n535), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n453), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n732));
  XOR2_X1   g531(.A(KEYINPUT49), .B(G64gat), .Z(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n731), .B2(new_n733), .ZN(G1333gat));
  NAND2_X1  g533(.A1(new_n727), .A2(new_n704), .ZN(new_n735));
  INV_X1    g534(.A(new_n546), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(G71gat), .ZN(new_n737));
  AOI22_X1  g536(.A1(new_n735), .A2(G71gat), .B1(new_n727), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g538(.A1(new_n727), .A2(new_n480), .ZN(new_n740));
  XOR2_X1   g539(.A(KEYINPUT110), .B(G78gat), .Z(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1335gat));
  AOI21_X1  g541(.A(new_n634), .B1(new_n538), .B2(new_n549), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n307), .A2(new_n591), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n743), .A2(KEYINPUT112), .A3(KEYINPUT51), .A4(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n678), .B(new_n744), .C1(new_n679), .C2(new_n548), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n748), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n747), .A2(KEYINPUT113), .A3(new_n748), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n750), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n755), .A2(new_n608), .A3(new_n728), .A4(new_n655), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n744), .A2(new_n655), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT111), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n684), .A2(new_n758), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n759), .A2(new_n728), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n756), .B1(new_n760), .B2(new_n608), .ZN(G1336gat));
  NAND3_X1  g560(.A1(new_n453), .A2(new_n609), .A3(new_n655), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT114), .Z(new_n763));
  AND3_X1   g562(.A1(new_n747), .A2(KEYINPUT115), .A3(new_n748), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT115), .B1(new_n747), .B2(new_n748), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n763), .B1(new_n766), .B2(new_n750), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n682), .A2(new_n453), .A3(new_n683), .A4(new_n758), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n768), .A2(G92gat), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT52), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n763), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n745), .A2(new_n749), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n753), .A2(new_n754), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT52), .B1(new_n768), .B2(G92gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n770), .A2(new_n776), .ZN(G1337gat));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n704), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G99gat), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n736), .A2(G99gat), .A3(new_n656), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n755), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(G1338gat));
  NOR3_X1   g581(.A1(new_n481), .A2(G106gat), .A3(new_n656), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n784), .B1(new_n766), .B2(new_n750), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n682), .A2(new_n480), .A3(new_n683), .A4(new_n758), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n786), .A2(G106gat), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT53), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n783), .B1(new_n772), .B2(new_n773), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT53), .B1(new_n786), .B2(G106gat), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n791), .ZN(G1339gat));
  NOR2_X1   g591(.A1(new_n657), .A2(new_n307), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n642), .A2(new_n643), .A3(new_n636), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n652), .A2(KEYINPUT54), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n649), .B1(new_n644), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n795), .A2(KEYINPUT55), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n654), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT55), .B1(new_n795), .B2(new_n797), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n627), .A2(new_n801), .A3(new_n633), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n203), .B1(new_n283), .B2(new_n263), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n264), .A2(new_n205), .A3(new_n266), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n299), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n306), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n655), .A2(new_n306), .A3(new_n805), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n307), .B2(new_n801), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n808), .B1(new_n811), .B2(new_n678), .ZN(new_n812));
  INV_X1    g611(.A(new_n591), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n793), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n480), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n815), .A2(new_n728), .A3(new_n536), .A4(new_n546), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n816), .A2(new_n318), .A3(new_n308), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n814), .A2(new_n535), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n542), .A2(new_n453), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(new_n307), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n817), .B1(new_n318), .B2(new_n820), .ZN(G1340gat));
  OAI21_X1  g620(.A(G120gat), .B1(new_n816), .B2(new_n656), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n818), .A2(new_n819), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n656), .A2(new_n320), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(G1341gat));
  OAI21_X1  g624(.A(G127gat), .B1(new_n816), .B2(new_n813), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n813), .A2(G127gat), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n826), .B1(new_n823), .B2(new_n827), .ZN(G1342gat));
  OR3_X1    g627(.A1(new_n823), .A2(G134gat), .A3(new_n634), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n829), .A2(KEYINPUT56), .ZN(new_n830));
  OAI21_X1  g629(.A(G134gat), .B1(new_n816), .B2(new_n634), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(KEYINPUT56), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(G1343gat));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n658), .A2(new_n308), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n306), .B1(new_n304), .B2(KEYINPUT94), .ZN(new_n836));
  AOI211_X1 g635(.A(new_n202), .B(new_n302), .C1(new_n286), .C2(new_n293), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n801), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n809), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n807), .B1(new_n839), .B2(new_n634), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n835), .B1(new_n840), .B2(new_n591), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n480), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n842), .A2(KEYINPUT57), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n795), .A2(new_n797), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT55), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n795), .A2(KEYINPUT116), .A3(new_n797), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n799), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n848), .B1(new_n836), .B2(new_n837), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n809), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n807), .B1(new_n850), .B2(new_n634), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n835), .B1(new_n851), .B2(new_n591), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT57), .B1(new_n853), .B2(new_n481), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n670), .A2(new_n728), .A3(new_n536), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n843), .A2(new_n854), .A3(new_n307), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(G141gat), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n818), .A2(new_n480), .A3(new_n670), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n858), .A2(KEYINPUT118), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(KEYINPUT118), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n536), .A3(new_n860), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n308), .A2(G141gat), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n834), .B(new_n857), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n857), .A2(KEYINPUT117), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n865), .B1(new_n856), .B2(G141gat), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n858), .A2(new_n453), .A3(new_n862), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n864), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n863), .B1(new_n868), .B2(new_n834), .ZN(G1344gat));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n843), .A2(new_n855), .A3(new_n854), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n870), .B(G148gat), .C1(new_n871), .C2(new_n656), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n873));
  INV_X1    g672(.A(G148gat), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n852), .A2(KEYINPUT119), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n876), .B(new_n835), .C1(new_n851), .C2(new_n591), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n481), .A2(KEYINPUT57), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT57), .B1(new_n814), .B2(new_n481), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n879), .A2(new_n655), .A3(new_n855), .A4(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n874), .B1(new_n881), .B2(KEYINPUT120), .ZN(new_n882));
  INV_X1    g681(.A(new_n878), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n883), .B1(new_n852), .B2(KEYINPUT119), .ZN(new_n884));
  AOI22_X1  g683(.A1(new_n884), .A2(new_n877), .B1(new_n842), .B2(KEYINPUT57), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n885), .A2(new_n886), .A3(new_n655), .A4(new_n855), .ZN(new_n887));
  AOI211_X1 g686(.A(new_n873), .B(new_n870), .C1(new_n882), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n881), .A2(KEYINPUT120), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n887), .A3(G148gat), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT121), .B1(new_n890), .B2(KEYINPUT59), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n872), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  OR3_X1    g691(.A1(new_n861), .A2(G148gat), .A3(new_n656), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1345gat));
  OAI21_X1  g693(.A(G155gat), .B1(new_n871), .B2(new_n813), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n813), .A2(G155gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n861), .B2(new_n896), .ZN(G1346gat));
  OAI21_X1  g696(.A(new_n333), .B1(new_n871), .B2(new_n634), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n634), .A2(new_n333), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n898), .B1(new_n861), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT122), .ZN(G1347gat));
  NOR2_X1   g701(.A1(new_n814), .A2(new_n728), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n903), .A2(new_n453), .A3(new_n481), .A4(new_n546), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(G169gat), .B1(new_n905), .B2(new_n307), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n728), .A2(new_n536), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n815), .A2(new_n546), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT123), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n308), .A2(new_n396), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n906), .B1(new_n909), .B2(new_n910), .ZN(G1348gat));
  NAND3_X1  g710(.A1(new_n905), .A2(new_n397), .A3(new_n655), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n909), .A2(new_n655), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(new_n397), .ZN(G1349gat));
  AOI21_X1  g713(.A(new_n378), .B1(new_n909), .B2(new_n591), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n905), .A2(new_n374), .A3(new_n591), .ZN(new_n916));
  OR3_X1    g715(.A1(new_n915), .A2(KEYINPUT60), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT60), .B1(new_n915), .B2(new_n916), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1350gat));
  AOI21_X1  g718(.A(new_n387), .B1(new_n909), .B2(new_n678), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT124), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n921), .A2(KEYINPUT124), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n905), .A2(new_n373), .A3(new_n678), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n924), .B(new_n925), .C1(new_n920), .C2(new_n922), .ZN(G1351gat));
  AND2_X1   g725(.A1(new_n907), .A2(new_n670), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n885), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(G197gat), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n928), .A2(new_n929), .A3(new_n308), .ZN(new_n930));
  AND4_X1   g729(.A1(new_n453), .A2(new_n903), .A3(new_n480), .A4(new_n670), .ZN(new_n931));
  AOI21_X1  g730(.A(G197gat), .B1(new_n931), .B2(new_n307), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n930), .A2(new_n932), .ZN(G1352gat));
  INV_X1    g732(.A(G204gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n931), .A2(new_n934), .A3(new_n655), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT62), .Z(new_n936));
  AND3_X1   g735(.A1(new_n885), .A2(new_n655), .A3(new_n927), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n934), .B2(new_n937), .ZN(G1353gat));
  NAND3_X1  g737(.A1(new_n885), .A2(new_n591), .A3(new_n927), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT63), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n421), .B1(KEYINPUT125), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(new_n943), .A3(KEYINPUT63), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n939), .B(new_n941), .C1(KEYINPUT125), .C2(new_n940), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n931), .A2(new_n421), .A3(new_n591), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(G1354gat));
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n634), .B1(new_n928), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n949), .B1(new_n948), .B2(new_n928), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G218gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n931), .A2(new_n422), .A3(new_n678), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1355gat));
endmodule


