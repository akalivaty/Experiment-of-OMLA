

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582;

  XOR2_X1 U320 ( .A(n358), .B(n357), .Z(n465) );
  XNOR2_X1 U321 ( .A(n412), .B(KEYINPUT31), .ZN(n413) );
  XNOR2_X1 U322 ( .A(n414), .B(n413), .ZN(n417) );
  INV_X1 U323 ( .A(KEYINPUT95), .ZN(n388) );
  XNOR2_X1 U324 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U325 ( .A(KEYINPUT37), .B(KEYINPUT102), .ZN(n408) );
  XNOR2_X1 U326 ( .A(n425), .B(n424), .ZN(n571) );
  XNOR2_X1 U327 ( .A(n409), .B(n408), .ZN(n505) );
  NOR2_X1 U328 ( .A1(n382), .A2(n467), .ZN(n559) );
  XNOR2_X1 U329 ( .A(n445), .B(KEYINPUT38), .ZN(n492) );
  XNOR2_X1 U330 ( .A(G183GAT), .B(KEYINPUT120), .ZN(n468) );
  XNOR2_X1 U331 ( .A(n446), .B(G29GAT), .ZN(n447) );
  XNOR2_X1 U332 ( .A(n469), .B(n468), .ZN(G1350GAT) );
  XNOR2_X1 U333 ( .A(n448), .B(n447), .ZN(G1328GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT2), .B(G162GAT), .Z(n289) );
  XNOR2_X1 U335 ( .A(G155GAT), .B(G141GAT), .ZN(n288) );
  XNOR2_X1 U336 ( .A(n289), .B(n288), .ZN(n290) );
  XNOR2_X1 U337 ( .A(KEYINPUT3), .B(n290), .ZN(n350) );
  XOR2_X1 U338 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n292) );
  XNOR2_X1 U339 ( .A(KEYINPUT6), .B(KEYINPUT86), .ZN(n291) );
  XNOR2_X1 U340 ( .A(n292), .B(n291), .ZN(n303) );
  XOR2_X1 U341 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n294) );
  XNOR2_X1 U342 ( .A(G85GAT), .B(KEYINPUT4), .ZN(n293) );
  XNOR2_X1 U343 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U344 ( .A(G113GAT), .B(G1GAT), .Z(n431) );
  XOR2_X1 U345 ( .A(n295), .B(n431), .Z(n301) );
  XOR2_X1 U346 ( .A(G29GAT), .B(G134GAT), .Z(n318) );
  XNOR2_X1 U347 ( .A(G148GAT), .B(G120GAT), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n296), .B(G57GAT), .ZN(n415) );
  XOR2_X1 U349 ( .A(n318), .B(n415), .Z(n298) );
  NAND2_X1 U350 ( .A1(G225GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U352 ( .A(KEYINPUT0), .B(G127GAT), .Z(n332) );
  XNOR2_X1 U353 ( .A(n299), .B(n332), .ZN(n300) );
  XNOR2_X1 U354 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U355 ( .A(n303), .B(n302), .Z(n304) );
  XNOR2_X1 U356 ( .A(n350), .B(n304), .ZN(n379) );
  XNOR2_X1 U357 ( .A(KEYINPUT87), .B(n379), .ZN(n476) );
  INV_X1 U358 ( .A(n476), .ZN(n506) );
  XOR2_X1 U359 ( .A(KEYINPUT11), .B(G92GAT), .Z(n306) );
  XNOR2_X1 U360 ( .A(G162GAT), .B(KEYINPUT74), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n322) );
  XOR2_X1 U362 ( .A(G106GAT), .B(G218GAT), .Z(n308) );
  XOR2_X1 U363 ( .A(G190GAT), .B(G36GAT), .Z(n370) );
  XOR2_X1 U364 ( .A(G85GAT), .B(G99GAT), .Z(n410) );
  XNOR2_X1 U365 ( .A(n370), .B(n410), .ZN(n307) );
  XNOR2_X1 U366 ( .A(n308), .B(n307), .ZN(n314) );
  XOR2_X1 U367 ( .A(G43GAT), .B(G50GAT), .Z(n310) );
  XNOR2_X1 U368 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n309) );
  XNOR2_X1 U369 ( .A(n310), .B(n309), .ZN(n440) );
  XOR2_X1 U370 ( .A(KEYINPUT10), .B(n440), .Z(n312) );
  NAND2_X1 U371 ( .A1(G232GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U372 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U373 ( .A(n314), .B(n313), .Z(n320) );
  XOR2_X1 U374 ( .A(KEYINPUT65), .B(KEYINPUT73), .Z(n316) );
  XNOR2_X1 U375 ( .A(KEYINPUT9), .B(KEYINPUT64), .ZN(n315) );
  XNOR2_X1 U376 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U377 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U379 ( .A(n322), .B(n321), .ZN(n545) );
  XNOR2_X1 U380 ( .A(KEYINPUT36), .B(n545), .ZN(n579) );
  XOR2_X1 U381 ( .A(G176GAT), .B(G15GAT), .Z(n324) );
  XNOR2_X1 U382 ( .A(G183GAT), .B(G71GAT), .ZN(n323) );
  XNOR2_X1 U383 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U384 ( .A(KEYINPUT20), .B(KEYINPUT79), .Z(n326) );
  XNOR2_X1 U385 ( .A(KEYINPUT78), .B(KEYINPUT80), .ZN(n325) );
  XNOR2_X1 U386 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U387 ( .A(n328), .B(n327), .ZN(n341) );
  XOR2_X1 U388 ( .A(G99GAT), .B(G190GAT), .Z(n330) );
  XNOR2_X1 U389 ( .A(G134GAT), .B(G43GAT), .ZN(n329) );
  XNOR2_X1 U390 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U391 ( .A(n332), .B(n331), .Z(n334) );
  NAND2_X1 U392 ( .A1(G227GAT), .A2(G233GAT), .ZN(n333) );
  XOR2_X1 U393 ( .A(n334), .B(n333), .Z(n337) );
  XOR2_X1 U394 ( .A(G169GAT), .B(KEYINPUT19), .Z(n336) );
  XNOR2_X1 U395 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n336), .B(n335), .ZN(n365) );
  XNOR2_X1 U397 ( .A(n337), .B(n365), .ZN(n339) );
  XNOR2_X1 U398 ( .A(G120GAT), .B(G113GAT), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U400 ( .A(n341), .B(n340), .ZN(n382) );
  XOR2_X1 U401 ( .A(KEYINPUT23), .B(KEYINPUT81), .Z(n343) );
  XNOR2_X1 U402 ( .A(G22GAT), .B(G204GAT), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U404 ( .A(G106GAT), .B(G78GAT), .Z(n420) );
  XOR2_X1 U405 ( .A(n344), .B(n420), .Z(n346) );
  XNOR2_X1 U406 ( .A(G148GAT), .B(G50GAT), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n358) );
  XOR2_X1 U408 ( .A(KEYINPUT82), .B(KEYINPUT22), .Z(n348) );
  NAND2_X1 U409 ( .A1(G228GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U411 ( .A(n349), .B(KEYINPUT24), .Z(n356) );
  INV_X1 U412 ( .A(n350), .ZN(n354) );
  XOR2_X1 U413 ( .A(KEYINPUT83), .B(G197GAT), .Z(n352) );
  XNOR2_X1 U414 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n351) );
  XNOR2_X1 U415 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U416 ( .A(G211GAT), .B(n353), .Z(n369) );
  XNOR2_X1 U417 ( .A(n354), .B(n369), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n357) );
  NAND2_X1 U419 ( .A1(n382), .A2(n465), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n359), .B(KEYINPUT26), .ZN(n565) );
  XOR2_X1 U421 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n361) );
  NAND2_X1 U422 ( .A1(G226GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U424 ( .A(n362), .B(KEYINPUT90), .Z(n367) );
  XOR2_X1 U425 ( .A(G176GAT), .B(G204GAT), .Z(n364) );
  XNOR2_X1 U426 ( .A(G92GAT), .B(G64GAT), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n411) );
  XNOR2_X1 U428 ( .A(n365), .B(n411), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U430 ( .A(n369), .B(n368), .Z(n372) );
  XOR2_X1 U431 ( .A(G183GAT), .B(G8GAT), .Z(n394) );
  XNOR2_X1 U432 ( .A(n370), .B(n394), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n372), .B(n371), .ZN(n480) );
  XOR2_X1 U434 ( .A(n480), .B(KEYINPUT91), .Z(n373) );
  XNOR2_X1 U435 ( .A(KEYINPUT27), .B(n373), .ZN(n383) );
  NOR2_X1 U436 ( .A1(n565), .A2(n383), .ZN(n374) );
  XNOR2_X1 U437 ( .A(KEYINPUT93), .B(n374), .ZN(n378) );
  NOR2_X1 U438 ( .A1(n382), .A2(n480), .ZN(n375) );
  NOR2_X1 U439 ( .A1(n465), .A2(n375), .ZN(n376) );
  XNOR2_X1 U440 ( .A(KEYINPUT25), .B(n376), .ZN(n377) );
  AND2_X1 U441 ( .A1(n378), .A2(n377), .ZN(n380) );
  NOR2_X1 U442 ( .A1(n380), .A2(n379), .ZN(n381) );
  XNOR2_X1 U443 ( .A(n381), .B(KEYINPUT94), .ZN(n387) );
  INV_X1 U444 ( .A(n382), .ZN(n520) );
  NOR2_X1 U445 ( .A1(n476), .A2(n383), .ZN(n517) );
  XNOR2_X1 U446 ( .A(KEYINPUT28), .B(n465), .ZN(n519) );
  INV_X1 U447 ( .A(n519), .ZN(n486) );
  NAND2_X1 U448 ( .A1(n517), .A2(n486), .ZN(n384) );
  NOR2_X1 U449 ( .A1(n520), .A2(n384), .ZN(n385) );
  XNOR2_X1 U450 ( .A(KEYINPUT92), .B(n385), .ZN(n386) );
  NOR2_X1 U451 ( .A1(n387), .A2(n386), .ZN(n389) );
  XNOR2_X1 U452 ( .A(n389), .B(n388), .ZN(n473) );
  XOR2_X1 U453 ( .A(G211GAT), .B(G78GAT), .Z(n391) );
  XNOR2_X1 U454 ( .A(G155GAT), .B(G127GAT), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n391), .B(n390), .ZN(n405) );
  XOR2_X1 U456 ( .A(G22GAT), .B(G15GAT), .Z(n430) );
  XOR2_X1 U457 ( .A(G71GAT), .B(KEYINPUT13), .Z(n421) );
  XOR2_X1 U458 ( .A(n430), .B(n421), .Z(n393) );
  NAND2_X1 U459 ( .A1(G231GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n393), .B(n392), .ZN(n395) );
  XOR2_X1 U461 ( .A(n395), .B(n394), .Z(n403) );
  XOR2_X1 U462 ( .A(KEYINPUT12), .B(G64GAT), .Z(n397) );
  XNOR2_X1 U463 ( .A(G57GAT), .B(G1GAT), .ZN(n396) );
  XNOR2_X1 U464 ( .A(n397), .B(n396), .ZN(n401) );
  XOR2_X1 U465 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n399) );
  XNOR2_X1 U466 ( .A(KEYINPUT76), .B(KEYINPUT75), .ZN(n398) );
  XNOR2_X1 U467 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U468 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U469 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U470 ( .A(n405), .B(n404), .ZN(n576) );
  NOR2_X1 U471 ( .A1(n473), .A2(n576), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n406), .B(KEYINPUT101), .ZN(n407) );
  NOR2_X1 U473 ( .A1(n579), .A2(n407), .ZN(n409) );
  XOR2_X1 U474 ( .A(n411), .B(n410), .Z(n414) );
  NAND2_X1 U475 ( .A1(G230GAT), .A2(G233GAT), .ZN(n412) );
  XOR2_X1 U476 ( .A(n415), .B(KEYINPUT71), .Z(n416) );
  XNOR2_X1 U477 ( .A(n417), .B(n416), .ZN(n425) );
  XOR2_X1 U478 ( .A(KEYINPUT72), .B(KEYINPUT70), .Z(n419) );
  XNOR2_X1 U479 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n418) );
  XOR2_X1 U480 ( .A(n419), .B(n418), .Z(n423) );
  XNOR2_X1 U481 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U482 ( .A(G169GAT), .B(G197GAT), .Z(n427) );
  XNOR2_X1 U483 ( .A(G141GAT), .B(G8GAT), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n444) );
  XOR2_X1 U485 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n429) );
  XNOR2_X1 U486 ( .A(KEYINPUT69), .B(KEYINPUT67), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n435) );
  XOR2_X1 U488 ( .A(n430), .B(G36GAT), .Z(n433) );
  XNOR2_X1 U489 ( .A(G29GAT), .B(n431), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U491 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U492 ( .A1(G229GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n439) );
  INV_X1 U494 ( .A(KEYINPUT29), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n440), .B(KEYINPUT68), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X2 U498 ( .A(n444), .B(n443), .Z(n566) );
  NAND2_X1 U499 ( .A1(n571), .A2(n566), .ZN(n474) );
  NOR2_X1 U500 ( .A1(n505), .A2(n474), .ZN(n445) );
  NAND2_X1 U501 ( .A1(n506), .A2(n492), .ZN(n448) );
  XOR2_X1 U502 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n446) );
  INV_X1 U503 ( .A(n480), .ZN(n509) );
  XNOR2_X1 U504 ( .A(KEYINPUT45), .B(KEYINPUT108), .ZN(n450) );
  INV_X1 U505 ( .A(n576), .ZN(n531) );
  NOR2_X1 U506 ( .A1(n579), .A2(n531), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n450), .B(n449), .ZN(n451) );
  NAND2_X1 U508 ( .A1(n571), .A2(n451), .ZN(n452) );
  NOR2_X1 U509 ( .A1(n566), .A2(n452), .ZN(n453) );
  XOR2_X1 U510 ( .A(KEYINPUT109), .B(n453), .Z(n461) );
  INV_X1 U511 ( .A(KEYINPUT41), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n571), .B(n454), .ZN(n525) );
  INV_X1 U513 ( .A(n525), .ZN(n553) );
  NAND2_X1 U514 ( .A1(n553), .A2(n566), .ZN(n456) );
  XOR2_X1 U515 ( .A(KEYINPUT46), .B(KEYINPUT107), .Z(n455) );
  XNOR2_X1 U516 ( .A(n456), .B(n455), .ZN(n457) );
  NAND2_X1 U517 ( .A1(n457), .A2(n545), .ZN(n458) );
  NOR2_X1 U518 ( .A1(n576), .A2(n458), .ZN(n459) );
  XOR2_X1 U519 ( .A(KEYINPUT47), .B(n459), .Z(n460) );
  NOR2_X1 U520 ( .A1(n461), .A2(n460), .ZN(n462) );
  XOR2_X1 U521 ( .A(KEYINPUT48), .B(n462), .Z(n516) );
  AND2_X1 U522 ( .A1(n509), .A2(n516), .ZN(n463) );
  XNOR2_X1 U523 ( .A(n463), .B(KEYINPUT54), .ZN(n464) );
  NAND2_X1 U524 ( .A1(n464), .A2(n476), .ZN(n564) );
  NOR2_X1 U525 ( .A1(n465), .A2(n564), .ZN(n466) );
  XNOR2_X1 U526 ( .A(n466), .B(KEYINPUT55), .ZN(n467) );
  NAND2_X1 U527 ( .A1(n576), .A2(n559), .ZN(n469) );
  XOR2_X1 U528 ( .A(KEYINPUT77), .B(KEYINPUT16), .Z(n471) );
  NAND2_X1 U529 ( .A1(n576), .A2(n545), .ZN(n470) );
  XNOR2_X1 U530 ( .A(n471), .B(n470), .ZN(n472) );
  OR2_X1 U531 ( .A1(n473), .A2(n472), .ZN(n495) );
  NOR2_X1 U532 ( .A1(n474), .A2(n495), .ZN(n475) );
  XOR2_X1 U533 ( .A(KEYINPUT96), .B(n475), .Z(n485) );
  NOR2_X1 U534 ( .A1(n485), .A2(n476), .ZN(n478) );
  XNOR2_X1 U535 ( .A(KEYINPUT34), .B(KEYINPUT97), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U537 ( .A(G1GAT), .B(n479), .ZN(G1324GAT) );
  NOR2_X1 U538 ( .A1(n480), .A2(n485), .ZN(n481) );
  XOR2_X1 U539 ( .A(G8GAT), .B(n481), .Z(G1325GAT) );
  XNOR2_X1 U540 ( .A(KEYINPUT98), .B(KEYINPUT35), .ZN(n483) );
  NOR2_X1 U541 ( .A1(n382), .A2(n485), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U543 ( .A(G15GAT), .B(n484), .ZN(G1326GAT) );
  XNOR2_X1 U544 ( .A(G22GAT), .B(KEYINPUT99), .ZN(n488) );
  NOR2_X1 U545 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(G1327GAT) );
  NAND2_X1 U547 ( .A1(n509), .A2(n492), .ZN(n489) );
  XNOR2_X1 U548 ( .A(G36GAT), .B(n489), .ZN(G1329GAT) );
  NAND2_X1 U549 ( .A1(n492), .A2(n520), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n490), .B(KEYINPUT40), .ZN(n491) );
  XNOR2_X1 U551 ( .A(G43GAT), .B(n491), .ZN(G1330GAT) );
  XOR2_X1 U552 ( .A(G50GAT), .B(KEYINPUT103), .Z(n494) );
  NAND2_X1 U553 ( .A1(n492), .A2(n519), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(G1331GAT) );
  XNOR2_X1 U555 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n497) );
  INV_X1 U556 ( .A(n566), .ZN(n522) );
  NAND2_X1 U557 ( .A1(n522), .A2(n553), .ZN(n504) );
  NOR2_X1 U558 ( .A1(n504), .A2(n495), .ZN(n501) );
  NAND2_X1 U559 ( .A1(n506), .A2(n501), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n497), .B(n496), .ZN(G1332GAT) );
  NAND2_X1 U561 ( .A1(n509), .A2(n501), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n498), .B(KEYINPUT104), .ZN(n499) );
  XNOR2_X1 U563 ( .A(G64GAT), .B(n499), .ZN(G1333GAT) );
  NAND2_X1 U564 ( .A1(n520), .A2(n501), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n500), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U566 ( .A(G78GAT), .B(KEYINPUT43), .Z(n503) );
  NAND2_X1 U567 ( .A1(n501), .A2(n519), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(G1335GAT) );
  XOR2_X1 U569 ( .A(G85GAT), .B(KEYINPUT105), .Z(n508) );
  NOR2_X1 U570 ( .A1(n505), .A2(n504), .ZN(n512) );
  NAND2_X1 U571 ( .A1(n512), .A2(n506), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(G1336GAT) );
  NAND2_X1 U573 ( .A1(n509), .A2(n512), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n510), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U575 ( .A1(n520), .A2(n512), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n511), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT44), .B(KEYINPUT106), .Z(n514) );
  NAND2_X1 U578 ( .A1(n512), .A2(n519), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U580 ( .A(G106GAT), .B(n515), .Z(G1339GAT) );
  NAND2_X1 U581 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U582 ( .A(KEYINPUT110), .B(n518), .ZN(n537) );
  NOR2_X1 U583 ( .A1(n537), .A2(n519), .ZN(n521) );
  NAND2_X1 U584 ( .A1(n521), .A2(n520), .ZN(n534) );
  NOR2_X1 U585 ( .A1(n522), .A2(n534), .ZN(n524) );
  XNOR2_X1 U586 ( .A(G113GAT), .B(KEYINPUT111), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n524), .B(n523), .ZN(G1340GAT) );
  NOR2_X1 U588 ( .A1(n525), .A2(n534), .ZN(n527) );
  XNOR2_X1 U589 ( .A(KEYINPUT49), .B(KEYINPUT112), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G120GAT), .B(n528), .ZN(G1341GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n530) );
  XNOR2_X1 U593 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(n533) );
  NOR2_X1 U595 ( .A1(n531), .A2(n534), .ZN(n532) );
  XOR2_X1 U596 ( .A(n533), .B(n532), .Z(G1342GAT) );
  NOR2_X1 U597 ( .A1(n545), .A2(n534), .ZN(n536) );
  XNOR2_X1 U598 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n536), .B(n535), .ZN(G1343GAT) );
  XOR2_X1 U600 ( .A(G141GAT), .B(KEYINPUT115), .Z(n539) );
  NOR2_X1 U601 ( .A1(n565), .A2(n537), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n546), .A2(n566), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(G1344GAT) );
  XNOR2_X1 U604 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n543) );
  XOR2_X1 U605 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n541) );
  NAND2_X1 U606 ( .A1(n546), .A2(n553), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(G1345GAT) );
  NAND2_X1 U609 ( .A1(n576), .A2(n546), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n544), .B(G155GAT), .ZN(G1346GAT) );
  INV_X1 U611 ( .A(n545), .ZN(n558) );
  NAND2_X1 U612 ( .A1(n546), .A2(n558), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n547), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U614 ( .A(G169GAT), .B(KEYINPUT117), .Z(n549) );
  NAND2_X1 U615 ( .A1(n559), .A2(n566), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1348GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT57), .B(KEYINPUT119), .Z(n551) );
  XNOR2_X1 U618 ( .A(G176GAT), .B(KEYINPUT118), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U620 ( .A(KEYINPUT56), .B(n552), .Z(n555) );
  NAND2_X1 U621 ( .A1(n559), .A2(n553), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1349GAT) );
  XNOR2_X1 U623 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(KEYINPUT121), .ZN(n557) );
  XOR2_X1 U625 ( .A(KEYINPUT122), .B(n557), .Z(n561) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1351GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT125), .B(KEYINPUT124), .Z(n563) );
  XNOR2_X1 U629 ( .A(KEYINPUT59), .B(KEYINPUT60), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n570) );
  XOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT123), .Z(n568) );
  NOR2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n575) );
  NAND2_X1 U633 ( .A1(n575), .A2(n566), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U635 ( .A(n570), .B(n569), .Z(G1352GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n573) );
  INV_X1 U637 ( .A(n575), .ZN(n578) );
  OR2_X1 U638 ( .A1(n578), .A2(n571), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(n574), .ZN(G1353GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

