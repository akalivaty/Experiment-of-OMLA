

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U553 ( .A1(n695), .A2(n770), .ZN(n739) );
  XNOR2_X2 U554 ( .A(n782), .B(n693), .ZN(n697) );
  AND2_X1 U555 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U556 ( .A1(n701), .A2(n700), .ZN(n718) );
  BUF_X1 U557 ( .A(n617), .Z(n896) );
  INV_X1 U558 ( .A(G2104), .ZN(n546) );
  INV_X1 U559 ( .A(KEYINPUT97), .ZN(n763) );
  NOR2_X1 U560 ( .A1(n762), .A2(KEYINPUT33), .ZN(n764) );
  XNOR2_X1 U561 ( .A(n547), .B(KEYINPUT65), .ZN(n617) );
  NOR2_X1 U562 ( .A1(G2105), .A2(n546), .ZN(n572) );
  INV_X1 U563 ( .A(G301), .ZN(G171) );
  NOR2_X2 U564 ( .A1(n653), .A2(G651), .ZN(n592) );
  OR2_X1 U565 ( .A1(n810), .A2(n523), .ZN(n520) );
  XOR2_X1 U566 ( .A(KEYINPUT32), .B(KEYINPUT96), .Z(n521) );
  NOR2_X2 U567 ( .A1(n579), .A2(n578), .ZN(G160) );
  XOR2_X1 U568 ( .A(KEYINPUT68), .B(n537), .Z(n522) );
  AND2_X1 U569 ( .A1(n826), .A2(n919), .ZN(n523) );
  INV_X1 U570 ( .A(n995), .ZN(n758) );
  NOR2_X1 U571 ( .A1(n778), .A2(n758), .ZN(n759) );
  XNOR2_X1 U572 ( .A(n764), .B(n763), .ZN(n765) );
  XNOR2_X1 U573 ( .A(KEYINPUT12), .B(KEYINPUT72), .ZN(n583) );
  NOR2_X1 U574 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U575 ( .A(n584), .B(n583), .ZN(n586) );
  NOR2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n543) );
  NOR2_X1 U577 ( .A1(G651), .A2(G543), .ZN(n656) );
  NOR2_X2 U578 ( .A1(n653), .A2(n525), .ZN(n657) );
  XNOR2_X1 U579 ( .A(n542), .B(KEYINPUT69), .ZN(G301) );
  XOR2_X1 U580 ( .A(KEYINPUT71), .B(n533), .Z(G299) );
  XOR2_X1 U581 ( .A(G543), .B(KEYINPUT0), .Z(n653) );
  NAND2_X1 U582 ( .A1(n592), .A2(G53), .ZN(n532) );
  INV_X1 U583 ( .A(G651), .ZN(n525) );
  NOR2_X1 U584 ( .A1(G543), .A2(n525), .ZN(n524) );
  XOR2_X2 U585 ( .A(KEYINPUT1), .B(n524), .Z(n660) );
  NAND2_X1 U586 ( .A1(G65), .A2(n660), .ZN(n527) );
  NAND2_X1 U587 ( .A1(G78), .A2(n657), .ZN(n526) );
  NAND2_X1 U588 ( .A1(n527), .A2(n526), .ZN(n530) );
  NAND2_X1 U589 ( .A1(n656), .A2(G91), .ZN(n528) );
  XOR2_X1 U590 ( .A(KEYINPUT70), .B(n528), .Z(n529) );
  NOR2_X1 U591 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U592 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U593 ( .A1(G64), .A2(n660), .ZN(n535) );
  NAND2_X1 U594 ( .A1(G52), .A2(n592), .ZN(n534) );
  NAND2_X1 U595 ( .A1(n535), .A2(n534), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n656), .A2(G90), .ZN(n536) );
  XNOR2_X1 U597 ( .A(KEYINPUT67), .B(n536), .ZN(n538) );
  NAND2_X1 U598 ( .A1(n657), .A2(G77), .ZN(n537) );
  NOR2_X1 U599 ( .A1(n538), .A2(n522), .ZN(n539) );
  XNOR2_X1 U600 ( .A(n539), .B(KEYINPUT9), .ZN(n540) );
  NOR2_X1 U601 ( .A1(n541), .A2(n540), .ZN(n542) );
  BUF_X1 U602 ( .A(n572), .Z(n892) );
  NAND2_X1 U603 ( .A1(G102), .A2(n892), .ZN(n545) );
  XOR2_X1 U604 ( .A(KEYINPUT17), .B(n543), .Z(n619) );
  NAND2_X1 U605 ( .A1(G138), .A2(n619), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n551) );
  AND2_X1 U607 ( .A1(G2104), .A2(G2105), .ZN(n898) );
  NAND2_X1 U608 ( .A1(G114), .A2(n898), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n546), .A2(G2105), .ZN(n547) );
  NAND2_X1 U610 ( .A1(G126), .A2(n617), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U612 ( .A1(n551), .A2(n550), .ZN(G164) );
  XOR2_X1 U613 ( .A(G2443), .B(G2446), .Z(n553) );
  XNOR2_X1 U614 ( .A(G2427), .B(G2451), .ZN(n552) );
  XNOR2_X1 U615 ( .A(n553), .B(n552), .ZN(n559) );
  XOR2_X1 U616 ( .A(G2430), .B(G2454), .Z(n555) );
  XNOR2_X1 U617 ( .A(G1341), .B(G1348), .ZN(n554) );
  XNOR2_X1 U618 ( .A(n555), .B(n554), .ZN(n557) );
  XOR2_X1 U619 ( .A(G2435), .B(G2438), .Z(n556) );
  XNOR2_X1 U620 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U621 ( .A(n559), .B(n558), .Z(n560) );
  AND2_X1 U622 ( .A1(G14), .A2(n560), .ZN(G401) );
  AND2_X1 U623 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U624 ( .A(G57), .ZN(G237) );
  NAND2_X1 U625 ( .A1(n656), .A2(G89), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(KEYINPUT4), .ZN(n563) );
  NAND2_X1 U627 ( .A1(G76), .A2(n657), .ZN(n562) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(KEYINPUT5), .B(n564), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G63), .A2(n660), .ZN(n566) );
  NAND2_X1 U631 ( .A1(G51), .A2(n592), .ZN(n565) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n568) );
  XOR2_X1 U633 ( .A(KEYINPUT6), .B(KEYINPUT76), .Z(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(KEYINPUT7), .B(n571), .ZN(G168) );
  XOR2_X1 U637 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U638 ( .A1(n898), .A2(G113), .ZN(n575) );
  NAND2_X1 U639 ( .A1(G101), .A2(n572), .ZN(n573) );
  XOR2_X1 U640 ( .A(KEYINPUT23), .B(n573), .Z(n574) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U642 ( .A1(G137), .A2(n619), .ZN(n577) );
  NAND2_X1 U643 ( .A1(G125), .A2(n617), .ZN(n576) );
  NAND2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U645 ( .A1(G7), .A2(G661), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n580), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U647 ( .A(G223), .ZN(n831) );
  NAND2_X1 U648 ( .A1(n831), .A2(G567), .ZN(n581) );
  XOR2_X1 U649 ( .A(KEYINPUT11), .B(n581), .Z(G234) );
  NAND2_X1 U650 ( .A1(G56), .A2(n660), .ZN(n582) );
  XOR2_X1 U651 ( .A(KEYINPUT14), .B(n582), .Z(n589) );
  NAND2_X1 U652 ( .A1(G81), .A2(n656), .ZN(n584) );
  NAND2_X1 U653 ( .A1(G68), .A2(n657), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U655 ( .A(KEYINPUT13), .B(n587), .Z(n588) );
  NOR2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U657 ( .A1(n592), .A2(G43), .ZN(n590) );
  NAND2_X1 U658 ( .A1(n591), .A2(n590), .ZN(n997) );
  INV_X1 U659 ( .A(G860), .ZN(n607) );
  OR2_X1 U660 ( .A1(n997), .A2(n607), .ZN(G153) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n604) );
  NAND2_X1 U662 ( .A1(n592), .A2(G54), .ZN(n593) );
  XOR2_X1 U663 ( .A(n593), .B(KEYINPUT73), .Z(n595) );
  NAND2_X1 U664 ( .A1(n657), .A2(G79), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U666 ( .A(n596), .B(KEYINPUT74), .ZN(n600) );
  NAND2_X1 U667 ( .A1(G92), .A2(n656), .ZN(n598) );
  NAND2_X1 U668 ( .A1(G66), .A2(n660), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U670 ( .A(KEYINPUT15), .B(n601), .ZN(n602) );
  XNOR2_X1 U671 ( .A(KEYINPUT75), .B(n602), .ZN(n713) );
  BUF_X1 U672 ( .A(n713), .Z(n1004) );
  OR2_X1 U673 ( .A1(n1004), .A2(G868), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n604), .A2(n603), .ZN(G284) );
  NAND2_X1 U675 ( .A1(G286), .A2(G868), .ZN(n606) );
  INV_X1 U676 ( .A(G299), .ZN(n717) );
  OR2_X1 U677 ( .A1(n717), .A2(G868), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(G297) );
  NAND2_X1 U679 ( .A1(n607), .A2(G559), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n608), .A2(n1004), .ZN(n609) );
  XNOR2_X1 U681 ( .A(n609), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U682 ( .A1(G868), .A2(n997), .ZN(n612) );
  NAND2_X1 U683 ( .A1(G868), .A2(n1004), .ZN(n610) );
  NOR2_X1 U684 ( .A1(G559), .A2(n610), .ZN(n611) );
  NOR2_X1 U685 ( .A1(n612), .A2(n611), .ZN(G282) );
  NAND2_X1 U686 ( .A1(n898), .A2(G111), .ZN(n613) );
  XOR2_X1 U687 ( .A(KEYINPUT77), .B(n613), .Z(n615) );
  NAND2_X1 U688 ( .A1(n892), .A2(G99), .ZN(n614) );
  NAND2_X1 U689 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U690 ( .A(KEYINPUT78), .B(n616), .ZN(n623) );
  NAND2_X1 U691 ( .A1(G123), .A2(n896), .ZN(n618) );
  XNOR2_X1 U692 ( .A(n618), .B(KEYINPUT18), .ZN(n621) );
  BUF_X1 U693 ( .A(n619), .Z(n890) );
  NAND2_X1 U694 ( .A1(n890), .A2(G135), .ZN(n620) );
  NAND2_X1 U695 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U696 ( .A1(n623), .A2(n622), .ZN(n924) );
  XNOR2_X1 U697 ( .A(G2096), .B(n924), .ZN(n625) );
  INV_X1 U698 ( .A(G2100), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n625), .A2(n624), .ZN(G156) );
  NAND2_X1 U700 ( .A1(G67), .A2(n660), .ZN(n627) );
  NAND2_X1 U701 ( .A1(G55), .A2(n592), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U703 ( .A1(G93), .A2(n656), .ZN(n629) );
  NAND2_X1 U704 ( .A1(G80), .A2(n657), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n670) );
  NAND2_X1 U707 ( .A1(G559), .A2(n1004), .ZN(n632) );
  XNOR2_X1 U708 ( .A(n632), .B(n997), .ZN(n673) );
  NOR2_X1 U709 ( .A1(G860), .A2(n673), .ZN(n633) );
  XOR2_X1 U710 ( .A(KEYINPUT79), .B(n633), .Z(n634) );
  XNOR2_X1 U711 ( .A(n670), .B(n634), .ZN(G145) );
  NAND2_X1 U712 ( .A1(G60), .A2(n660), .ZN(n636) );
  NAND2_X1 U713 ( .A1(G47), .A2(n592), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U715 ( .A1(G85), .A2(n656), .ZN(n637) );
  XOR2_X1 U716 ( .A(KEYINPUT66), .B(n637), .Z(n638) );
  NOR2_X1 U717 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n657), .A2(G72), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n641), .A2(n640), .ZN(G290) );
  NAND2_X1 U720 ( .A1(G48), .A2(n592), .ZN(n648) );
  NAND2_X1 U721 ( .A1(G86), .A2(n656), .ZN(n643) );
  NAND2_X1 U722 ( .A1(G61), .A2(n660), .ZN(n642) );
  NAND2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U724 ( .A1(n657), .A2(G73), .ZN(n644) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(n644), .Z(n645) );
  NOR2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U728 ( .A(n649), .B(KEYINPUT80), .ZN(G305) );
  NAND2_X1 U729 ( .A1(G49), .A2(n592), .ZN(n651) );
  NAND2_X1 U730 ( .A1(G74), .A2(G651), .ZN(n650) );
  NAND2_X1 U731 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U732 ( .A1(n660), .A2(n652), .ZN(n655) );
  NAND2_X1 U733 ( .A1(n653), .A2(G87), .ZN(n654) );
  NAND2_X1 U734 ( .A1(n655), .A2(n654), .ZN(G288) );
  NAND2_X1 U735 ( .A1(G88), .A2(n656), .ZN(n659) );
  NAND2_X1 U736 ( .A1(G75), .A2(n657), .ZN(n658) );
  NAND2_X1 U737 ( .A1(n659), .A2(n658), .ZN(n665) );
  NAND2_X1 U738 ( .A1(G62), .A2(n660), .ZN(n662) );
  NAND2_X1 U739 ( .A1(G50), .A2(n592), .ZN(n661) );
  NAND2_X1 U740 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U741 ( .A(KEYINPUT81), .B(n663), .Z(n664) );
  NOR2_X1 U742 ( .A1(n665), .A2(n664), .ZN(G166) );
  NOR2_X1 U743 ( .A1(n670), .A2(G868), .ZN(n666) );
  XNOR2_X1 U744 ( .A(KEYINPUT83), .B(n666), .ZN(n677) );
  XNOR2_X1 U745 ( .A(n717), .B(KEYINPUT19), .ZN(n668) );
  XNOR2_X1 U746 ( .A(G290), .B(G305), .ZN(n667) );
  XNOR2_X1 U747 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U748 ( .A(n670), .B(n669), .ZN(n672) );
  XNOR2_X1 U749 ( .A(G288), .B(G166), .ZN(n671) );
  XNOR2_X1 U750 ( .A(n672), .B(n671), .ZN(n907) );
  XNOR2_X1 U751 ( .A(n907), .B(n673), .ZN(n674) );
  NAND2_X1 U752 ( .A1(n674), .A2(G868), .ZN(n675) );
  XNOR2_X1 U753 ( .A(KEYINPUT82), .B(n675), .ZN(n676) );
  NAND2_X1 U754 ( .A1(n677), .A2(n676), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n678) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n678), .Z(n679) );
  NAND2_X1 U757 ( .A1(G2090), .A2(n679), .ZN(n680) );
  XNOR2_X1 U758 ( .A(KEYINPUT21), .B(n680), .ZN(n681) );
  NAND2_X1 U759 ( .A1(n681), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U760 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U761 ( .A1(G661), .A2(G483), .ZN(n691) );
  XOR2_X1 U762 ( .A(KEYINPUT22), .B(KEYINPUT84), .Z(n683) );
  NAND2_X1 U763 ( .A1(G132), .A2(G82), .ZN(n682) );
  XNOR2_X1 U764 ( .A(n683), .B(n682), .ZN(n684) );
  NAND2_X1 U765 ( .A1(n684), .A2(G96), .ZN(n685) );
  NOR2_X1 U766 ( .A1(n685), .A2(G218), .ZN(n686) );
  XNOR2_X1 U767 ( .A(n686), .B(KEYINPUT85), .ZN(n838) );
  NAND2_X1 U768 ( .A1(G2106), .A2(n838), .ZN(n690) );
  NAND2_X1 U769 ( .A1(G69), .A2(G120), .ZN(n687) );
  NOR2_X1 U770 ( .A1(G237), .A2(n687), .ZN(n688) );
  NAND2_X1 U771 ( .A1(G108), .A2(n688), .ZN(n837) );
  NAND2_X1 U772 ( .A1(G567), .A2(n837), .ZN(n689) );
  NAND2_X1 U773 ( .A1(n690), .A2(n689), .ZN(n859) );
  NOR2_X1 U774 ( .A1(n691), .A2(n859), .ZN(n692) );
  XNOR2_X1 U775 ( .A(n692), .B(KEYINPUT86), .ZN(n836) );
  NAND2_X1 U776 ( .A1(G36), .A2(n836), .ZN(G176) );
  XNOR2_X1 U777 ( .A(KEYINPUT87), .B(G166), .ZN(G303) );
  XNOR2_X1 U778 ( .A(G1981), .B(G305), .ZN(n1008) );
  NAND2_X1 U779 ( .A1(G160), .A2(G40), .ZN(n782) );
  INV_X1 U780 ( .A(KEYINPUT90), .ZN(n693) );
  NOR2_X1 U781 ( .A1(G164), .A2(G1384), .ZN(n783) );
  NAND2_X2 U782 ( .A1(n697), .A2(n783), .ZN(n745) );
  NOR2_X1 U783 ( .A1(G2084), .A2(n745), .ZN(n729) );
  NAND2_X1 U784 ( .A1(n729), .A2(G8), .ZN(n741) );
  INV_X1 U785 ( .A(G1966), .ZN(n695) );
  NAND2_X1 U786 ( .A1(n745), .A2(G8), .ZN(n694) );
  XNOR2_X2 U787 ( .A(n694), .B(KEYINPUT91), .ZN(n770) );
  NAND2_X1 U788 ( .A1(G1956), .A2(n745), .ZN(n696) );
  XNOR2_X1 U789 ( .A(KEYINPUT93), .B(n696), .ZN(n701) );
  XOR2_X1 U790 ( .A(KEYINPUT27), .B(KEYINPUT92), .Z(n699) );
  AND2_X1 U791 ( .A1(n783), .A2(n697), .ZN(n724) );
  NAND2_X1 U792 ( .A1(n724), .A2(G2072), .ZN(n698) );
  XOR2_X1 U793 ( .A(n699), .B(n698), .Z(n700) );
  NOR2_X1 U794 ( .A1(n718), .A2(n717), .ZN(n703) );
  XOR2_X1 U795 ( .A(KEYINPUT28), .B(KEYINPUT94), .Z(n702) );
  XNOR2_X1 U796 ( .A(n703), .B(n702), .ZN(n722) );
  NAND2_X1 U797 ( .A1(n724), .A2(G1996), .ZN(n704) );
  XNOR2_X1 U798 ( .A(n704), .B(KEYINPUT26), .ZN(n706) );
  NAND2_X1 U799 ( .A1(n745), .A2(G1341), .ZN(n705) );
  NAND2_X1 U800 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X2 U801 ( .A1(n997), .A2(n707), .ZN(n714) );
  NAND2_X1 U802 ( .A1(n713), .A2(n714), .ZN(n712) );
  AND2_X1 U803 ( .A1(n724), .A2(G2067), .ZN(n708) );
  XNOR2_X1 U804 ( .A(n708), .B(KEYINPUT95), .ZN(n710) );
  NAND2_X1 U805 ( .A1(n745), .A2(G1348), .ZN(n709) );
  NAND2_X1 U806 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U807 ( .A1(n712), .A2(n711), .ZN(n716) );
  OR2_X1 U808 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U809 ( .A1(n716), .A2(n715), .ZN(n720) );
  NAND2_X1 U810 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U811 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U812 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U813 ( .A(n723), .B(KEYINPUT29), .ZN(n728) );
  XOR2_X1 U814 ( .A(KEYINPUT25), .B(G2078), .Z(n947) );
  NOR2_X1 U815 ( .A1(n947), .A2(n745), .ZN(n726) );
  NOR2_X1 U816 ( .A1(n724), .A2(G1961), .ZN(n725) );
  NOR2_X1 U817 ( .A1(n726), .A2(n725), .ZN(n733) );
  NOR2_X1 U818 ( .A1(G301), .A2(n733), .ZN(n727) );
  NOR2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n738) );
  NOR2_X1 U820 ( .A1(n739), .A2(n729), .ZN(n730) );
  NAND2_X1 U821 ( .A1(n730), .A2(G8), .ZN(n731) );
  XNOR2_X1 U822 ( .A(n731), .B(KEYINPUT30), .ZN(n732) );
  NOR2_X1 U823 ( .A1(G168), .A2(n732), .ZN(n735) );
  AND2_X1 U824 ( .A1(G301), .A2(n733), .ZN(n734) );
  NOR2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U826 ( .A(n736), .B(KEYINPUT31), .ZN(n737) );
  NOR2_X2 U827 ( .A1(n738), .A2(n737), .ZN(n742) );
  NOR2_X1 U828 ( .A1(n739), .A2(n742), .ZN(n740) );
  NAND2_X1 U829 ( .A1(n741), .A2(n740), .ZN(n755) );
  INV_X1 U830 ( .A(n742), .ZN(n744) );
  AND2_X1 U831 ( .A1(G286), .A2(G8), .ZN(n743) );
  NAND2_X1 U832 ( .A1(n744), .A2(n743), .ZN(n752) );
  INV_X1 U833 ( .A(G8), .ZN(n750) );
  INV_X1 U834 ( .A(n770), .ZN(n778) );
  NOR2_X1 U835 ( .A1(G1971), .A2(n778), .ZN(n747) );
  NOR2_X1 U836 ( .A1(G2090), .A2(n745), .ZN(n746) );
  NOR2_X1 U837 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U838 ( .A1(n748), .A2(G303), .ZN(n749) );
  OR2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U841 ( .A(n753), .B(n521), .ZN(n754) );
  NAND2_X1 U842 ( .A1(n755), .A2(n754), .ZN(n776) );
  NOR2_X1 U843 ( .A1(G1971), .A2(G303), .ZN(n756) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n994) );
  NOR2_X1 U845 ( .A1(n756), .A2(n994), .ZN(n757) );
  NAND2_X1 U846 ( .A1(n776), .A2(n757), .ZN(n760) );
  NAND2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n995) );
  XNOR2_X1 U848 ( .A(n761), .B(KEYINPUT64), .ZN(n762) );
  NOR2_X1 U849 ( .A1(n1008), .A2(n765), .ZN(n768) );
  AND2_X1 U850 ( .A1(n994), .A2(KEYINPUT33), .ZN(n766) );
  NAND2_X1 U851 ( .A1(n766), .A2(n770), .ZN(n767) );
  NAND2_X1 U852 ( .A1(n768), .A2(n767), .ZN(n773) );
  NOR2_X1 U853 ( .A1(G1981), .A2(G305), .ZN(n769) );
  XNOR2_X1 U854 ( .A(n769), .B(KEYINPUT24), .ZN(n771) );
  NAND2_X1 U855 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U856 ( .A1(n773), .A2(n772), .ZN(n781) );
  NOR2_X1 U857 ( .A1(G2090), .A2(G303), .ZN(n774) );
  NAND2_X1 U858 ( .A1(G8), .A2(n774), .ZN(n775) );
  NAND2_X1 U859 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U860 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U861 ( .A(KEYINPUT98), .B(n779), .Z(n780) );
  NOR2_X1 U862 ( .A1(n781), .A2(n780), .ZN(n811) );
  NOR2_X1 U863 ( .A1(n783), .A2(n782), .ZN(n826) );
  NAND2_X1 U864 ( .A1(G104), .A2(n892), .ZN(n785) );
  NAND2_X1 U865 ( .A1(G140), .A2(n890), .ZN(n784) );
  NAND2_X1 U866 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U867 ( .A(KEYINPUT34), .B(n786), .ZN(n791) );
  NAND2_X1 U868 ( .A1(G116), .A2(n898), .ZN(n788) );
  NAND2_X1 U869 ( .A1(G128), .A2(n896), .ZN(n787) );
  NAND2_X1 U870 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U871 ( .A(KEYINPUT35), .B(n789), .Z(n790) );
  NOR2_X1 U872 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U873 ( .A(KEYINPUT36), .B(n792), .ZN(n871) );
  XNOR2_X1 U874 ( .A(G2067), .B(KEYINPUT37), .ZN(n822) );
  NOR2_X1 U875 ( .A1(n871), .A2(n822), .ZN(n925) );
  NAND2_X1 U876 ( .A1(n826), .A2(n925), .ZN(n820) );
  INV_X1 U877 ( .A(n820), .ZN(n810) );
  NAND2_X1 U878 ( .A1(G117), .A2(n898), .ZN(n794) );
  NAND2_X1 U879 ( .A1(G129), .A2(n896), .ZN(n793) );
  NAND2_X1 U880 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U881 ( .A1(n892), .A2(G105), .ZN(n795) );
  XOR2_X1 U882 ( .A(KEYINPUT38), .B(n795), .Z(n796) );
  NOR2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n799) );
  NAND2_X1 U884 ( .A1(n890), .A2(G141), .ZN(n798) );
  NAND2_X1 U885 ( .A1(n799), .A2(n798), .ZN(n873) );
  NAND2_X1 U886 ( .A1(G1996), .A2(n873), .ZN(n808) );
  NAND2_X1 U887 ( .A1(G107), .A2(n898), .ZN(n801) );
  NAND2_X1 U888 ( .A1(G119), .A2(n896), .ZN(n800) );
  NAND2_X1 U889 ( .A1(n801), .A2(n800), .ZN(n804) );
  NAND2_X1 U890 ( .A1(n892), .A2(G95), .ZN(n802) );
  XOR2_X1 U891 ( .A(KEYINPUT88), .B(n802), .Z(n803) );
  NOR2_X1 U892 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U893 ( .A1(n890), .A2(G131), .ZN(n805) );
  NAND2_X1 U894 ( .A1(n806), .A2(n805), .ZN(n870) );
  NAND2_X1 U895 ( .A1(G1991), .A2(n870), .ZN(n807) );
  NAND2_X1 U896 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U897 ( .A(KEYINPUT89), .B(n809), .Z(n919) );
  OR2_X2 U898 ( .A1(n811), .A2(n520), .ZN(n812) );
  XNOR2_X1 U899 ( .A(n812), .B(KEYINPUT99), .ZN(n814) );
  XNOR2_X1 U900 ( .A(G1986), .B(G290), .ZN(n993) );
  NAND2_X1 U901 ( .A1(n826), .A2(n993), .ZN(n813) );
  NAND2_X1 U902 ( .A1(n814), .A2(n813), .ZN(n829) );
  NOR2_X1 U903 ( .A1(n873), .A2(G1996), .ZN(n815) );
  XNOR2_X1 U904 ( .A(n815), .B(KEYINPUT100), .ZN(n934) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n870), .ZN(n923) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U907 ( .A1(n923), .A2(n816), .ZN(n817) );
  NOR2_X1 U908 ( .A1(n919), .A2(n817), .ZN(n818) );
  NOR2_X1 U909 ( .A1(n934), .A2(n818), .ZN(n819) );
  XNOR2_X1 U910 ( .A(n819), .B(KEYINPUT39), .ZN(n821) );
  NAND2_X1 U911 ( .A1(n821), .A2(n820), .ZN(n823) );
  NAND2_X1 U912 ( .A1(n871), .A2(n822), .ZN(n920) );
  NAND2_X1 U913 ( .A1(n823), .A2(n920), .ZN(n824) );
  XOR2_X1 U914 ( .A(KEYINPUT101), .B(n824), .Z(n825) );
  NAND2_X1 U915 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U916 ( .A(n827), .B(KEYINPUT102), .ZN(n828) );
  NAND2_X1 U917 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U918 ( .A(KEYINPUT40), .B(n830), .ZN(G329) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n831), .ZN(G217) );
  NAND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n833) );
  INV_X1 U921 ( .A(G661), .ZN(n832) );
  NOR2_X1 U922 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U923 ( .A(n834), .B(KEYINPUT103), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U925 ( .A1(n836), .A2(n835), .ZN(G188) );
  INV_X1 U927 ( .A(G132), .ZN(G219) );
  INV_X1 U928 ( .A(G120), .ZN(G236) );
  INV_X1 U929 ( .A(G96), .ZN(G221) );
  INV_X1 U930 ( .A(G82), .ZN(G220) );
  INV_X1 U931 ( .A(G69), .ZN(G235) );
  NOR2_X1 U932 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  XOR2_X1 U934 ( .A(KEYINPUT105), .B(G2084), .Z(n840) );
  XNOR2_X1 U935 ( .A(G2090), .B(G2072), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U937 ( .A(n841), .B(G2096), .Z(n843) );
  XNOR2_X1 U938 ( .A(G2078), .B(G2067), .ZN(n842) );
  XNOR2_X1 U939 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U940 ( .A(KEYINPUT43), .B(G2678), .Z(n845) );
  XNOR2_X1 U941 ( .A(G2100), .B(KEYINPUT42), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U943 ( .A(n847), .B(n846), .Z(G227) );
  XOR2_X1 U944 ( .A(KEYINPUT41), .B(G1966), .Z(n849) );
  XNOR2_X1 U945 ( .A(G1981), .B(G1961), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U947 ( .A(n850), .B(KEYINPUT106), .Z(n852) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U950 ( .A(G1956), .B(G1971), .Z(n854) );
  XNOR2_X1 U951 ( .A(G1986), .B(G1976), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U953 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U954 ( .A(KEYINPUT107), .B(G2474), .ZN(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(G229) );
  XOR2_X1 U956 ( .A(KEYINPUT104), .B(n859), .Z(G319) );
  NAND2_X1 U957 ( .A1(n890), .A2(G136), .ZN(n860) );
  XNOR2_X1 U958 ( .A(KEYINPUT108), .B(n860), .ZN(n863) );
  NAND2_X1 U959 ( .A1(n896), .A2(G124), .ZN(n861) );
  XNOR2_X1 U960 ( .A(KEYINPUT44), .B(n861), .ZN(n862) );
  NAND2_X1 U961 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U962 ( .A(n864), .B(KEYINPUT109), .ZN(n866) );
  NAND2_X1 U963 ( .A1(G112), .A2(n898), .ZN(n865) );
  NAND2_X1 U964 ( .A1(n866), .A2(n865), .ZN(n869) );
  NAND2_X1 U965 ( .A1(n892), .A2(G100), .ZN(n867) );
  XOR2_X1 U966 ( .A(KEYINPUT110), .B(n867), .Z(n868) );
  NOR2_X1 U967 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U968 ( .A(n871), .B(n870), .Z(n872) );
  XNOR2_X1 U969 ( .A(n873), .B(n872), .ZN(n882) );
  NAND2_X1 U970 ( .A1(G118), .A2(n898), .ZN(n875) );
  NAND2_X1 U971 ( .A1(G130), .A2(n896), .ZN(n874) );
  NAND2_X1 U972 ( .A1(n875), .A2(n874), .ZN(n880) );
  NAND2_X1 U973 ( .A1(G106), .A2(n892), .ZN(n877) );
  NAND2_X1 U974 ( .A1(G142), .A2(n890), .ZN(n876) );
  NAND2_X1 U975 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U976 ( .A(n878), .B(KEYINPUT45), .Z(n879) );
  NOR2_X1 U977 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U978 ( .A(n882), .B(n881), .Z(n889) );
  XOR2_X1 U979 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n884) );
  XNOR2_X1 U980 ( .A(KEYINPUT114), .B(KEYINPUT48), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U982 ( .A(n885), .B(n924), .Z(n887) );
  XNOR2_X1 U983 ( .A(G164), .B(G160), .ZN(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U985 ( .A(n889), .B(n888), .Z(n905) );
  NAND2_X1 U986 ( .A1(G139), .A2(n890), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n891), .B(KEYINPUT112), .ZN(n895) );
  NAND2_X1 U988 ( .A1(G103), .A2(n892), .ZN(n893) );
  XOR2_X1 U989 ( .A(KEYINPUT111), .B(n893), .Z(n894) );
  NAND2_X1 U990 ( .A1(n895), .A2(n894), .ZN(n903) );
  NAND2_X1 U991 ( .A1(n896), .A2(G127), .ZN(n897) );
  XOR2_X1 U992 ( .A(KEYINPUT113), .B(n897), .Z(n900) );
  NAND2_X1 U993 ( .A1(n898), .A2(G115), .ZN(n899) );
  NAND2_X1 U994 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U995 ( .A(KEYINPUT47), .B(n901), .Z(n902) );
  NOR2_X1 U996 ( .A1(n903), .A2(n902), .ZN(n929) );
  XNOR2_X1 U997 ( .A(n929), .B(G162), .ZN(n904) );
  XNOR2_X1 U998 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U999 ( .A1(G37), .A2(n906), .ZN(G395) );
  XNOR2_X1 U1000 ( .A(n997), .B(n907), .ZN(n909) );
  XNOR2_X1 U1001 ( .A(G171), .B(n1004), .ZN(n908) );
  XNOR2_X1 U1002 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1003 ( .A(G286), .B(n910), .Z(n911) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n911), .ZN(G397) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(n912), .B(KEYINPUT49), .ZN(n916) );
  INV_X1 U1007 ( .A(G319), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(n913), .A2(G401), .ZN(n914) );
  XOR2_X1 U1009 ( .A(KEYINPUT116), .B(n914), .Z(n915) );
  NOR2_X1 U1010 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1015 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n1025) );
  INV_X1 U1016 ( .A(n919), .ZN(n921) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n941) );
  XOR2_X1 U1018 ( .A(G2084), .B(G160), .Z(n922) );
  NOR2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n927) );
  NOR2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1021 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1022 ( .A(KEYINPUT117), .B(n928), .ZN(n939) );
  XOR2_X1 U1023 ( .A(G2072), .B(n929), .Z(n931) );
  XOR2_X1 U1024 ( .A(G164), .B(G2078), .Z(n930) );
  NOR2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1026 ( .A(KEYINPUT50), .B(n932), .Z(n937) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n933) );
  NOR2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1029 ( .A(KEYINPUT51), .B(n935), .ZN(n936) );
  NOR2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1031 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1032 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1033 ( .A(KEYINPUT52), .B(n942), .ZN(n944) );
  INV_X1 U1034 ( .A(KEYINPUT55), .ZN(n943) );
  NAND2_X1 U1035 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1036 ( .A1(n945), .A2(G29), .ZN(n946) );
  XNOR2_X1 U1037 ( .A(KEYINPUT118), .B(n946), .ZN(n1023) );
  XNOR2_X1 U1038 ( .A(G1991), .B(G25), .ZN(n958) );
  XOR2_X1 U1039 ( .A(G2072), .B(G33), .Z(n952) );
  XNOR2_X1 U1040 ( .A(n947), .B(G27), .ZN(n949) );
  XNOR2_X1 U1041 ( .A(G32), .B(G1996), .ZN(n948) );
  NOR2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(KEYINPUT120), .B(n950), .ZN(n951) );
  NAND2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n955) );
  XOR2_X1 U1045 ( .A(G26), .B(G2067), .Z(n953) );
  XNOR2_X1 U1046 ( .A(KEYINPUT119), .B(n953), .ZN(n954) );
  NOR2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(KEYINPUT121), .B(n956), .ZN(n957) );
  NOR2_X1 U1049 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1050 ( .A1(G28), .A2(n959), .ZN(n960) );
  XNOR2_X1 U1051 ( .A(n960), .B(KEYINPUT53), .ZN(n963) );
  XOR2_X1 U1052 ( .A(G2084), .B(G34), .Z(n961) );
  XNOR2_X1 U1053 ( .A(KEYINPUT54), .B(n961), .ZN(n962) );
  NAND2_X1 U1054 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1055 ( .A(G35), .B(G2090), .ZN(n964) );
  NOR2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1057 ( .A(KEYINPUT55), .B(n966), .Z(n967) );
  NOR2_X1 U1058 ( .A1(G29), .A2(n967), .ZN(n1021) );
  XOR2_X1 U1059 ( .A(G1961), .B(G5), .Z(n977) );
  XNOR2_X1 U1060 ( .A(G1348), .B(KEYINPUT59), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(n968), .B(G4), .ZN(n972) );
  XNOR2_X1 U1062 ( .A(G1981), .B(G6), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(G1341), .B(G19), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(G20), .B(G1956), .ZN(n973) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(KEYINPUT60), .B(n975), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(G21), .B(G1966), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1072 ( .A(KEYINPUT123), .B(n980), .Z(n988) );
  XOR2_X1 U1073 ( .A(G1971), .B(G22), .Z(n983) );
  XOR2_X1 U1074 ( .A(G24), .B(KEYINPUT124), .Z(n981) );
  XNOR2_X1 U1075 ( .A(n981), .B(G1986), .ZN(n982) );
  NAND2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(G23), .B(G1976), .ZN(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(KEYINPUT58), .B(n986), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1081 ( .A(n989), .B(KEYINPUT125), .Z(n990) );
  XNOR2_X1 U1082 ( .A(KEYINPUT61), .B(n990), .ZN(n991) );
  NOR2_X1 U1083 ( .A1(G16), .A2(n991), .ZN(n1017) );
  XOR2_X1 U1084 ( .A(G16), .B(KEYINPUT56), .Z(n1015) );
  XNOR2_X1 U1085 ( .A(G1971), .B(KEYINPUT122), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(n992), .B(G303), .ZN(n1013) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n996) );
  NAND2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(G1341), .B(n997), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(G301), .B(G1961), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(G299), .B(G1956), .ZN(n1000) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1006) );
  XOR2_X1 U1095 ( .A(G1348), .B(n1004), .Z(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1011) );
  XOR2_X1 U1097 ( .A(G168), .B(G1966), .Z(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1099 ( .A(KEYINPUT57), .B(n1009), .Z(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(n1018), .B(KEYINPUT126), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(G11), .A2(n1019), .ZN(n1020) );
  NOR2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(n1025), .B(n1024), .ZN(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

