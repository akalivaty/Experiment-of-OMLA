//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1263, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G107), .ZN(new_n227));
  INV_X1    g0027(.A(G264), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n212), .B1(new_n215), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT64), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n202), .A2(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n219), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n244), .B(new_n249), .ZN(G351));
  NAND2_X1  g0050(.A1(new_n206), .A2(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G50), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT68), .ZN(new_n253));
  INV_X1    g0053(.A(G13), .ZN(new_n254));
  NOR3_X1   g0054(.A1(new_n254), .A2(new_n207), .A3(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n213), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n255), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n253), .A2(new_n259), .B1(G50), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n257), .ZN(new_n262));
  XOR2_X1   g0062(.A(KEYINPUT8), .B(G58), .Z(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n263), .A2(new_n265), .B1(G150), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n203), .A2(G20), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n262), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n261), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT65), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n213), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(KEYINPUT65), .A2(G33), .A3(G41), .ZN(new_n275));
  AOI21_X1  g0075(.A(KEYINPUT66), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(new_n272), .ZN(new_n277));
  INV_X1    g0077(.A(new_n213), .ZN(new_n278));
  AND4_X1   g0078(.A1(KEYINPUT66), .A2(new_n277), .A3(new_n278), .A4(new_n275), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n271), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT67), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n277), .A2(new_n278), .A3(new_n275), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT66), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n274), .A2(KEYINPUT66), .A3(new_n275), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT67), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(new_n287), .A3(new_n271), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n281), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G226), .ZN(new_n290));
  INV_X1    g0090(.A(new_n271), .ZN(new_n291));
  OAI211_X1 g0091(.A(G274), .B(new_n291), .C1(new_n276), .C2(new_n279), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT3), .B(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G222), .A2(G1698), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(G223), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n294), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n278), .A2(new_n273), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT3), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n299), .B1(new_n303), .B2(new_n225), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n293), .B1(new_n298), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n290), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n270), .B1(new_n307), .B2(G169), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n308), .A2(KEYINPUT69), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(KEYINPUT69), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n306), .A2(G179), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n311), .A2(KEYINPUT70), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(KEYINPUT70), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n309), .A2(new_n310), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n270), .B(KEYINPUT9), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n306), .A2(G200), .ZN(new_n316));
  INV_X1    g0116(.A(G190), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n315), .B(new_n316), .C1(new_n317), .C2(new_n306), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT10), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n263), .A2(new_n251), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n259), .A2(new_n321), .B1(new_n260), .B2(new_n263), .ZN(new_n322));
  INV_X1    g0122(.A(G58), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n219), .ZN(new_n324));
  OR2_X1    g0124(.A1(new_n324), .A2(new_n201), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n325), .A2(G20), .B1(G159), .B2(new_n266), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT7), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT75), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n264), .B2(KEYINPUT3), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n300), .A2(KEYINPUT75), .A3(G33), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n330), .A2(new_n331), .A3(new_n302), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n328), .B1(new_n332), .B2(G20), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n330), .A2(new_n331), .A3(new_n302), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(KEYINPUT76), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT7), .B1(new_n334), .B2(new_n207), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT76), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n219), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n327), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n262), .B1(new_n340), .B2(KEYINPUT16), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT16), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n328), .B1(new_n294), .B2(G20), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n303), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n219), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n326), .B1(new_n345), .B2(KEYINPUT77), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT77), .ZN(new_n347));
  AOI211_X1 g0147(.A(new_n347), .B(new_n219), .C1(new_n343), .C2(new_n344), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n342), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n322), .B1(new_n341), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n286), .A2(G232), .A3(new_n271), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G87), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT78), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n352), .B(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G226), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G1698), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(G223), .B2(G1698), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n354), .B1(new_n334), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n299), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n351), .A2(new_n292), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G169), .ZN(new_n362));
  INV_X1    g0162(.A(G179), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n362), .B1(new_n363), .B2(new_n361), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT18), .B1(new_n350), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G200), .ZN(new_n367));
  INV_X1    g0167(.A(G274), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n284), .B2(new_n285), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n369), .A2(new_n291), .B1(new_n359), .B2(new_n358), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n367), .B1(new_n370), .B2(new_n351), .ZN(new_n371));
  AND4_X1   g0171(.A1(G190), .A2(new_n351), .A3(new_n292), .A4(new_n360), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n335), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n374), .A2(new_n337), .A3(new_n338), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n338), .B(new_n328), .C1(new_n332), .C2(G20), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G68), .ZN(new_n377));
  OAI211_X1 g0177(.A(KEYINPUT16), .B(new_n326), .C1(new_n375), .C2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n378), .A2(new_n349), .A3(new_n257), .ZN(new_n379));
  INV_X1    g0179(.A(new_n322), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n373), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT17), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n379), .A2(new_n380), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT18), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(new_n364), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n373), .A2(new_n379), .A3(KEYINPUT17), .A4(new_n380), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n366), .A2(new_n383), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n289), .A2(G244), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n294), .A2(G232), .A3(new_n296), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n294), .A2(G238), .A3(G1698), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n390), .B(new_n391), .C1(new_n227), .C2(new_n294), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n293), .B1(new_n359), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n363), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n258), .A2(G77), .A3(new_n251), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(G77), .B2(new_n260), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n263), .A2(new_n266), .B1(G20), .B2(G77), .ZN(new_n399));
  XNOR2_X1  g0199(.A(KEYINPUT15), .B(G87), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n265), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n262), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G169), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n394), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n396), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n394), .A2(new_n317), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT71), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n404), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n411), .B1(new_n394), .B2(G200), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n413), .A2(new_n409), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n408), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  OR3_X1    g0215(.A1(new_n320), .A2(new_n388), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n220), .B1(new_n281), .B2(new_n288), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n301), .A2(new_n302), .A3(G232), .A4(G1698), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G97), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT72), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n355), .A2(G1698), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n294), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n301), .A3(new_n302), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT72), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n420), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n292), .B1(new_n426), .B2(new_n299), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT13), .B1(new_n417), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n287), .B1(new_n286), .B2(new_n271), .ZN(new_n429));
  AOI211_X1 g0229(.A(KEYINPUT67), .B(new_n291), .C1(new_n284), .C2(new_n285), .ZN(new_n430));
  OAI21_X1  g0230(.A(G238), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT13), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n425), .A2(new_n423), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n433), .A2(new_n419), .A3(new_n418), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n434), .A2(new_n359), .B1(new_n369), .B2(new_n291), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n431), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n428), .A2(KEYINPUT73), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n427), .B1(new_n289), .B2(G238), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT73), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n439), .A3(new_n432), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n437), .A2(G200), .A3(new_n440), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n266), .A2(G50), .B1(G20), .B2(new_n219), .ZN(new_n442));
  INV_X1    g0242(.A(new_n265), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n443), .B2(new_n225), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n257), .ZN(new_n445));
  XOR2_X1   g0245(.A(new_n445), .B(KEYINPUT11), .Z(new_n446));
  NAND3_X1  g0246(.A1(new_n258), .A2(G68), .A3(new_n251), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n254), .A2(G1), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(G20), .A3(new_n219), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT74), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT12), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n450), .A2(KEYINPUT12), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n447), .B(new_n453), .C1(new_n451), .C2(new_n449), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n446), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n317), .B1(new_n438), .B2(new_n432), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(new_n428), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n441), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n428), .A2(G179), .A3(new_n436), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n437), .A2(G169), .A3(new_n440), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT14), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n437), .A2(KEYINPUT14), .A3(G169), .A4(new_n440), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n459), .B1(new_n466), .B2(new_n455), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n416), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n222), .A2(new_n296), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n470), .B1(G257), .B2(new_n296), .ZN(new_n471));
  INV_X1    g0271(.A(G294), .ZN(new_n472));
  OAI22_X1  g0272(.A1(new_n334), .A2(new_n471), .B1(new_n264), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT88), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI221_X1 g0275(.A(KEYINPUT88), .B1(new_n264), .B2(new_n472), .C1(new_n334), .C2(new_n471), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n359), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT89), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n475), .A2(KEYINPUT89), .A3(new_n476), .A4(new_n359), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n206), .A2(G45), .ZN(new_n482));
  OR2_X1    g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  NAND2_X1  g0283(.A1(KEYINPUT5), .A2(G41), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n369), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n485), .B1(new_n284), .B2(new_n285), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G264), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n481), .A2(new_n317), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n477), .A2(new_n486), .A3(new_n488), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n367), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n255), .A2(new_n227), .ZN(new_n494));
  XNOR2_X1  g0294(.A(new_n494), .B(KEYINPUT25), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n258), .B1(G1), .B2(new_n264), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n495), .B1(new_n497), .B2(G107), .ZN(new_n498));
  NOR4_X1   g0298(.A1(new_n303), .A2(KEYINPUT22), .A3(G20), .A4(new_n221), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT22), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n330), .A2(new_n331), .A3(new_n207), .A4(new_n302), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n221), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT85), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n500), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(KEYINPUT85), .B1(new_n501), .B2(new_n221), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n499), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT23), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(new_n227), .A3(G20), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n507), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  XNOR2_X1  g0311(.A(new_n511), .B(KEYINPUT86), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT24), .B1(new_n506), .B2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n332), .A2(new_n503), .A3(new_n207), .A4(G87), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(KEYINPUT22), .A3(new_n505), .ZN(new_n515));
  INV_X1    g0315(.A(new_n499), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT24), .ZN(new_n518));
  INV_X1    g0318(.A(new_n512), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT87), .B1(new_n521), .B2(new_n257), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT87), .ZN(new_n523));
  AOI211_X1 g0323(.A(new_n523), .B(new_n262), .C1(new_n513), .C2(new_n520), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n493), .B(new_n498), .C1(new_n522), .C2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n260), .A2(G97), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(new_n497), .B2(G97), .ZN(new_n527));
  INV_X1    g0327(.A(G97), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n227), .B1(new_n528), .B2(KEYINPUT6), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT6), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(G97), .A3(G107), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n528), .A2(KEYINPUT79), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT79), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G97), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n535), .A3(KEYINPUT6), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n532), .A2(new_n536), .A3(G20), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n266), .A2(G77), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT80), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT80), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n537), .A2(new_n541), .A3(new_n538), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n343), .A2(new_n344), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G107), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n540), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n545), .A2(KEYINPUT81), .A3(new_n257), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT81), .B1(new_n545), .B2(new_n257), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n527), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT4), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n296), .A2(G244), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n334), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G283), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n549), .A2(new_n226), .A3(G1698), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n222), .A2(new_n296), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n294), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n551), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n359), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n487), .A2(G257), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n486), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G169), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n363), .B2(new_n559), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n548), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n548), .A2(KEYINPUT82), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT81), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n537), .A2(new_n541), .A3(new_n538), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n541), .B1(new_n537), .B2(new_n538), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n227), .B1(new_n343), .B2(new_n344), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n564), .B1(new_n568), .B2(new_n262), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n545), .A2(KEYINPUT81), .A3(new_n257), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT82), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n572), .A3(new_n527), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n559), .A2(new_n317), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(G200), .B2(new_n559), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n563), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n332), .A2(KEYINPUT84), .A3(new_n207), .A4(G68), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT84), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n501), .B2(new_n219), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT83), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n533), .A2(new_n535), .A3(new_n221), .A4(new_n227), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT19), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n207), .B1(new_n419), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n581), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n582), .A2(new_n581), .A3(new_n584), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n533), .A2(new_n535), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT19), .B1(new_n588), .B2(new_n265), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n586), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n257), .B1(new_n580), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n401), .A2(new_n260), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n497), .A2(G87), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(G238), .A2(G1698), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n226), .B2(G1698), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n598), .A2(new_n330), .A3(new_n331), .A4(new_n302), .ZN(new_n599));
  NAND2_X1  g0399(.A1(G33), .A2(G116), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n299), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n482), .A2(new_n222), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(G274), .B2(new_n482), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(new_n284), .B2(new_n285), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n601), .A2(new_n604), .A3(new_n317), .ZN(new_n605));
  INV_X1    g0405(.A(new_n603), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n286), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n226), .A2(G1698), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(G238), .B2(G1698), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n600), .B1(new_n334), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n359), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n367), .B1(new_n607), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n497), .A2(new_n401), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n592), .A2(new_n594), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(G169), .B1(new_n607), .B2(new_n611), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n601), .A2(new_n604), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n616), .B1(new_n363), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n596), .A2(new_n613), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n525), .A2(new_n562), .A3(new_n576), .A4(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n533), .A2(new_n535), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n207), .B(new_n552), .C1(new_n621), .C2(G33), .ZN(new_n622));
  INV_X1    g0422(.A(G116), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n262), .B1(G20), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT20), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n622), .A2(new_n624), .A3(KEYINPUT20), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n255), .A2(new_n623), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n496), .B2(new_n623), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n487), .A2(G270), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n228), .A2(G1698), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(G257), .B2(G1698), .ZN(new_n636));
  INV_X1    g0436(.A(G303), .ZN(new_n637));
  OAI22_X1  g0437(.A1(new_n334), .A2(new_n636), .B1(new_n637), .B2(new_n294), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n359), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n486), .A2(new_n634), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n633), .A2(G169), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT21), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n633), .A2(KEYINPUT21), .A3(G169), .A4(new_n640), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n631), .B1(new_n627), .B2(new_n628), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n486), .A2(new_n634), .A3(G179), .A4(new_n639), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n640), .A2(G200), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n648), .B(new_n645), .C1(new_n317), .C2(new_n640), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n643), .A2(new_n644), .A3(new_n647), .A4(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n498), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n518), .B1(new_n517), .B2(new_n519), .ZN(new_n652));
  AOI211_X1 g0452(.A(KEYINPUT24), .B(new_n512), .C1(new_n515), .C2(new_n516), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n257), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n523), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n521), .A2(KEYINPUT87), .A3(new_n257), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OR3_X1    g0457(.A1(new_n491), .A2(KEYINPUT90), .A3(new_n363), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT90), .B1(new_n491), .B2(new_n363), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n406), .B1(new_n481), .B2(new_n489), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n650), .B1(new_n657), .B2(new_n662), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n469), .A2(new_n620), .A3(new_n663), .ZN(G372));
  NOR2_X1   g0464(.A1(new_n466), .A2(new_n455), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n408), .B1(new_n441), .B2(new_n458), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n383), .B(new_n387), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n366), .A2(new_n386), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n319), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n670), .A2(new_n314), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n643), .A2(new_n644), .A3(new_n647), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n498), .B1(new_n522), .B2(new_n524), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n481), .A2(new_n489), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n659), .B(new_n658), .C1(new_n674), .C2(new_n406), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n672), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n620), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n615), .A2(new_n618), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n613), .A2(new_n594), .A3(new_n592), .A4(new_n595), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n548), .A2(new_n678), .A3(new_n561), .A4(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n679), .B1(new_n681), .B2(KEYINPUT26), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n572), .B1(new_n571), .B2(new_n527), .ZN(new_n683));
  INV_X1    g0483(.A(new_n527), .ZN(new_n684));
  AOI211_X1 g0484(.A(KEYINPUT82), .B(new_n684), .C1(new_n569), .C2(new_n570), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n561), .B(new_n619), .C1(new_n683), .C2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n682), .B1(new_n686), .B2(KEYINPUT26), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n468), .B1(new_n677), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n671), .A2(new_n688), .ZN(G369));
  NAND2_X1  g0489(.A1(new_n448), .A2(new_n207), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G213), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n645), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n672), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n643), .A2(new_n644), .A3(new_n647), .A4(new_n649), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n698), .B(KEYINPUT91), .C1(new_n699), .C2(new_n697), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(KEYINPUT91), .B2(new_n698), .ZN(new_n701));
  INV_X1    g0501(.A(G330), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n525), .B1(new_n657), .B2(new_n696), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n673), .A2(new_n675), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n673), .A2(new_n675), .A3(new_n696), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n707), .ZN(new_n711));
  INV_X1    g0511(.A(new_n672), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n695), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n711), .B1(new_n706), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n710), .A2(new_n714), .ZN(G399));
  INV_X1    g0515(.A(new_n210), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n582), .A2(G116), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G1), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n217), .B2(new_n718), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n576), .A2(new_n562), .A3(new_n619), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n699), .B1(new_n673), .B2(new_n675), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n723), .A2(new_n724), .A3(new_n525), .A4(new_n696), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n617), .A2(new_n557), .A3(new_n558), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n491), .A2(new_n726), .A3(new_n646), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT92), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT30), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n557), .A2(new_n558), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(new_n489), .A3(new_n477), .A4(new_n617), .ZN(new_n732));
  OAI211_X1 g0532(.A(KEYINPUT92), .B(new_n730), .C1(new_n732), .C2(new_n646), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n617), .A2(G179), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n491), .A2(new_n734), .A3(new_n559), .A4(new_n640), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n729), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT31), .B1(new_n736), .B2(new_n695), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n702), .B1(new_n725), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n696), .B1(new_n677), .B2(new_n687), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT93), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT29), .ZN(new_n744));
  OAI211_X1 g0544(.A(KEYINPUT93), .B(new_n696), .C1(new_n677), .C2(new_n687), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT26), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT94), .B1(new_n681), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(new_n686), .B2(new_n747), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n731), .A2(G179), .A3(new_n486), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n563), .A2(new_n573), .B1(new_n560), .B2(new_n750), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n751), .A2(KEYINPUT94), .A3(KEYINPUT26), .A4(new_n619), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n749), .A2(new_n678), .A3(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT95), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n749), .A2(new_n752), .A3(KEYINPUT95), .A4(new_n678), .ZN(new_n756));
  INV_X1    g0556(.A(new_n620), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT96), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n676), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n712), .B1(new_n657), .B2(new_n662), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(KEYINPUT96), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n757), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n755), .A2(new_n756), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(KEYINPUT29), .A3(new_n696), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n740), .B1(new_n746), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n722), .B1(new_n765), .B2(G1), .ZN(G364));
  NOR2_X1   g0566(.A1(new_n254), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n206), .B1(new_n767), .B2(G45), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n717), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n703), .A2(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n701), .A2(new_n702), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n701), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n210), .A2(G355), .A3(new_n294), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n716), .A2(new_n332), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(G45), .B2(new_n217), .ZN(new_n780));
  INV_X1    g0580(.A(G45), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n249), .A2(new_n781), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n778), .B1(G116), .B2(new_n210), .C1(new_n780), .C2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n207), .B1(KEYINPUT97), .B2(new_n406), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n406), .A2(KEYINPUT97), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n213), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n776), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n771), .B1(new_n783), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n207), .A2(new_n363), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n789), .A2(new_n317), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(KEYINPUT33), .B(G317), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n207), .A2(G179), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n793), .A2(G190), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n791), .A2(new_n792), .B1(new_n795), .B2(G303), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n317), .A2(G200), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n207), .B1(new_n797), .B2(new_n363), .ZN(new_n798));
  INV_X1    g0598(.A(G326), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n789), .A2(G190), .A3(G200), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n796), .B1(new_n472), .B2(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n789), .A2(new_n797), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G190), .A2(G200), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n793), .A2(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G322), .A2(new_n802), .B1(new_n804), .B2(G329), .ZN(new_n805));
  INV_X1    g0605(.A(G311), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n789), .A2(new_n803), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n805), .B(new_n303), .C1(new_n806), .C2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n801), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n793), .A2(new_n317), .A3(G200), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT98), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G283), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n804), .A2(G159), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n815), .A2(KEYINPUT32), .B1(new_n795), .B2(G87), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n219), .B2(new_n790), .ZN(new_n817));
  INV_X1    g0617(.A(new_n802), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n294), .B1(new_n808), .B2(new_n225), .C1(new_n323), .C2(new_n818), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n815), .A2(KEYINPUT32), .B1(new_n202), .B2(new_n800), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n812), .A2(new_n227), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n798), .B(KEYINPUT99), .Z(new_n823));
  AOI21_X1  g0623(.A(new_n822), .B1(G97), .B2(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n810), .A2(new_n814), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n786), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n788), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n772), .A2(new_n773), .B1(new_n777), .B2(new_n827), .ZN(G396));
  NOR2_X1   g0628(.A1(new_n408), .A2(new_n695), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n412), .A2(new_n414), .B1(new_n404), .B2(new_n696), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n829), .B1(new_n830), .B2(new_n408), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n743), .A2(new_n745), .A3(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n831), .B(new_n696), .C1(new_n677), .C2(new_n687), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n740), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n770), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n833), .A2(new_n740), .A3(new_n834), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n786), .A2(new_n774), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n771), .B1(new_n839), .B2(new_n225), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n800), .A2(new_n637), .B1(new_n794), .B2(new_n227), .ZN(new_n841));
  INV_X1    g0641(.A(new_n804), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n303), .B1(new_n842), .B2(new_n806), .C1(new_n818), .C2(new_n472), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n841), .B(new_n843), .C1(G97), .C2(new_n823), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n813), .A2(G87), .ZN(new_n845));
  XNOR2_X1  g0645(.A(KEYINPUT100), .B(G283), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n808), .A2(new_n623), .B1(new_n790), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n845), .B1(KEYINPUT101), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(KEYINPUT101), .B2(new_n847), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G143), .A2(new_n802), .B1(new_n807), .B2(G159), .ZN(new_n850));
  INV_X1    g0650(.A(G137), .ZN(new_n851));
  INV_X1    g0651(.A(G150), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n850), .B1(new_n851), .B2(new_n800), .C1(new_n852), .C2(new_n790), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT34), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n813), .A2(G68), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n334), .B1(G132), .B2(new_n804), .ZN(new_n857));
  INV_X1    g0657(.A(new_n798), .ZN(new_n858));
  AOI22_X1  g0658(.A1(G58), .A2(new_n858), .B1(new_n795), .B2(G50), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n853), .A2(new_n854), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n844), .A2(new_n849), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n840), .B1(new_n826), .B2(new_n863), .C1(new_n831), .C2(new_n775), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n838), .A2(new_n864), .ZN(G384));
  INV_X1    g0665(.A(KEYINPUT40), .ZN(new_n866));
  AOI221_X4 g0666(.A(new_n461), .B1(new_n441), .B2(new_n458), .C1(new_n464), .C2(new_n465), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n455), .A2(new_n696), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT102), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n459), .B(new_n869), .C1(new_n466), .C2(new_n455), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n464), .A2(new_n465), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(new_n460), .A3(new_n459), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT102), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n873), .A2(new_n874), .A3(new_n868), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n870), .A2(new_n871), .A3(new_n875), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n620), .A2(new_n663), .A3(new_n695), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n736), .A2(new_n695), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT31), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT104), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT104), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n725), .A2(new_n739), .A3(new_n884), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n876), .A2(new_n831), .A3(new_n883), .A4(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n326), .B1(new_n375), .B2(new_n377), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n342), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n322), .B1(new_n341), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n381), .B1(new_n889), .B2(new_n693), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n365), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n384), .A2(new_n364), .ZN(new_n893));
  INV_X1    g0693(.A(new_n693), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n384), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n893), .A2(new_n895), .A3(new_n896), .A4(new_n381), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n889), .A2(new_n693), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n388), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n898), .A2(new_n900), .A3(KEYINPUT38), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n866), .B1(new_n886), .B2(new_n906), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n898), .A2(KEYINPUT38), .A3(new_n900), .ZN(new_n908));
  XOR2_X1   g0708(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n381), .B1(new_n350), .B2(new_n365), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n350), .A2(new_n693), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT37), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n897), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n388), .A2(new_n912), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n910), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT105), .B1(new_n908), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT105), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n897), .A2(new_n913), .B1(new_n388), .B2(new_n912), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n904), .B(new_n918), .C1(new_n919), .C2(new_n910), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n917), .A2(KEYINPUT40), .A3(new_n920), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n725), .A2(new_n884), .A3(new_n739), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n884), .B1(new_n725), .B2(new_n739), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n875), .A2(new_n871), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n874), .B1(new_n873), .B2(new_n868), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n831), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n921), .A2(new_n924), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n907), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n468), .A2(new_n924), .ZN(new_n931));
  OAI21_X1  g0731(.A(G330), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n931), .B2(new_n930), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n746), .A2(new_n764), .A3(new_n468), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n671), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n875), .A2(new_n871), .ZN(new_n936));
  INV_X1    g0736(.A(new_n829), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n936), .A2(new_n870), .B1(new_n834), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n905), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT39), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n908), .B2(new_n916), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n903), .A2(KEYINPUT39), .A3(new_n904), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n665), .A2(new_n696), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n668), .A2(new_n894), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n939), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n935), .B(new_n947), .Z(new_n948));
  OAI22_X1  g0748(.A1(new_n933), .A2(new_n948), .B1(new_n206), .B2(new_n767), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n948), .B2(new_n933), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n532), .A2(new_n536), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT35), .ZN(new_n952));
  OAI211_X1 g0752(.A(G116), .B(new_n214), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n952), .B2(new_n951), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT36), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n217), .A2(new_n225), .A3(new_n324), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n206), .B(G13), .C1(new_n956), .C2(new_n245), .ZN(new_n957));
  OR3_X1    g0757(.A1(new_n950), .A2(new_n955), .A3(new_n957), .ZN(G367));
  NOR2_X1   g0758(.A1(new_n562), .A2(new_n695), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n711), .B1(new_n705), .B2(new_n704), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n751), .A2(new_n695), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n576), .A2(new_n562), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n696), .B1(new_n563), .B2(new_n573), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n960), .A2(new_n713), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n959), .B1(new_n965), .B2(KEYINPUT42), .ZN(new_n966));
  INV_X1    g0766(.A(new_n964), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n707), .A2(KEYINPUT42), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n714), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT109), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n966), .A2(KEYINPUT109), .A3(new_n969), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n619), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n596), .A2(new_n696), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(new_n679), .ZN(new_n978));
  OR3_X1    g0778(.A1(new_n977), .A2(new_n978), .A3(KEYINPUT106), .ZN(new_n979));
  OAI21_X1  g0779(.A(KEYINPUT106), .B1(new_n977), .B2(new_n978), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n981), .B(KEYINPUT107), .ZN(new_n984));
  XNOR2_X1  g0784(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n974), .A2(new_n983), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n988), .B1(new_n974), .B2(new_n983), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n989), .A2(new_n709), .A3(new_n964), .A4(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n989), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n993), .A2(new_n990), .B1(new_n710), .B2(new_n967), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n717), .B(KEYINPUT41), .Z(new_n995));
  OAI21_X1  g0795(.A(new_n708), .B1(new_n712), .B2(new_n695), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n960), .A2(new_n713), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(new_n703), .Z(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n765), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n714), .A2(new_n964), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT45), .Z(new_n1003));
  NOR2_X1   g0803(.A1(new_n714), .A2(new_n964), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT44), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1003), .A2(new_n710), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n709), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1001), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n995), .B1(new_n1009), .B2(new_n765), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n992), .B(new_n994), .C1(new_n1010), .C2(new_n769), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n779), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n236), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n787), .B1(new_n210), .B2(new_n400), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n770), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n818), .A2(new_n852), .B1(new_n808), .B2(new_n202), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n303), .B(new_n1016), .C1(G137), .C2(new_n804), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n823), .A2(G68), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n800), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n811), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G143), .A2(new_n1019), .B1(new_n1020), .B2(G77), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G159), .A2(new_n791), .B1(new_n795), .B2(G58), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1017), .A2(new_n1018), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n846), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G303), .A2(new_n802), .B1(new_n807), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(G317), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1025), .B1(new_n1026), .B2(new_n842), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n472), .A2(new_n790), .B1(new_n800), .B2(new_n806), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n588), .B2(new_n1020), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n795), .A2(G116), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT46), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n332), .B1(new_n858), .B2(G107), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1028), .A2(new_n1030), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1023), .A2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT47), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1015), .B1(new_n1036), .B2(new_n786), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n776), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1037), .B1(new_n982), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1011), .A2(new_n1039), .ZN(G387));
  NAND2_X1  g0840(.A1(new_n999), .A2(new_n769), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n787), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n779), .B1(new_n240), .B2(new_n781), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n210), .A2(new_n294), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1043), .B1(new_n719), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n263), .ZN(new_n1046));
  OR3_X1    g0846(.A1(new_n1046), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1047));
  AOI21_X1  g0847(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT50), .B1(new_n1046), .B2(G50), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1047), .A2(new_n719), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1045), .A2(new_n1050), .B1(new_n227), .B2(new_n716), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G303), .A2(new_n807), .B1(new_n802), .B2(G317), .ZN(new_n1052));
  INV_X1    g0852(.A(G322), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1052), .B1(new_n806), .B2(new_n790), .C1(new_n1053), .C2(new_n800), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT48), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n858), .A2(new_n1024), .B1(new_n795), .B2(G294), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT112), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1060), .A2(KEYINPUT49), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n334), .B1(new_n623), .B2(new_n811), .C1(new_n842), .C2(new_n799), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n1060), .B2(KEYINPUT49), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n823), .A2(new_n401), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n202), .B2(new_n818), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT111), .Z(new_n1066));
  INV_X1    g0866(.A(G159), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n808), .A2(new_n219), .B1(new_n1067), .B2(new_n800), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n334), .B1(G150), .B2(new_n804), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n225), .B2(new_n794), .C1(new_n812), .C2(new_n528), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT110), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1068), .B(new_n1071), .C1(new_n263), .C2(new_n791), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1061), .A2(new_n1063), .B1(new_n1066), .B2(new_n1072), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n770), .B1(new_n1042), .B2(new_n1051), .C1(new_n1073), .C2(new_n826), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n708), .B2(new_n776), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT113), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1000), .A2(new_n717), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n999), .A2(new_n765), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1041), .B(new_n1076), .C1(new_n1077), .C2(new_n1078), .ZN(G393));
  AND2_X1   g0879(.A1(new_n1008), .A2(new_n1006), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n769), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1012), .A2(new_n244), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n787), .B1(new_n210), .B2(new_n621), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n770), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1019), .A2(G317), .B1(new_n802), .B2(G311), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT52), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G116), .A2(new_n858), .B1(new_n795), .B2(new_n1024), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n637), .B2(new_n790), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n303), .B1(new_n842), .B2(new_n1053), .C1(new_n472), .C2(new_n808), .ZN(new_n1089));
  NOR4_X1   g0889(.A1(new_n1086), .A2(new_n1088), .A3(new_n822), .A4(new_n1089), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1090), .A2(KEYINPUT114), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(KEYINPUT114), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n263), .A2(new_n807), .B1(new_n804), .B2(G143), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G50), .A2(new_n791), .B1(new_n795), .B2(G68), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n845), .A2(new_n332), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n823), .A2(G77), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1019), .A2(G150), .B1(new_n802), .B2(G159), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1097), .A2(KEYINPUT51), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(KEYINPUT51), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1096), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1091), .B(new_n1092), .C1(new_n1095), .C2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1084), .B1(new_n1101), .B2(new_n786), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n964), .B2(new_n1038), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1009), .A2(new_n717), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1080), .A2(new_n1001), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1081), .B(new_n1103), .C1(new_n1104), .C2(new_n1105), .ZN(G390));
  NAND4_X1  g0906(.A1(new_n883), .A2(G330), .A3(new_n831), .A4(new_n885), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n876), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n830), .A2(new_n408), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n763), .A2(new_n696), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n876), .A2(new_n740), .A3(new_n831), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1109), .A2(new_n937), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(G330), .B(new_n831), .C1(new_n877), .C2(new_n882), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(new_n936), .A3(new_n870), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n883), .A2(G330), .A3(new_n885), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n927), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n834), .A2(new_n937), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n1117), .A2(KEYINPUT115), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(KEYINPUT115), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1113), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n934), .B(new_n671), .C1(new_n469), .C2(new_n1116), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n941), .A2(new_n942), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n938), .B2(new_n944), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1108), .B1(new_n1111), .B2(new_n937), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n917), .A2(new_n920), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n943), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1126), .B(new_n1112), .C1(new_n1127), .C2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1118), .A2(new_n876), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1131), .A2(new_n943), .B1(new_n941), .B2(new_n942), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1111), .A2(new_n937), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n876), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1129), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1132), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1116), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n928), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1130), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n718), .B1(new_n1124), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1126), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1141), .A2(new_n928), .A3(new_n1137), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1121), .A2(new_n1142), .A3(new_n1130), .A4(new_n1123), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1139), .A2(new_n768), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1125), .A2(new_n774), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n623), .A2(new_n818), .B1(new_n808), .B2(new_n621), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n294), .B(new_n1147), .C1(G294), .C2(new_n804), .ZN(new_n1148));
  INV_X1    g0948(.A(G283), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n800), .A2(new_n1149), .B1(new_n794), .B2(new_n221), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G107), .B2(new_n791), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1148), .A2(new_n856), .A3(new_n1096), .A4(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n804), .A2(G125), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1153), .B1(new_n808), .B2(new_n1154), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n303), .B(new_n1155), .C1(G132), .C2(new_n802), .ZN(new_n1156));
  INV_X1    g0956(.A(G128), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n1157), .A2(new_n800), .B1(new_n790), .B2(new_n851), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G50), .B2(new_n1020), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n794), .A2(new_n852), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT53), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n823), .A2(G159), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1156), .A2(new_n1159), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n826), .B1(new_n1152), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n839), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n770), .B1(new_n1165), .B2(new_n263), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1166), .B(KEYINPUT116), .Z(new_n1167));
  NOR2_X1   g0967(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1146), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1145), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1144), .A2(new_n1171), .ZN(G378));
  NAND2_X1  g0972(.A1(new_n270), .A2(new_n894), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n320), .B(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1174), .B(new_n1175), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n924), .A2(new_n831), .A3(new_n905), .A4(new_n876), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n883), .A2(new_n885), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n927), .A2(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1177), .A2(new_n866), .B1(new_n1179), .B2(new_n921), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1176), .B1(new_n1180), .B2(G330), .ZN(new_n1181));
  AND4_X1   g0981(.A1(G330), .A2(new_n907), .A3(new_n929), .A4(new_n1176), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n947), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1176), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n930), .B2(new_n702), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n947), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1180), .A2(G330), .A3(new_n1176), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1183), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1113), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT115), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1117), .A2(KEYINPUT115), .A3(new_n1118), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1190), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1123), .B1(new_n1139), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1189), .A2(new_n1196), .A3(KEYINPUT57), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1143), .A2(new_n1123), .B1(new_n1183), .B2(new_n1188), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(new_n717), .C1(new_n1198), .C2(KEYINPUT57), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1189), .A2(new_n769), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n771), .B1(new_n839), .B2(new_n202), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n794), .A2(new_n1154), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1202), .A2(KEYINPUT117), .B1(G128), .B2(new_n802), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(KEYINPUT117), .B2(new_n1202), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT118), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1019), .A2(G125), .B1(new_n807), .B2(G137), .ZN(new_n1206));
  INV_X1    g1006(.A(G132), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1206), .B1(new_n1207), .B2(new_n790), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G150), .B2(new_n823), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1205), .A2(new_n1209), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT59), .Z(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1212), .A2(KEYINPUT119), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(KEYINPUT119), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1020), .A2(G159), .ZN(new_n1215));
  AOI211_X1 g1015(.A(G33), .B(G41), .C1(new_n804), .C2(G124), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G107), .A2(new_n802), .B1(new_n807), .B2(new_n401), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n1149), .B2(new_n842), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n811), .A2(new_n323), .B1(new_n794), .B2(new_n225), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n528), .A2(new_n790), .B1(new_n800), .B2(new_n623), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n332), .A2(G41), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NOR4_X1   g1023(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .A4(new_n1223), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1224), .A2(new_n1018), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(KEYINPUT58), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1223), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1225), .A2(KEYINPUT58), .ZN(new_n1228));
  AND4_X1   g1028(.A1(new_n1217), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1201), .B1(new_n826), .B2(new_n1229), .C1(new_n1176), .C2(new_n775), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1200), .A2(new_n1230), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1199), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(G375));
  OAI21_X1  g1033(.A(KEYINPUT120), .B1(new_n1195), .B2(new_n768), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1108), .A2(new_n774), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT121), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n818), .A2(new_n1149), .B1(new_n808), .B2(new_n227), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n294), .B(new_n1237), .C1(G303), .C2(new_n804), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n790), .A2(new_n623), .B1(new_n794), .B2(new_n528), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G294), .B2(new_n1019), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n813), .A2(G77), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1238), .A2(new_n1064), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n808), .A2(new_n852), .B1(new_n842), .B2(new_n1157), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G137), .B2(new_n802), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n823), .A2(G50), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n800), .A2(new_n1207), .B1(new_n794), .B2(new_n1067), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1154), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1246), .B1(new_n791), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n334), .B1(new_n1020), .B2(G58), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1244), .A2(new_n1245), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n826), .B1(new_n1242), .B2(new_n1250), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n771), .B(new_n1251), .C1(new_n219), .C2(new_n839), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1236), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1234), .A2(new_n1253), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1195), .A2(KEYINPUT120), .A3(new_n768), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n995), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1122), .B(new_n1113), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1124), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1256), .A2(new_n1259), .ZN(G381));
  OR2_X1    g1060(.A1(G393), .A2(G396), .ZN(new_n1261));
  OR3_X1    g1061(.A1(G390), .A2(new_n1261), .A3(G384), .ZN(new_n1262));
  NOR4_X1   g1062(.A1(new_n1262), .A2(G387), .A3(G378), .A4(G381), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1232), .ZN(G407));
  AOI211_X1 g1064(.A(new_n1145), .B(new_n1170), .C1(new_n1140), .C2(new_n1143), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n694), .A2(G213), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1232), .A2(new_n1265), .A3(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(G407), .A2(G213), .A3(new_n1268), .ZN(G409));
  NAND3_X1  g1069(.A1(new_n1199), .A2(G378), .A3(new_n1231), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1189), .A2(new_n1196), .A3(new_n1257), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1200), .A2(new_n1230), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1265), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1267), .B1(new_n1270), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT123), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT122), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT60), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1278), .B1(new_n1258), .B2(new_n1279), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1195), .A2(KEYINPUT122), .A3(KEYINPUT60), .A4(new_n1122), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1258), .A2(new_n1279), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n718), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G384), .B1(new_n1285), .B2(new_n1256), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1256), .A3(G384), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1267), .A2(G2897), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1289), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1276), .B(new_n1277), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1285), .A2(new_n1256), .A3(G384), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1294), .A2(new_n1286), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1293), .A2(new_n1266), .A3(new_n1295), .ZN(new_n1296));
  OR2_X1    g1096(.A1(new_n1296), .A2(KEYINPUT63), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(KEYINPUT63), .ZN(new_n1298));
  INV_X1    g1098(.A(G390), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G393), .A2(G396), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1261), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(G390), .A2(new_n1261), .A3(new_n1300), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT124), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1011), .A2(new_n1305), .A3(new_n1039), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1305), .B1(new_n1011), .B2(new_n1039), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1304), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1308), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1310), .A2(new_n1306), .A3(new_n1303), .A4(new_n1302), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1309), .A2(new_n1311), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1312), .A2(KEYINPUT61), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1292), .A2(new_n1297), .A3(new_n1298), .A4(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT61), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1315), .B1(new_n1316), .B2(new_n1274), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1318), .B1(new_n1274), .B2(new_n1295), .ZN(new_n1319));
  AOI22_X1  g1119(.A1(KEYINPUT126), .A2(new_n1319), .B1(new_n1296), .B2(KEYINPUT62), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT126), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1321), .B1(new_n1296), .B2(new_n1318), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1317), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1309), .A2(new_n1311), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1314), .B1(new_n1323), .B2(new_n1324), .ZN(G405));
  INV_X1    g1125(.A(new_n1295), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(KEYINPUT127), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1324), .A2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1312), .A2(KEYINPUT127), .A3(new_n1326), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1270), .B1(new_n1326), .B2(KEYINPUT127), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1331), .B1(new_n1265), .B2(G375), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1330), .B(new_n1332), .ZN(G402));
endmodule


