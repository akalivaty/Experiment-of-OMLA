

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763;

  INV_X1 U375 ( .A(n719), .ZN(n395) );
  NAND2_X1 U376 ( .A1(n377), .A2(n373), .ZN(n565) );
  NAND2_X1 U377 ( .A1(n726), .A2(n395), .ZN(n394) );
  XNOR2_X1 U378 ( .A(n367), .B(KEYINPUT97), .ZN(n528) );
  AND2_X1 U379 ( .A1(n528), .A2(KEYINPUT66), .ZN(n527) );
  XNOR2_X1 U380 ( .A(n368), .B(n391), .ZN(n401) );
  OR2_X1 U381 ( .A1(n396), .A2(n572), .ZN(n597) );
  NOR2_X2 U382 ( .A1(n597), .A2(n563), .ZN(n718) );
  OR2_X1 U383 ( .A1(n611), .A2(n612), .ZN(n353) );
  INV_X1 U384 ( .A(n636), .ZN(n518) );
  NAND2_X1 U385 ( .A1(n518), .A2(n634), .ZN(n533) );
  XNOR2_X2 U386 ( .A(n750), .B(n429), .ZN(n737) );
  AND2_X1 U387 ( .A1(n401), .A2(n618), .ZN(n620) );
  NAND2_X1 U388 ( .A1(n401), .A2(n617), .ZN(n749) );
  NOR2_X1 U389 ( .A1(n565), .A2(n605), .ZN(n404) );
  NAND2_X1 U390 ( .A1(n639), .A2(n568), .ZN(n585) );
  XNOR2_X1 U391 ( .A(n750), .B(n439), .ZN(n673) );
  XNOR2_X1 U392 ( .A(n487), .B(G134), .ZN(n469) );
  NOR2_X1 U393 ( .A1(n685), .A2(KEYINPUT44), .ZN(n525) );
  NAND2_X1 U394 ( .A1(n666), .A2(n665), .ZN(n367) );
  AND2_X1 U395 ( .A1(n371), .A2(n370), .ZN(n730) );
  NAND2_X1 U396 ( .A1(n577), .A2(n576), .ZN(n722) );
  NOR2_X1 U397 ( .A1(n593), .A2(n592), .ZN(n596) );
  XNOR2_X1 U398 ( .A(n404), .B(n567), .ZN(n403) );
  NOR2_X1 U399 ( .A1(n565), .A2(n585), .ZN(n561) );
  XNOR2_X1 U400 ( .A(n565), .B(n413), .ZN(n586) );
  XNOR2_X1 U401 ( .A(n499), .B(n498), .ZN(n570) );
  XNOR2_X1 U402 ( .A(n594), .B(KEYINPUT39), .ZN(n595) );
  NOR2_X1 U403 ( .A1(n611), .A2(n354), .ZN(n383) );
  OR2_X1 U404 ( .A1(n612), .A2(KEYINPUT87), .ZN(n354) );
  XNOR2_X1 U405 ( .A(n524), .B(KEYINPUT35), .ZN(n355) );
  XNOR2_X1 U406 ( .A(n524), .B(KEYINPUT35), .ZN(n685) );
  AND2_X2 U407 ( .A1(n668), .A2(n752), .ZN(n669) );
  XNOR2_X1 U408 ( .A(n601), .B(n361), .ZN(n393) );
  OR2_X2 U409 ( .A1(n570), .A2(n605), .ZN(n587) );
  XNOR2_X1 U410 ( .A(n469), .B(n416), .ZN(n420) );
  INV_X1 U411 ( .A(G137), .ZN(n416) );
  NOR2_X1 U412 ( .A1(n410), .A2(n726), .ZN(n603) );
  XNOR2_X1 U413 ( .A(n412), .B(n411), .ZN(n410) );
  INV_X1 U414 ( .A(KEYINPUT108), .ZN(n411) );
  NOR2_X1 U415 ( .A1(n586), .A2(n585), .ZN(n412) );
  XNOR2_X1 U416 ( .A(n580), .B(n579), .ZN(n581) );
  INV_X1 U417 ( .A(KEYINPUT48), .ZN(n391) );
  NOR2_X1 U418 ( .A1(G237), .A2(G953), .ZN(n432) );
  NOR2_X1 U419 ( .A1(n614), .A2(n613), .ZN(n615) );
  OR2_X1 U420 ( .A1(n673), .A2(n378), .ZN(n377) );
  AND2_X1 U421 ( .A1(n374), .A2(n376), .ZN(n373) );
  INV_X1 U422 ( .A(G110), .ZN(n421) );
  XNOR2_X1 U423 ( .A(n466), .B(n398), .ZN(n700) );
  XNOR2_X1 U424 ( .A(n400), .B(n399), .ZN(n398) );
  XNOR2_X1 U425 ( .A(n463), .B(G113), .ZN(n399) );
  INV_X1 U426 ( .A(KEYINPUT64), .ZN(n422) );
  NOR2_X1 U427 ( .A1(n615), .A2(n616), .ZN(n381) );
  XNOR2_X1 U428 ( .A(n598), .B(n362), .ZN(n656) );
  INV_X1 U429 ( .A(KEYINPUT41), .ZN(n362) );
  NAND2_X1 U430 ( .A1(n603), .A2(n588), .ZN(n372) );
  OR2_X1 U431 ( .A1(n737), .A2(n387), .ZN(n386) );
  AND2_X1 U432 ( .A1(n385), .A2(n389), .ZN(n388) );
  NAND2_X1 U433 ( .A1(n430), .A2(n440), .ZN(n387) );
  XNOR2_X1 U434 ( .A(n456), .B(n455), .ZN(n457) );
  NOR2_X1 U435 ( .A1(n624), .A2(n638), .ZN(n510) );
  XNOR2_X1 U436 ( .A(n394), .B(KEYINPUT106), .ZN(n625) );
  XNOR2_X1 U437 ( .A(KEYINPUT2), .B(KEYINPUT88), .ZN(n612) );
  XNOR2_X1 U438 ( .A(n607), .B(KEYINPUT38), .ZN(n622) );
  XNOR2_X1 U439 ( .A(n460), .B(n359), .ZN(n400) );
  XNOR2_X1 U440 ( .A(G146), .B(KEYINPUT74), .ZN(n417) );
  XOR2_X1 U441 ( .A(G131), .B(KEYINPUT75), .Z(n418) );
  XNOR2_X1 U442 ( .A(n497), .B(n496), .ZN(n498) );
  AND2_X1 U443 ( .A1(n569), .A2(n568), .ZN(n402) );
  NAND2_X1 U444 ( .A1(G469), .A2(G902), .ZN(n389) );
  XNOR2_X1 U445 ( .A(G116), .B(G113), .ZN(n435) );
  XNOR2_X1 U446 ( .A(G128), .B(G110), .ZN(n446) );
  XNOR2_X1 U447 ( .A(n447), .B(n364), .ZN(n448) );
  XNOR2_X1 U448 ( .A(G137), .B(KEYINPUT102), .ZN(n447) );
  XNOR2_X1 U449 ( .A(n365), .B(KEYINPUT23), .ZN(n364) );
  INV_X1 U450 ( .A(KEYINPUT24), .ZN(n365) );
  XOR2_X1 U451 ( .A(G116), .B(KEYINPUT7), .Z(n471) );
  XNOR2_X1 U452 ( .A(G107), .B(G122), .ZN(n470) );
  INV_X1 U453 ( .A(G128), .ZN(n414) );
  NAND2_X1 U454 ( .A1(n671), .A2(n670), .ZN(n408) );
  INV_X1 U455 ( .A(G953), .ZN(n503) );
  XNOR2_X1 U456 ( .A(n467), .B(n356), .ZN(n541) );
  INV_X1 U457 ( .A(KEYINPUT0), .ZN(n508) );
  INV_X1 U458 ( .A(KEYINPUT6), .ZN(n413) );
  BUF_X1 U459 ( .A(n733), .Z(n744) );
  XNOR2_X1 U460 ( .A(n428), .B(n427), .ZN(n429) );
  NAND2_X1 U461 ( .A1(n353), .A2(n381), .ZN(n380) );
  NAND2_X1 U462 ( .A1(n599), .A2(n656), .ZN(n600) );
  XNOR2_X1 U463 ( .A(n407), .B(n405), .ZN(n762) );
  XNOR2_X1 U464 ( .A(n406), .B(KEYINPUT40), .ZN(n405) );
  INV_X1 U465 ( .A(KEYINPUT111), .ZN(n406) );
  INV_X1 U466 ( .A(n589), .ZN(n370) );
  XNOR2_X1 U467 ( .A(n372), .B(n360), .ZN(n371) );
  INV_X1 U468 ( .A(n726), .ZN(n723) );
  INV_X1 U469 ( .A(KEYINPUT67), .ZN(n515) );
  INV_X1 U470 ( .A(G122), .ZN(n684) );
  NAND2_X1 U471 ( .A1(n441), .A2(G902), .ZN(n376) );
  OR2_X1 U472 ( .A1(G902), .A2(n700), .ZN(n356) );
  XOR2_X1 U473 ( .A(KEYINPUT8), .B(KEYINPUT72), .Z(n357) );
  XOR2_X1 U474 ( .A(G146), .B(G119), .Z(n358) );
  AND2_X1 U475 ( .A1(G214), .A2(n464), .ZN(n359) );
  INV_X1 U476 ( .A(G469), .ZN(n430) );
  NAND2_X2 U477 ( .A1(n388), .A2(n386), .ZN(n591) );
  XOR2_X1 U478 ( .A(KEYINPUT112), .B(KEYINPUT36), .Z(n360) );
  XOR2_X1 U479 ( .A(KEYINPUT94), .B(KEYINPUT46), .Z(n361) );
  INV_X2 U480 ( .A(G104), .ZN(n390) );
  NAND2_X1 U481 ( .A1(n363), .A2(n512), .ZN(n513) );
  INV_X1 U482 ( .A(n544), .ZN(n363) );
  XNOR2_X2 U483 ( .A(n511), .B(KEYINPUT22), .ZN(n544) );
  NOR2_X2 U484 ( .A1(G902), .A2(n745), .ZN(n458) );
  XNOR2_X1 U485 ( .A(n584), .B(n583), .ZN(n392) );
  INV_X1 U486 ( .A(n668), .ZN(n686) );
  XNOR2_X2 U487 ( .A(n554), .B(KEYINPUT45), .ZN(n668) );
  NOR2_X1 U488 ( .A1(n383), .A2(n366), .ZN(n382) );
  NAND2_X1 U489 ( .A1(n379), .A2(n671), .ZN(n366) );
  XNOR2_X1 U490 ( .A(n384), .B(KEYINPUT92), .ZN(n662) );
  XNOR2_X1 U491 ( .A(n516), .B(n515), .ZN(n517) );
  NAND2_X1 U492 ( .A1(n369), .A2(n392), .ZN(n368) );
  AND2_X1 U493 ( .A1(n590), .A2(n393), .ZN(n369) );
  NAND2_X1 U494 ( .A1(n673), .A2(n375), .ZN(n374) );
  NOR2_X1 U495 ( .A1(n441), .A2(G902), .ZN(n375) );
  INV_X1 U496 ( .A(n441), .ZN(n378) );
  NAND2_X1 U497 ( .A1(n615), .A2(n616), .ZN(n379) );
  NAND2_X1 U498 ( .A1(n382), .A2(n380), .ZN(n384) );
  NAND2_X1 U499 ( .A1(n737), .A2(G469), .ZN(n385) );
  XNOR2_X2 U500 ( .A(n591), .B(n431), .ZN(n636) );
  XNOR2_X1 U501 ( .A(n520), .B(n519), .ZN(n631) );
  XNOR2_X2 U502 ( .A(n390), .B(G122), .ZN(n480) );
  NAND2_X1 U503 ( .A1(n718), .A2(n625), .ZN(n564) );
  XNOR2_X1 U504 ( .A(n561), .B(n397), .ZN(n396) );
  INV_X1 U505 ( .A(KEYINPUT28), .ZN(n397) );
  NAND2_X1 U506 ( .A1(n403), .A2(n402), .ZN(n593) );
  NAND2_X1 U507 ( .A1(n763), .A2(n762), .ZN(n601) );
  NAND2_X1 U508 ( .A1(n602), .A2(n723), .ZN(n407) );
  NOR2_X4 U509 ( .A1(n408), .A2(n672), .ZN(n733) );
  NAND2_X1 U510 ( .A1(n409), .A2(n668), .ZN(n671) );
  XNOR2_X1 U511 ( .A(n620), .B(n619), .ZN(n409) );
  NOR2_X2 U512 ( .A1(n582), .A2(n581), .ZN(n584) );
  INV_X1 U513 ( .A(KEYINPUT89), .ZN(n579) );
  INV_X1 U514 ( .A(KEYINPUT79), .ZN(n583) );
  XNOR2_X1 U515 ( .A(n566), .B(KEYINPUT109), .ZN(n567) );
  BUF_X1 U516 ( .A(n631), .Z(n657) );
  INV_X1 U517 ( .A(n639), .ZN(n569) );
  XNOR2_X1 U518 ( .A(n471), .B(n470), .ZN(n472) );
  INV_X1 U519 ( .A(KEYINPUT76), .ZN(n594) );
  XNOR2_X1 U520 ( .A(KEYINPUT83), .B(KEYINPUT25), .ZN(n455) );
  XNOR2_X1 U521 ( .A(n473), .B(n472), .ZN(n474) );
  OR2_X1 U522 ( .A1(n753), .A2(G952), .ZN(n703) );
  XNOR2_X2 U523 ( .A(G143), .B(KEYINPUT65), .ZN(n415) );
  XNOR2_X2 U524 ( .A(n415), .B(n414), .ZN(n487) );
  XNOR2_X1 U525 ( .A(n418), .B(n417), .ZN(n465) );
  XNOR2_X1 U526 ( .A(KEYINPUT4), .B(n465), .ZN(n419) );
  XNOR2_X2 U527 ( .A(n420), .B(n419), .ZN(n750) );
  XNOR2_X1 U528 ( .A(n421), .B(G107), .ZN(n481) );
  XOR2_X1 U529 ( .A(n481), .B(KEYINPUT101), .Z(n424) );
  XNOR2_X2 U530 ( .A(n422), .B(G953), .ZN(n753) );
  NAND2_X1 U531 ( .A1(G227), .A2(n753), .ZN(n423) );
  XNOR2_X1 U532 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U533 ( .A(KEYINPUT84), .B(G140), .Z(n426) );
  XNOR2_X1 U534 ( .A(G104), .B(G101), .ZN(n425) );
  XNOR2_X1 U535 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U536 ( .A(KEYINPUT68), .B(KEYINPUT1), .Z(n431) );
  XNOR2_X1 U537 ( .A(n636), .B(KEYINPUT98), .ZN(n589) );
  XNOR2_X1 U538 ( .A(n432), .B(KEYINPUT82), .ZN(n464) );
  NAND2_X1 U539 ( .A1(n464), .A2(G210), .ZN(n434) );
  XOR2_X1 U540 ( .A(KEYINPUT81), .B(KEYINPUT5), .Z(n433) );
  XNOR2_X1 U541 ( .A(n434), .B(n433), .ZN(n438) );
  XNOR2_X1 U542 ( .A(n435), .B(G119), .ZN(n437) );
  XNOR2_X1 U543 ( .A(G101), .B(KEYINPUT3), .ZN(n436) );
  XNOR2_X1 U544 ( .A(n437), .B(n436), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n438), .B(n483), .ZN(n439) );
  INV_X1 U546 ( .A(G902), .ZN(n440) );
  XNOR2_X1 U547 ( .A(KEYINPUT77), .B(G472), .ZN(n441) );
  XOR2_X1 U548 ( .A(G140), .B(KEYINPUT10), .Z(n443) );
  XNOR2_X1 U549 ( .A(G125), .B(KEYINPUT73), .ZN(n442) );
  XNOR2_X1 U550 ( .A(n443), .B(n442), .ZN(n751) );
  NAND2_X1 U551 ( .A1(G234), .A2(n753), .ZN(n445) );
  XNOR2_X1 U552 ( .A(n357), .B(KEYINPUT90), .ZN(n444) );
  XNOR2_X1 U553 ( .A(n445), .B(n444), .ZN(n468) );
  NAND2_X1 U554 ( .A1(G221), .A2(n468), .ZN(n451) );
  XNOR2_X1 U555 ( .A(n358), .B(n446), .ZN(n449) );
  XOR2_X1 U556 ( .A(n449), .B(n448), .Z(n450) );
  XNOR2_X1 U557 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U558 ( .A(n751), .B(n452), .Z(n745) );
  XOR2_X1 U559 ( .A(KEYINPUT103), .B(KEYINPUT20), .Z(n454) );
  XNOR2_X1 U560 ( .A(KEYINPUT15), .B(G902), .ZN(n493) );
  NAND2_X1 U561 ( .A1(G234), .A2(n493), .ZN(n453) );
  XNOR2_X1 U562 ( .A(n454), .B(n453), .ZN(n477) );
  NAND2_X1 U563 ( .A1(n477), .A2(G217), .ZN(n456) );
  XNOR2_X2 U564 ( .A(n458), .B(n457), .ZN(n639) );
  NAND2_X1 U565 ( .A1(n586), .A2(n639), .ZN(n459) );
  NOR2_X1 U566 ( .A1(n589), .A2(n459), .ZN(n512) );
  XNOR2_X1 U567 ( .A(KEYINPUT13), .B(G475), .ZN(n467) );
  XNOR2_X1 U568 ( .A(n480), .B(G143), .ZN(n460) );
  XOR2_X1 U569 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n462) );
  XNOR2_X1 U570 ( .A(KEYINPUT105), .B(KEYINPUT104), .ZN(n461) );
  XNOR2_X1 U571 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U572 ( .A(n465), .B(n751), .Z(n466) );
  NAND2_X1 U573 ( .A1(n468), .A2(G217), .ZN(n475) );
  XOR2_X1 U574 ( .A(KEYINPUT9), .B(n469), .Z(n473) );
  XNOR2_X1 U575 ( .A(n475), .B(n474), .ZN(n741) );
  NOR2_X1 U576 ( .A1(G902), .A2(n741), .ZN(n476) );
  XNOR2_X1 U577 ( .A(G478), .B(n476), .ZN(n539) );
  NAND2_X1 U578 ( .A1(n541), .A2(n539), .ZN(n624) );
  NAND2_X1 U579 ( .A1(G221), .A2(n477), .ZN(n478) );
  XNOR2_X1 U580 ( .A(n478), .B(KEYINPUT21), .ZN(n638) );
  XNOR2_X1 U581 ( .A(KEYINPUT78), .B(KEYINPUT16), .ZN(n479) );
  XNOR2_X1 U582 ( .A(n480), .B(n479), .ZN(n482) );
  XNOR2_X1 U583 ( .A(n482), .B(n481), .ZN(n484) );
  XNOR2_X1 U584 ( .A(n484), .B(n483), .ZN(n694) );
  XNOR2_X1 U585 ( .A(G146), .B(G125), .ZN(n485) );
  XNOR2_X1 U586 ( .A(n485), .B(KEYINPUT4), .ZN(n486) );
  XNOR2_X1 U587 ( .A(n487), .B(n486), .ZN(n491) );
  NAND2_X1 U588 ( .A1(n753), .A2(G224), .ZN(n489) );
  XNOR2_X1 U589 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n488) );
  XNOR2_X1 U590 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U591 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U592 ( .A(n694), .B(n492), .ZN(n679) );
  INV_X1 U593 ( .A(n493), .ZN(n670) );
  OR2_X2 U594 ( .A1(n679), .A2(n670), .ZN(n499) );
  NOR2_X1 U595 ( .A1(G902), .A2(G237), .ZN(n494) );
  XNOR2_X1 U596 ( .A(n494), .B(KEYINPUT80), .ZN(n501) );
  INV_X1 U597 ( .A(G210), .ZN(n495) );
  OR2_X1 U598 ( .A1(n501), .A2(n495), .ZN(n497) );
  INV_X1 U599 ( .A(KEYINPUT85), .ZN(n496) );
  INV_X1 U600 ( .A(G214), .ZN(n500) );
  OR2_X1 U601 ( .A1(n501), .A2(n500), .ZN(n502) );
  XNOR2_X1 U602 ( .A(n502), .B(KEYINPUT100), .ZN(n621) );
  INV_X1 U603 ( .A(n621), .ZN(n605) );
  XNOR2_X2 U604 ( .A(n587), .B(KEYINPUT19), .ZN(n562) );
  NAND2_X1 U605 ( .A1(G952), .A2(n503), .ZN(n557) );
  NOR2_X1 U606 ( .A1(G898), .A2(n503), .ZN(n695) );
  NAND2_X1 U607 ( .A1(n695), .A2(G902), .ZN(n504) );
  NAND2_X1 U608 ( .A1(n557), .A2(n504), .ZN(n506) );
  NAND2_X1 U609 ( .A1(G234), .A2(G237), .ZN(n505) );
  XNOR2_X1 U610 ( .A(n505), .B(KEYINPUT14), .ZN(n652) );
  AND2_X1 U611 ( .A1(n506), .A2(n652), .ZN(n507) );
  NAND2_X1 U612 ( .A1(n562), .A2(n507), .ZN(n509) );
  XNOR2_X2 U613 ( .A(n509), .B(n508), .ZN(n538) );
  NAND2_X1 U614 ( .A1(n510), .A2(n538), .ZN(n511) );
  XNOR2_X1 U615 ( .A(n513), .B(KEYINPUT32), .ZN(n665) );
  NAND2_X1 U616 ( .A1(n565), .A2(n636), .ZN(n514) );
  NOR2_X2 U617 ( .A1(n544), .A2(n514), .ZN(n516) );
  NAND2_X1 U618 ( .A1(n517), .A2(n639), .ZN(n666) );
  NOR2_X1 U619 ( .A1(n638), .A2(n639), .ZN(n634) );
  NOR2_X1 U620 ( .A1(n533), .A2(n586), .ZN(n520) );
  XNOR2_X1 U621 ( .A(KEYINPUT107), .B(KEYINPUT33), .ZN(n519) );
  NAND2_X1 U622 ( .A1(n631), .A2(n538), .ZN(n522) );
  INV_X1 U623 ( .A(KEYINPUT34), .ZN(n521) );
  XNOR2_X1 U624 ( .A(n522), .B(n521), .ZN(n523) );
  NOR2_X1 U625 ( .A1(n541), .A2(n539), .ZN(n576) );
  NAND2_X1 U626 ( .A1(n523), .A2(n576), .ZN(n524) );
  XNOR2_X1 U627 ( .A(n525), .B(KEYINPUT71), .ZN(n526) );
  NAND2_X1 U628 ( .A1(n527), .A2(n526), .ZN(n532) );
  INV_X1 U629 ( .A(n528), .ZN(n530) );
  NAND2_X1 U630 ( .A1(KEYINPUT66), .A2(KEYINPUT44), .ZN(n529) );
  NAND2_X1 U631 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U632 ( .A1(n532), .A2(n531), .ZN(n553) );
  NAND2_X1 U633 ( .A1(n355), .A2(KEYINPUT44), .ZN(n548) );
  OR2_X1 U634 ( .A1(n533), .A2(n565), .ZN(n633) );
  INV_X1 U635 ( .A(n538), .ZN(n534) );
  NOR2_X1 U636 ( .A1(n633), .A2(n534), .ZN(n535) );
  XNOR2_X1 U637 ( .A(n535), .B(KEYINPUT31), .ZN(n728) );
  INV_X1 U638 ( .A(n565), .ZN(n644) );
  NAND2_X1 U639 ( .A1(n591), .A2(n634), .ZN(n536) );
  NOR2_X1 U640 ( .A1(n644), .A2(n536), .ZN(n537) );
  NAND2_X1 U641 ( .A1(n538), .A2(n537), .ZN(n713) );
  NAND2_X1 U642 ( .A1(n728), .A2(n713), .ZN(n542) );
  INV_X1 U643 ( .A(n539), .ZN(n540) );
  OR2_X1 U644 ( .A1(n541), .A2(n540), .ZN(n726) );
  AND2_X1 U645 ( .A1(n541), .A2(n540), .ZN(n719) );
  AND2_X1 U646 ( .A1(n542), .A2(n625), .ZN(n546) );
  NOR2_X1 U647 ( .A1(n518), .A2(n639), .ZN(n543) );
  NAND2_X1 U648 ( .A1(n543), .A2(n586), .ZN(n545) );
  NOR2_X1 U649 ( .A1(n545), .A2(n544), .ZN(n707) );
  NOR2_X1 U650 ( .A1(n546), .A2(n707), .ZN(n547) );
  NAND2_X1 U651 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U652 ( .A(n549), .B(KEYINPUT96), .ZN(n551) );
  NOR2_X1 U653 ( .A1(KEYINPUT44), .A2(KEYINPUT66), .ZN(n550) );
  NOR2_X1 U654 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U655 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U656 ( .A1(n668), .A2(KEYINPUT91), .ZN(n610) );
  NOR2_X1 U657 ( .A1(n753), .A2(G900), .ZN(n555) );
  NAND2_X1 U658 ( .A1(G902), .A2(n555), .ZN(n556) );
  NAND2_X1 U659 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U660 ( .A1(n652), .A2(n558), .ZN(n559) );
  XNOR2_X1 U661 ( .A(KEYINPUT86), .B(n559), .ZN(n560) );
  NOR2_X1 U662 ( .A1(n638), .A2(n560), .ZN(n568) );
  INV_X1 U663 ( .A(n562), .ZN(n563) );
  NOR2_X1 U664 ( .A1(KEYINPUT47), .A2(n564), .ZN(n582) );
  NAND2_X1 U665 ( .A1(n564), .A2(KEYINPUT47), .ZN(n578) );
  INV_X1 U666 ( .A(KEYINPUT30), .ZN(n566) );
  INV_X1 U667 ( .A(n593), .ZN(n574) );
  INV_X1 U668 ( .A(n591), .ZN(n572) );
  INV_X1 U669 ( .A(n570), .ZN(n571) );
  INV_X1 U670 ( .A(n571), .ZN(n607) );
  NOR2_X1 U671 ( .A1(n572), .A2(n607), .ZN(n573) );
  NAND2_X1 U672 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U673 ( .A(KEYINPUT110), .B(n575), .Z(n577) );
  NAND2_X1 U674 ( .A1(n578), .A2(n722), .ZN(n580) );
  INV_X1 U675 ( .A(n587), .ZN(n588) );
  XNOR2_X1 U676 ( .A(KEYINPUT95), .B(n730), .ZN(n590) );
  NAND2_X1 U677 ( .A1(n591), .A2(n622), .ZN(n592) );
  XNOR2_X1 U678 ( .A(n596), .B(n595), .ZN(n602) );
  INV_X1 U679 ( .A(n597), .ZN(n599) );
  NAND2_X1 U680 ( .A1(n622), .A2(n621), .ZN(n627) );
  NOR2_X1 U681 ( .A1(n627), .A2(n624), .ZN(n598) );
  XNOR2_X1 U682 ( .A(n600), .B(KEYINPUT42), .ZN(n763) );
  NAND2_X1 U683 ( .A1(n719), .A2(n602), .ZN(n732) );
  INV_X1 U684 ( .A(n732), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n603), .A2(n636), .ZN(n604) );
  NOR2_X1 U686 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U687 ( .A(n606), .B(KEYINPUT43), .ZN(n608) );
  NOR2_X1 U688 ( .A1(n608), .A2(n571), .ZN(n667) );
  NOR2_X1 U689 ( .A1(n609), .A2(n667), .ZN(n617) );
  NOR2_X1 U690 ( .A1(n610), .A2(n749), .ZN(n611) );
  NOR2_X1 U691 ( .A1(n668), .A2(n612), .ZN(n614) );
  INV_X1 U692 ( .A(KEYINPUT91), .ZN(n613) );
  INV_X1 U693 ( .A(KEYINPUT87), .ZN(n616) );
  AND2_X1 U694 ( .A1(KEYINPUT2), .A2(n617), .ZN(n618) );
  INV_X1 U695 ( .A(KEYINPUT93), .ZN(n619) );
  NOR2_X1 U696 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n629) );
  INV_X1 U698 ( .A(n625), .ZN(n626) );
  NOR2_X1 U699 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U701 ( .A(n630), .B(KEYINPUT119), .ZN(n632) );
  NAND2_X1 U702 ( .A1(n632), .A2(n657), .ZN(n650) );
  INV_X1 U703 ( .A(n633), .ZN(n646) );
  INV_X1 U704 ( .A(n634), .ZN(n635) );
  NAND2_X1 U705 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U706 ( .A(n637), .B(KEYINPUT50), .ZN(n642) );
  AND2_X1 U707 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U708 ( .A(n640), .B(KEYINPUT49), .ZN(n641) );
  NAND2_X1 U709 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U710 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U711 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U712 ( .A(KEYINPUT51), .B(n647), .ZN(n648) );
  NAND2_X1 U713 ( .A1(n648), .A2(n656), .ZN(n649) );
  NAND2_X1 U714 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U715 ( .A(KEYINPUT52), .B(n651), .Z(n654) );
  NAND2_X1 U716 ( .A1(n652), .A2(G952), .ZN(n653) );
  NOR2_X1 U717 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U718 ( .A(n655), .B(KEYINPUT120), .ZN(n660) );
  NAND2_X1 U719 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U720 ( .A1(n658), .A2(n503), .ZN(n659) );
  NOR2_X1 U721 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U722 ( .A1(n662), .A2(n661), .ZN(n664) );
  INV_X1 U723 ( .A(KEYINPUT53), .ZN(n663) );
  XNOR2_X1 U724 ( .A(n664), .B(n663), .ZN(G75) );
  XNOR2_X1 U725 ( .A(n665), .B(G119), .ZN(G21) );
  XNOR2_X1 U726 ( .A(n666), .B(G110), .ZN(G12) );
  XOR2_X1 U727 ( .A(G140), .B(n667), .Z(G42) );
  NOR2_X1 U728 ( .A1(n669), .A2(KEYINPUT2), .ZN(n672) );
  NAND2_X1 U729 ( .A1(n733), .A2(G472), .ZN(n675) );
  XNOR2_X1 U730 ( .A(n673), .B(KEYINPUT62), .ZN(n674) );
  XNOR2_X1 U731 ( .A(n675), .B(n674), .ZN(n676) );
  NAND2_X1 U732 ( .A1(n676), .A2(n703), .ZN(n677) );
  XNOR2_X1 U733 ( .A(n677), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U734 ( .A1(n733), .A2(G210), .ZN(n681) );
  XOR2_X1 U735 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n678) );
  XNOR2_X1 U736 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U737 ( .A(n681), .B(n680), .ZN(n682) );
  INV_X1 U738 ( .A(n703), .ZN(n748) );
  NOR2_X2 U739 ( .A1(n682), .A2(n748), .ZN(n683) );
  XNOR2_X1 U740 ( .A(n683), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U741 ( .A(n355), .B(n684), .ZN(G24) );
  NOR2_X1 U742 ( .A1(n686), .A2(G953), .ZN(n687) );
  XNOR2_X1 U743 ( .A(n687), .B(KEYINPUT125), .ZN(n693) );
  XOR2_X1 U744 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n689) );
  NAND2_X1 U745 ( .A1(G224), .A2(G953), .ZN(n688) );
  XNOR2_X1 U746 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U747 ( .A(KEYINPUT123), .B(n690), .ZN(n691) );
  NAND2_X1 U748 ( .A1(n691), .A2(G898), .ZN(n692) );
  NAND2_X1 U749 ( .A1(n693), .A2(n692), .ZN(n697) );
  NOR2_X1 U750 ( .A1(n694), .A2(n695), .ZN(n696) );
  XNOR2_X1 U751 ( .A(n697), .B(n696), .ZN(G69) );
  NAND2_X1 U752 ( .A1(n733), .A2(G475), .ZN(n702) );
  XNOR2_X1 U753 ( .A(KEYINPUT69), .B(KEYINPUT99), .ZN(n698) );
  XNOR2_X1 U754 ( .A(n698), .B(KEYINPUT59), .ZN(n699) );
  XNOR2_X1 U755 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U756 ( .A(n702), .B(n701), .ZN(n704) );
  NAND2_X1 U757 ( .A1(n704), .A2(n703), .ZN(n706) );
  XOR2_X1 U758 ( .A(KEYINPUT70), .B(KEYINPUT60), .Z(n705) );
  XNOR2_X1 U759 ( .A(n706), .B(n705), .ZN(G60) );
  XNOR2_X1 U760 ( .A(n707), .B(G101), .ZN(n708) );
  XNOR2_X1 U761 ( .A(n708), .B(KEYINPUT113), .ZN(G3) );
  NOR2_X1 U762 ( .A1(n713), .A2(n726), .ZN(n709) );
  XOR2_X1 U763 ( .A(KEYINPUT114), .B(n709), .Z(n710) );
  XNOR2_X1 U764 ( .A(G104), .B(n710), .ZN(G6) );
  XOR2_X1 U765 ( .A(KEYINPUT117), .B(KEYINPUT27), .Z(n712) );
  XNOR2_X1 U766 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n711) );
  XNOR2_X1 U767 ( .A(n712), .B(n711), .ZN(n717) );
  NOR2_X1 U768 ( .A1(n713), .A2(n395), .ZN(n715) );
  XNOR2_X1 U769 ( .A(G107), .B(KEYINPUT26), .ZN(n714) );
  XNOR2_X1 U770 ( .A(n715), .B(n714), .ZN(n716) );
  XOR2_X1 U771 ( .A(n717), .B(n716), .Z(G9) );
  XOR2_X1 U772 ( .A(G128), .B(KEYINPUT29), .Z(n721) );
  NAND2_X1 U773 ( .A1(n718), .A2(n719), .ZN(n720) );
  XNOR2_X1 U774 ( .A(n721), .B(n720), .ZN(G30) );
  XNOR2_X1 U775 ( .A(G143), .B(n722), .ZN(G45) );
  NAND2_X1 U776 ( .A1(n718), .A2(n723), .ZN(n724) );
  XNOR2_X1 U777 ( .A(n724), .B(KEYINPUT118), .ZN(n725) );
  XNOR2_X1 U778 ( .A(G146), .B(n725), .ZN(G48) );
  NOR2_X1 U779 ( .A1(n726), .A2(n728), .ZN(n727) );
  XOR2_X1 U780 ( .A(G113), .B(n727), .Z(G15) );
  NOR2_X1 U781 ( .A1(n395), .A2(n728), .ZN(n729) );
  XOR2_X1 U782 ( .A(G116), .B(n729), .Z(G18) );
  XNOR2_X1 U783 ( .A(G125), .B(n730), .ZN(n731) );
  XNOR2_X1 U784 ( .A(n731), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U785 ( .A(G134), .B(n732), .ZN(G36) );
  NAND2_X1 U786 ( .A1(n744), .A2(G469), .ZN(n739) );
  XOR2_X1 U787 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n735) );
  XNOR2_X1 U788 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n734) );
  XNOR2_X1 U789 ( .A(n735), .B(n734), .ZN(n736) );
  XOR2_X1 U790 ( .A(n737), .B(n736), .Z(n738) );
  XNOR2_X1 U791 ( .A(n739), .B(n738), .ZN(n740) );
  NOR2_X1 U792 ( .A1(n748), .A2(n740), .ZN(G54) );
  NAND2_X1 U793 ( .A1(n744), .A2(G478), .ZN(n742) );
  XNOR2_X1 U794 ( .A(n742), .B(n741), .ZN(n743) );
  NOR2_X1 U795 ( .A1(n748), .A2(n743), .ZN(G63) );
  NAND2_X1 U796 ( .A1(n744), .A2(G217), .ZN(n746) );
  XNOR2_X1 U797 ( .A(n746), .B(n745), .ZN(n747) );
  NOR2_X1 U798 ( .A1(n748), .A2(n747), .ZN(G66) );
  INV_X1 U799 ( .A(n749), .ZN(n752) );
  XOR2_X1 U800 ( .A(n750), .B(n751), .Z(n756) );
  XNOR2_X1 U801 ( .A(n752), .B(n756), .ZN(n754) );
  NAND2_X1 U802 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U803 ( .A(KEYINPUT126), .B(n755), .ZN(n761) );
  XOR2_X1 U804 ( .A(G227), .B(n756), .Z(n757) );
  NAND2_X1 U805 ( .A1(n757), .A2(G900), .ZN(n758) );
  NAND2_X1 U806 ( .A1(G953), .A2(n758), .ZN(n759) );
  XOR2_X1 U807 ( .A(KEYINPUT127), .B(n759), .Z(n760) );
  NAND2_X1 U808 ( .A1(n761), .A2(n760), .ZN(G72) );
  XNOR2_X1 U809 ( .A(G131), .B(n762), .ZN(G33) );
  XNOR2_X1 U810 ( .A(G137), .B(n763), .ZN(G39) );
endmodule

