//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n606, new_n607, new_n609, new_n610, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1150, new_n1151;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(new_n455), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n458), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT70), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n465), .A2(new_n462), .A3(G101), .A4(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n469), .A2(new_n471), .A3(G137), .A4(new_n462), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT71), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n476), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n475), .B1(new_n477), .B2(new_n462), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT71), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n467), .A2(new_n479), .A3(new_n472), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n469), .A2(new_n471), .A3(G125), .ZN(new_n481));
  NAND2_X1  g056(.A1(G113), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n483), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n474), .A2(new_n478), .A3(new_n480), .A4(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  INV_X1    g061(.A(new_n476), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  OR2_X1    g063(.A1(new_n488), .A2(KEYINPUT72), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(KEYINPUT72), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n487), .A2(new_n462), .ZN(new_n494));
  OR2_X1    g069(.A1(G100), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G112), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n468), .B1(new_n496), .B2(G2105), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n494), .A2(G124), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G162));
  NAND4_X1  g075(.A1(new_n469), .A2(new_n471), .A3(G138), .A4(new_n462), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n476), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n469), .A2(new_n471), .A3(G126), .A4(G2105), .ZN(new_n506));
  INV_X1    g081(.A(G114), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G2105), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n508), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n505), .A2(new_n510), .ZN(G164));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(G50), .A3(G543), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(new_n514), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n515), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n520), .A2(G62), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n523), .A2(new_n527), .ZN(G166));
  XOR2_X1   g103(.A(KEYINPUT74), .B(KEYINPUT7), .Z(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G89), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n512), .A2(new_n513), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n516), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G51), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n533), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n538), .A2(new_n539), .ZN(new_n541));
  OAI221_X1 g116(.A(new_n531), .B1(new_n532), .B2(new_n521), .C1(new_n540), .C2(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  NAND2_X1  g118(.A1(new_n535), .A2(G52), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OAI221_X1 g121(.A(new_n544), .B1(new_n521), .B2(new_n545), .C1(new_n546), .C2(new_n524), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(KEYINPUT75), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(KEYINPUT75), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(G171));
  NAND2_X1  g125(.A1(new_n535), .A2(G43), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n552), .B2(new_n521), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT76), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n524), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(new_n559));
  XOR2_X1   g134(.A(new_n559), .B(KEYINPUT77), .Z(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(new_n535), .A2(G53), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT9), .ZN(new_n567));
  INV_X1    g142(.A(new_n521), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G91), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n520), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n570), .A2(new_n524), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n567), .A2(new_n569), .A3(new_n571), .ZN(G299));
  INV_X1    g147(.A(G171), .ZN(G301));
  INV_X1    g148(.A(G166), .ZN(G303));
  NAND2_X1  g149(.A1(new_n568), .A2(G87), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n535), .A2(G49), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  NAND3_X1  g153(.A1(new_n517), .A2(new_n519), .A3(G86), .ZN(new_n579));
  NAND2_X1  g154(.A1(G48), .A2(G543), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n534), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n517), .A2(new_n519), .A3(G61), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n524), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n581), .A2(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n535), .A2(G47), .ZN(new_n586));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n587), .B2(new_n521), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n524), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G290));
  AND3_X1   g167(.A1(new_n520), .A2(new_n514), .A3(G92), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n535), .A2(G54), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n520), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n524), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(G171), .B2(new_n599), .ZN(G284));
  OAI21_X1  g176(.A(new_n600), .B1(G171), .B2(new_n599), .ZN(G321));
  NAND2_X1  g177(.A1(G299), .A2(new_n599), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G168), .B2(new_n599), .ZN(G297));
  OAI21_X1  g179(.A(new_n603), .B1(G168), .B2(new_n599), .ZN(G280));
  INV_X1    g180(.A(new_n598), .ZN(new_n606));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n557), .A2(new_n599), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n598), .A2(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n599), .ZN(G323));
  XOR2_X1   g186(.A(KEYINPUT78), .B(KEYINPUT11), .Z(new_n612));
  XNOR2_X1  g187(.A(G323), .B(new_n612), .ZN(G282));
  NAND2_X1  g188(.A1(new_n492), .A2(G135), .ZN(new_n614));
  NOR3_X1   g189(.A1(new_n462), .A2(KEYINPUT79), .A3(G111), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(KEYINPUT79), .B1(new_n462), .B2(G111), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n618), .B(new_n619), .C1(new_n616), .C2(new_n617), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n494), .A2(G123), .ZN(new_n621));
  AND2_X1   g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n614), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NOR2_X1   g199(.A1(new_n468), .A2(G2105), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n476), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n624), .A2(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT15), .B(G2435), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(KEYINPUT14), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT81), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n637), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT82), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n641), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G14), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT83), .ZN(G401));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT84), .Z(new_n649));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  AOI21_X1  g225(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT85), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(KEYINPUT17), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n652), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n650), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n655), .A2(new_n647), .A3(new_n648), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT18), .Z(new_n657));
  NAND3_X1  g232(.A1(new_n649), .A2(new_n653), .A3(new_n647), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2096), .B(G2100), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT86), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(KEYINPUT86), .B1(new_n663), .B2(new_n665), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n662), .A2(new_n664), .ZN(new_n676));
  OR3_X1    g251(.A1(new_n671), .A2(new_n666), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n671), .A2(new_n676), .ZN(new_n679));
  NAND4_X1  g254(.A1(new_n675), .A2(new_n677), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1991), .B(G1996), .Z(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n680), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT87), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G229));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G25), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n492), .A2(G131), .ZN(new_n691));
  OR2_X1    g266(.A1(G95), .A2(G2105), .ZN(new_n692));
  INV_X1    g267(.A(G107), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n468), .B1(new_n693), .B2(G2105), .ZN(new_n694));
  AOI22_X1  g269(.A1(new_n494), .A2(G119), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n690), .B1(new_n697), .B2(new_n689), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT35), .B(G1991), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(G16), .A2(G24), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n591), .B(KEYINPUT88), .Z(new_n703));
  AOI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(G16), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(G1986), .Z(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G22), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n706), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1971), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n706), .A2(G23), .ZN(new_n710));
  INV_X1    g285(.A(G288), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n706), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT33), .Z(new_n713));
  AOI21_X1  g288(.A(new_n709), .B1(new_n713), .B2(G1976), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n706), .A2(G6), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n581), .A2(new_n584), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n706), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT32), .B(G1981), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n714), .B(new_n719), .C1(G1976), .C2(new_n713), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT34), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n701), .B(new_n705), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT89), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n720), .B(new_n721), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n727), .A2(KEYINPUT89), .A3(new_n701), .A4(new_n705), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n726), .A2(KEYINPUT36), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n724), .A2(KEYINPUT36), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n485), .A2(G29), .ZN(new_n733));
  INV_X1    g308(.A(G2084), .ZN(new_n734));
  OR2_X1    g309(.A1(KEYINPUT24), .A2(G34), .ZN(new_n735));
  NAND2_X1  g310(.A1(KEYINPUT24), .A2(G34), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n735), .A2(new_n689), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n733), .A2(new_n734), .A3(new_n737), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n726), .A2(new_n728), .A3(KEYINPUT90), .A4(KEYINPUT36), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT94), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G16), .B2(G21), .ZN(new_n741));
  NOR2_X1   g316(.A1(G286), .A2(new_n706), .ZN(new_n742));
  MUX2_X1   g317(.A(new_n741), .B(new_n740), .S(new_n742), .Z(new_n743));
  INV_X1    g318(.A(G1966), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n689), .A2(G35), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G162), .B2(new_n689), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n745), .B1(G2090), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n706), .A2(G20), .ZN(new_n751));
  INV_X1    g326(.A(G299), .ZN(new_n752));
  OAI211_X1 g327(.A(KEYINPUT23), .B(new_n751), .C1(new_n752), .C2(new_n706), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(KEYINPUT23), .B2(new_n751), .ZN(new_n754));
  INV_X1    g329(.A(G1956), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n734), .B1(new_n733), .B2(new_n737), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n750), .B(new_n758), .C1(G2090), .C2(new_n749), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n689), .A2(G26), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n492), .A2(G140), .ZN(new_n761));
  OR2_X1    g336(.A1(G104), .A2(G2105), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n762), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n494), .A2(G128), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT91), .Z(new_n765));
  NAND3_X1  g340(.A1(new_n761), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n760), .B1(new_n767), .B2(new_n689), .ZN(new_n768));
  MUX2_X1   g343(.A(new_n760), .B(new_n768), .S(KEYINPUT28), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G2067), .ZN(new_n770));
  OAI21_X1  g345(.A(KEYINPUT92), .B1(G29), .B2(G33), .ZN(new_n771));
  OR3_X1    g346(.A1(KEYINPUT92), .A2(G29), .A3(G33), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n625), .A2(G103), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT25), .Z(new_n774));
  AOI22_X1  g349(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n775));
  INV_X1    g350(.A(G139), .ZN(new_n776));
  OAI221_X1 g351(.A(new_n774), .B1(new_n462), .B2(new_n775), .C1(new_n491), .C2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT93), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n771), .B(new_n772), .C1(new_n778), .C2(new_n689), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2072), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n706), .A2(G19), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n558), .B2(new_n706), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1341), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT31), .B(G11), .Z(new_n784));
  INV_X1    g359(.A(new_n623), .ZN(new_n785));
  INV_X1    g360(.A(G28), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(KEYINPUT30), .ZN(new_n787));
  AOI21_X1  g362(.A(G29), .B1(new_n786), .B2(KEYINPUT30), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n785), .A2(G29), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT26), .Z(new_n791));
  AOI22_X1  g366(.A1(new_n494), .A2(G129), .B1(G105), .B2(new_n625), .ZN(new_n792));
  INV_X1    g367(.A(G141), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n791), .B(new_n792), .C1(new_n491), .C2(new_n793), .ZN(new_n794));
  MUX2_X1   g369(.A(G32), .B(new_n794), .S(G29), .Z(new_n795));
  XOR2_X1   g370(.A(KEYINPUT27), .B(G1996), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n689), .A2(G27), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G164), .B2(new_n689), .ZN(new_n799));
  INV_X1    g374(.A(G2078), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n789), .A2(new_n797), .A3(new_n801), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n783), .A2(new_n784), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n606), .A2(new_n706), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G4), .B2(new_n706), .ZN(new_n805));
  INV_X1    g380(.A(G1348), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI22_X1  g382(.A1(new_n805), .A2(new_n806), .B1(new_n795), .B2(new_n796), .ZN(new_n808));
  NOR2_X1   g383(.A1(G5), .A2(G16), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G171), .B2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT95), .B(G1961), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n780), .A2(new_n803), .A3(new_n807), .A4(new_n813), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n759), .A2(new_n770), .A3(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n732), .A2(new_n738), .A3(new_n739), .A4(new_n815), .ZN(G150));
  INV_X1    g391(.A(G150), .ZN(G311));
  NAND2_X1  g392(.A1(new_n535), .A2(G55), .ZN(new_n818));
  INV_X1    g393(.A(G93), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n521), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(new_n524), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G860), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT98), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT37), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n557), .A2(new_n823), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n554), .A2(new_n556), .A3(new_n824), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n598), .A2(new_n607), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT39), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n827), .B1(new_n835), .B2(G860), .ZN(G145));
  INV_X1    g411(.A(KEYINPUT99), .ZN(new_n837));
  AND3_X1   g412(.A1(new_n506), .A2(new_n509), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n837), .B1(new_n506), .B2(new_n509), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n503), .B(new_n504), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n794), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n766), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(new_n778), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n494), .A2(G130), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n462), .A2(G118), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n468), .B1(new_n847), .B2(KEYINPUT101), .ZN(new_n848));
  OAI221_X1 g423(.A(new_n848), .B1(KEYINPUT101), .B2(new_n847), .C1(G106), .C2(G2105), .ZN(new_n849));
  INV_X1    g424(.A(G142), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n846), .B(new_n849), .C1(new_n491), .C2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n627), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n697), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n844), .A2(new_n777), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n845), .A2(KEYINPUT102), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n623), .B(new_n499), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n485), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n853), .ZN(new_n859));
  INV_X1    g434(.A(new_n854), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n844), .A2(new_n778), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n845), .A2(new_n853), .A3(new_n854), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(G37), .B1(new_n858), .B2(new_n865), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n857), .A2(KEYINPUT103), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n857), .A2(KEYINPUT103), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n862), .A2(new_n863), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g446(.A1(new_n824), .A2(new_n599), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n830), .B(new_n610), .Z(new_n873));
  NAND2_X1  g448(.A1(new_n606), .A2(G299), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n752), .A2(new_n598), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT41), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n752), .A2(KEYINPUT104), .A3(new_n598), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n874), .A2(new_n876), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n873), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n881), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n883), .B1(new_n884), .B2(new_n873), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT42), .ZN(new_n886));
  XNOR2_X1  g461(.A(G288), .B(G166), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n716), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(G290), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n886), .B(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n872), .B1(new_n890), .B2(new_n599), .ZN(G295));
  OAI21_X1  g466(.A(new_n872), .B1(new_n890), .B2(new_n599), .ZN(G331));
  NAND3_X1  g467(.A1(new_n828), .A2(G171), .A3(new_n829), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(G171), .B1(new_n828), .B2(new_n829), .ZN(new_n895));
  OAI21_X1  g470(.A(G286), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n895), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(G168), .A3(new_n893), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n881), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n882), .A2(new_n898), .A3(new_n896), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n901), .A3(new_n889), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT105), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n900), .A2(new_n901), .A3(new_n904), .A4(new_n889), .ZN(new_n905));
  AOI21_X1  g480(.A(G37), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n907));
  INV_X1    g482(.A(new_n889), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n884), .A2(new_n878), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n877), .A2(KEYINPUT41), .A3(new_n879), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n896), .A2(new_n898), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT106), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n900), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n911), .A2(KEYINPUT106), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n908), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n906), .A2(new_n907), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n889), .B1(new_n900), .B2(new_n901), .ZN(new_n917));
  AOI211_X1 g492(.A(G37), .B(new_n917), .C1(new_n903), .C2(new_n905), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n916), .B1(new_n907), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n906), .A2(KEYINPUT43), .A3(new_n915), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT44), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n921), .A2(new_n924), .ZN(G397));
  INV_X1    g500(.A(G1384), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n842), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n467), .A2(new_n479), .A3(new_n472), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n479), .B1(new_n467), .B2(new_n472), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT69), .B1(new_n483), .B2(G2105), .ZN(new_n933));
  AOI211_X1 g508(.A(new_n475), .B(new_n462), .C1(new_n481), .C2(new_n482), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n932), .A2(new_n935), .A3(G40), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n929), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(G2067), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n766), .B(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n937), .B1(new_n940), .B2(new_n794), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n942));
  INV_X1    g517(.A(new_n937), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n942), .B1(new_n943), .B2(G1996), .ZN(new_n944));
  INV_X1    g519(.A(G1996), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n937), .A2(KEYINPUT46), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n941), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  XOR2_X1   g522(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n948));
  XNOR2_X1  g523(.A(new_n947), .B(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n794), .B(G1996), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n940), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n696), .A2(new_n699), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n767), .A2(new_n938), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n943), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT125), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n943), .A2(G1986), .A3(G290), .ZN(new_n957));
  XOR2_X1   g532(.A(new_n957), .B(KEYINPUT48), .Z(new_n958));
  NOR2_X1   g533(.A1(new_n697), .A2(new_n700), .ZN(new_n959));
  NOR4_X1   g534(.A1(new_n940), .A2(new_n952), .A3(new_n959), .A4(new_n950), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n960), .A2(new_n943), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT127), .Z(new_n962));
  AOI211_X1 g537(.A(new_n949), .B(new_n956), .C1(new_n958), .C2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(G8), .B1(new_n523), .B2(new_n527), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT55), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n964), .A2(KEYINPUT108), .A3(new_n965), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n840), .A2(new_n841), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n510), .A2(KEYINPUT99), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n506), .A2(new_n509), .A3(new_n837), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n505), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT100), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(KEYINPUT45), .B(new_n926), .C1(new_n972), .C2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G40), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n485), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n926), .B1(new_n505), .B2(new_n510), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n928), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n978), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1971), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(new_n840), .B2(new_n926), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT117), .B1(new_n987), .B2(new_n936), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n505), .B1(new_n973), .B2(new_n974), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT50), .B1(new_n989), .B2(G1384), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT117), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n980), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n981), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n986), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n988), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n985), .B1(G2090), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n971), .B1(new_n996), .B2(G8), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n840), .A2(new_n926), .ZN(new_n998));
  OAI21_X1  g573(.A(G8), .B1(new_n936), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g576(.A(KEYINPUT111), .B(G8), .C1(new_n936), .C2(new_n998), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT49), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(G305), .B2(G1981), .ZN(new_n1006));
  INV_X1    g581(.A(G1981), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n716), .A2(KEYINPUT113), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(G305), .A2(KEYINPUT114), .A3(G1981), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(new_n716), .B2(new_n1007), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(new_n1014), .B2(new_n1004), .ZN(new_n1016));
  AOI211_X1 g591(.A(KEYINPUT115), .B(KEYINPUT49), .C1(new_n1009), .C2(new_n1013), .ZN(new_n1017));
  OAI221_X1 g592(.A(new_n1003), .B1(new_n1004), .B2(new_n1014), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n711), .A2(G1976), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1019), .B(KEYINPUT112), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1003), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT52), .ZN(new_n1022));
  INV_X1    g597(.A(G1976), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT52), .B1(G288), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1003), .A2(new_n1020), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1018), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT109), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n971), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n968), .A2(new_n969), .A3(KEYINPUT109), .A4(new_n970), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n983), .A2(new_n984), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n840), .A2(new_n986), .A3(new_n926), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n1032), .A2(KEYINPUT107), .B1(KEYINPUT50), .B2(new_n981), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT107), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n993), .A2(new_n1034), .A3(new_n986), .ZN(new_n1035));
  NOR4_X1   g610(.A1(new_n1033), .A2(new_n1035), .A3(G2090), .A4(new_n936), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1030), .B(G8), .C1(new_n1031), .C2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1032), .A2(KEYINPUT107), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n986), .B2(new_n993), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1035), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n980), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n985), .B1(new_n1043), .B2(G2090), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1044), .A2(KEYINPUT110), .A3(G8), .A4(new_n1030), .ZN(new_n1045));
  AOI211_X1 g620(.A(new_n997), .B(new_n1026), .C1(new_n1039), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1041), .A2(new_n734), .A3(new_n980), .A4(new_n1042), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n993), .A2(KEYINPUT45), .ZN(new_n1049));
  INV_X1    g624(.A(new_n998), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n980), .B(new_n1049), .C1(new_n1050), .C2(KEYINPUT45), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n744), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1048), .A2(G168), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1047), .B1(new_n1053), .B2(G8), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G286), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT51), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1053), .A2(G8), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1054), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT62), .ZN(new_n1060));
  AOI21_X1  g635(.A(G301), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OR2_X1    g636(.A1(new_n983), .A2(G2078), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n1063));
  INV_X1    g638(.A(G1961), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1062), .A2(new_n1063), .B1(new_n1064), .B2(new_n1043), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n800), .A2(KEYINPUT53), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1065), .B1(new_n1066), .B2(new_n1051), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1046), .A2(new_n1061), .A3(KEYINPUT124), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT124), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1039), .A2(new_n1045), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1026), .ZN(new_n1071));
  INV_X1    g646(.A(new_n997), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .A4(new_n1067), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1054), .ZN(new_n1074));
  AOI21_X1  g649(.A(G168), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1075));
  OAI211_X1 g650(.A(G8), .B(new_n1053), .C1(new_n1075), .C2(new_n1047), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1074), .A2(new_n1076), .A3(new_n1060), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G171), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1069), .B1(new_n1073), .B2(new_n1078), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1068), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1055), .A2(G8), .A3(G168), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1044), .A2(G8), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1082), .B1(new_n1083), .B2(new_n971), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT63), .B1(new_n1084), .B2(new_n1026), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1018), .A2(new_n1023), .A3(new_n711), .ZN(new_n1086));
  XOR2_X1   g661(.A(new_n1009), .B(KEYINPUT116), .Z(new_n1087));
  OAI21_X1  g662(.A(new_n1003), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT63), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1072), .A2(new_n1090), .A3(new_n1082), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1026), .B1(new_n1091), .B2(new_n1070), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1081), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT61), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n995), .A2(new_n755), .ZN(new_n1096));
  XOR2_X1   g671(.A(G299), .B(KEYINPUT57), .Z(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT56), .B(G2072), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n978), .A2(new_n980), .A3(new_n982), .A4(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1096), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1097), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1095), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n978), .A2(new_n945), .A3(new_n980), .A4(new_n982), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1050), .A2(new_n980), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT58), .B(G1341), .Z(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(new_n1108), .A3(new_n558), .ZN(new_n1109));
  AOI211_X1 g684(.A(KEYINPUT119), .B(new_n557), .C1(new_n1103), .C2(new_n1106), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1109), .B(KEYINPUT59), .C1(new_n1110), .C2(new_n1108), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1107), .A2(new_n558), .ZN(new_n1113));
  OAI211_X1 g688(.A(KEYINPUT118), .B(new_n1112), .C1(new_n1113), .C2(KEYINPUT119), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1102), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT120), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1096), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1095), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1116), .A2(new_n1117), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1117), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1115), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT122), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1115), .B(new_n1125), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1104), .A2(G2067), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(new_n1043), .B2(new_n806), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(KEYINPUT60), .B2(new_n606), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n606), .A2(KEYINPUT60), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1129), .B(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1124), .A2(new_n1126), .A3(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1128), .A2(new_n598), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1118), .B1(new_n1133), .B2(new_n1101), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  XOR2_X1   g710(.A(G171), .B(KEYINPUT54), .Z(new_n1136));
  AOI21_X1  g711(.A(new_n1059), .B1(new_n1136), .B2(new_n1067), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1136), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n932), .B(G40), .C1(new_n462), .C2(new_n477), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n1139), .A2(KEYINPUT123), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1066), .B1(new_n1139), .B2(KEYINPUT123), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n929), .A2(new_n978), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1065), .A2(new_n1138), .A3(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1137), .A2(new_n1046), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1094), .B1(new_n1135), .B2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n591), .B(G1986), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n943), .B1(new_n960), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n963), .B1(new_n1145), .B2(new_n1147), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g723(.A1(new_n645), .A2(new_n460), .ZN(new_n1150));
  AOI211_X1 g724(.A(G227), .B(new_n1150), .C1(new_n866), .C2(new_n869), .ZN(new_n1151));
  AND3_X1   g725(.A1(new_n1151), .A2(new_n687), .A3(new_n919), .ZN(G308));
  NAND3_X1  g726(.A1(new_n1151), .A2(new_n687), .A3(new_n919), .ZN(G225));
endmodule


