//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n187));
  INV_X1    g001(.A(G137), .ZN(new_n188));
  AOI21_X1  g002(.A(KEYINPUT11), .B1(new_n188), .B2(G134), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(G134), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G131), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n191), .A2(KEYINPUT64), .A3(new_n192), .A4(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n195));
  INV_X1    g009(.A(G134), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(G137), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(G137), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n197), .A2(new_n193), .A3(new_n192), .A4(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n194), .A2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n197), .A2(new_n193), .A3(new_n198), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G131), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n202), .A2(KEYINPUT67), .A3(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT67), .B1(new_n202), .B2(new_n204), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT0), .A4(G128), .ZN(new_n211));
  XNOR2_X1  g025(.A(G143), .B(G146), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT0), .B(G128), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n205), .A2(new_n206), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n188), .A2(G134), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n192), .B1(new_n216), .B2(new_n198), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n208), .A2(new_n210), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT65), .B(G128), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n220), .B1(G143), .B2(new_n207), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n218), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n212), .A2(new_n220), .A3(G128), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n217), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n202), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n187), .B1(new_n215), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g041(.A(KEYINPUT2), .B(G113), .Z(new_n228));
  XNOR2_X1  g042(.A(G116), .B(G119), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(KEYINPUT66), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT2), .B(G113), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n232));
  INV_X1    g046(.A(G116), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G119), .ZN(new_n234));
  INV_X1    g048(.A(G119), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(G116), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n231), .B(new_n232), .C1(new_n234), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n230), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n199), .A2(new_n200), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n199), .A2(new_n200), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n204), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n202), .A2(KEYINPUT67), .A3(new_n204), .ZN(new_n245));
  INV_X1    g059(.A(new_n214), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT69), .A3(new_n225), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n227), .A2(new_n239), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT28), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(G237), .A2(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G210), .ZN(new_n253));
  XOR2_X1   g067(.A(new_n253), .B(KEYINPUT27), .Z(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(G101), .ZN(new_n255));
  XOR2_X1   g069(.A(new_n254), .B(new_n255), .Z(new_n256));
  NAND2_X1  g070(.A1(new_n242), .A2(new_n246), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n225), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n238), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n247), .A2(new_n225), .A3(new_n239), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n247), .A2(KEYINPUT68), .A3(new_n225), .A4(new_n239), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n260), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n251), .B(new_n256), .C1(new_n250), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n264), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n258), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n247), .A2(new_n225), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n238), .B(new_n269), .C1(new_n270), .C2(new_n268), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n256), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT29), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n266), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n256), .A2(KEYINPUT29), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n239), .B1(new_n247), .B2(new_n225), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n277), .B1(new_n263), .B2(new_n264), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n251), .B(new_n276), .C1(new_n250), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT71), .ZN(new_n280));
  INV_X1    g094(.A(new_n277), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n267), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT28), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n283), .A2(new_n284), .A3(new_n251), .A4(new_n276), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n275), .A2(new_n280), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G472), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT32), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n267), .A2(new_n256), .A3(new_n271), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n267), .A2(KEYINPUT31), .A3(new_n256), .A4(new_n271), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n250), .B1(new_n267), .B2(new_n259), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n238), .B1(new_n270), .B2(new_n187), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT28), .B1(new_n296), .B2(new_n248), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n273), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G472), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(new_n286), .A3(KEYINPUT70), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n302), .B1(G472), .B2(G902), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n289), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n304), .ZN(new_n306));
  AOI211_X1 g120(.A(KEYINPUT32), .B(new_n306), .C1(new_n294), .C2(new_n298), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n288), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT23), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n309), .B1(new_n235), .B2(G128), .ZN(new_n310));
  INV_X1    g124(.A(G128), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(G119), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n219), .A2(KEYINPUT23), .A3(G119), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n313), .A2(KEYINPUT72), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(KEYINPUT72), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n312), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G110), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G125), .ZN(new_n322));
  OR2_X1    g136(.A1(new_n322), .A2(KEYINPUT16), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(G146), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(G146), .B1(new_n320), .B2(new_n323), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n219), .A2(G119), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n327), .B1(G119), .B2(new_n311), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT24), .B(G110), .ZN(new_n329));
  OAI22_X1  g143(.A1(new_n325), .A2(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n318), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT22), .B(G137), .ZN(new_n332));
  INV_X1    g146(.A(G953), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(G221), .A3(G234), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n332), .B(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n316), .A2(new_n317), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n328), .A2(new_n329), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n319), .A2(new_n207), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n324), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n331), .B(new_n335), .C1(new_n338), .C2(new_n340), .ZN(new_n341));
  XOR2_X1   g155(.A(new_n335), .B(KEYINPUT73), .Z(new_n342));
  AOI21_X1  g156(.A(new_n340), .B1(new_n336), .B2(new_n337), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n318), .A2(new_n330), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G217), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(G234), .B2(new_n286), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(G902), .ZN(new_n348));
  XOR2_X1   g162(.A(KEYINPUT74), .B(KEYINPUT75), .Z(new_n349));
  XNOR2_X1  g163(.A(new_n348), .B(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n341), .A2(new_n345), .A3(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(KEYINPUT76), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n347), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n341), .A2(new_n345), .A3(new_n286), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT25), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n341), .A2(new_n345), .A3(KEYINPUT25), .A4(new_n286), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n354), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT9), .B(G234), .ZN(new_n361));
  OAI21_X1  g175(.A(G221), .B1(new_n361), .B2(G902), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(G110), .B(G140), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT77), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n333), .A2(G227), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n365), .B(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G104), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT3), .B1(new_n368), .B2(G107), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT3), .ZN(new_n370));
  INV_X1    g184(.A(G107), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(G104), .ZN(new_n372));
  INV_X1    g186(.A(G101), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n368), .A2(G107), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n369), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n368), .A2(G107), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n371), .A2(G104), .ZN(new_n377));
  OAI21_X1  g191(.A(G101), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n218), .B1(new_n221), .B2(new_n311), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n223), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n379), .A2(new_n222), .A3(new_n223), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(KEYINPUT12), .A3(new_n242), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n244), .A2(new_n385), .A3(new_n245), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT12), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n387), .A2(KEYINPUT80), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT80), .B1(new_n387), .B2(new_n388), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n369), .A2(new_n372), .A3(new_n374), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G101), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT4), .A3(new_n375), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n395), .A3(G101), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n246), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n222), .A2(new_n223), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n380), .A2(new_n398), .A3(KEYINPUT10), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n383), .A2(KEYINPUT79), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT79), .B1(new_n383), .B2(new_n401), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n205), .A2(new_n206), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n367), .B1(new_n391), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(new_n405), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n367), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n410), .A2(new_n406), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n286), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G469), .ZN(new_n414));
  XOR2_X1   g228(.A(KEYINPUT81), .B(G469), .Z(new_n415));
  NOR2_X1   g229(.A1(new_n406), .A2(new_n411), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n416), .A2(new_n391), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n367), .B1(new_n407), .B2(new_n409), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n286), .B(new_n415), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n363), .B1(new_n414), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(G475), .A2(G902), .ZN(new_n421));
  XNOR2_X1  g235(.A(G113), .B(G122), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT88), .B(G104), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n319), .A2(KEYINPUT19), .ZN(new_n425));
  INV_X1    g239(.A(G125), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G140), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n322), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT85), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT85), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n319), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n425), .B1(new_n432), .B2(KEYINPUT19), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT87), .B1(new_n433), .B2(G146), .ZN(new_n434));
  INV_X1    g248(.A(G237), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(new_n333), .A3(G214), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n209), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n252), .A2(G143), .A3(G214), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G131), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT86), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT86), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(new_n442), .A3(G131), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n437), .A2(new_n192), .A3(new_n438), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT87), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT19), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n429), .B2(new_n431), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n446), .B(new_n207), .C1(new_n448), .C2(new_n425), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n434), .A2(new_n324), .A3(new_n445), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(KEYINPUT18), .A2(G131), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n439), .B(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n339), .B1(new_n432), .B2(new_n207), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n424), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT17), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n441), .A2(new_n456), .A3(new_n443), .A4(new_n444), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n442), .B1(new_n439), .B2(G131), .ZN(new_n458));
  AOI211_X1 g272(.A(KEYINPUT86), .B(new_n192), .C1(new_n437), .C2(new_n438), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT17), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n325), .A2(new_n326), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n462), .A2(new_n424), .A3(new_n454), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n421), .B1(new_n455), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT20), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n466));
  INV_X1    g280(.A(new_n421), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT89), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n468), .B2(new_n467), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n470), .B1(new_n455), .B2(new_n463), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT90), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g287(.A(KEYINPUT90), .B(new_n470), .C1(new_n455), .C2(new_n463), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n465), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n424), .B1(new_n462), .B2(new_n454), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n286), .B1(new_n463), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G475), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT91), .B1(new_n233), .B2(G122), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT91), .ZN(new_n481));
  INV_X1    g295(.A(G122), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n482), .A3(G116), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n233), .A2(G122), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(KEYINPUT14), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n487), .A3(G107), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n484), .B(new_n485), .C1(KEYINPUT14), .C2(new_n371), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n311), .A2(KEYINPUT65), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT65), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G128), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n492), .A3(G143), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n209), .A2(G128), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n196), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n196), .B1(new_n493), .B2(new_n494), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n488), .B(new_n489), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT13), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n494), .A2(new_n499), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n493), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n500), .B1(new_n502), .B2(KEYINPUT92), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT92), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n493), .A2(new_n504), .A3(new_n501), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n196), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n486), .A2(G107), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n371), .B1(new_n484), .B2(new_n485), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n495), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n498), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n361), .A2(new_n346), .A3(G953), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n498), .B(new_n511), .C1(new_n506), .C2(new_n509), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n286), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT93), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G478), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(KEYINPUT15), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n515), .A2(KEYINPUT93), .A3(new_n286), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(G952), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(G953), .ZN(new_n524));
  INV_X1    g338(.A(G234), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n524), .B1(new_n525), .B2(new_n435), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(G902), .B(G953), .C1(new_n525), .C2(new_n435), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT94), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT21), .B(G898), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n516), .A2(new_n520), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n522), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(G214), .B1(G237), .B2(G902), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n394), .A2(new_n238), .A3(new_n396), .ZN(new_n536));
  OR2_X1    g350(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n537));
  NAND2_X1  g351(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n234), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT83), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n537), .A2(new_n538), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n229), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT83), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n234), .A2(new_n537), .A3(new_n543), .A4(new_n538), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n540), .A2(G113), .A3(new_n542), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n228), .A2(new_n229), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n380), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(G110), .B(G122), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n536), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n214), .A2(G125), .ZN(new_n550));
  INV_X1    g364(.A(G224), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT7), .B1(new_n551), .B2(G953), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  OAI221_X1 g367(.A(new_n550), .B1(KEYINPUT84), .B2(new_n553), .C1(G125), .C2(new_n398), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n553), .B1(new_n550), .B2(KEYINPUT84), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n550), .B1(G125), .B2(new_n398), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n549), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  XOR2_X1   g373(.A(new_n548), .B(KEYINPUT8), .Z(new_n560));
  NAND2_X1  g374(.A1(new_n229), .A2(KEYINPUT5), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n540), .A2(G113), .A3(new_n544), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n546), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n560), .B1(new_n563), .B2(new_n380), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n545), .A2(new_n379), .A3(new_n546), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(G902), .B1(new_n559), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n536), .A2(new_n547), .ZN(new_n568));
  INV_X1    g382(.A(new_n548), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(KEYINPUT6), .A3(new_n549), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n551), .A2(G953), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n556), .B(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT6), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n568), .A2(new_n574), .A3(new_n569), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n571), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(G210), .B1(G237), .B2(G902), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n567), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n577), .B1(new_n567), .B2(new_n576), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n535), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n479), .A2(new_n534), .A3(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n308), .A2(new_n360), .A3(new_n420), .A4(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(G101), .ZN(G3));
  NAND3_X1  g397(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n515), .A2(KEYINPUT33), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT33), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n513), .B2(new_n514), .ZN(new_n587));
  OAI211_X1 g401(.A(G478), .B(new_n286), .C1(new_n585), .C2(new_n587), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n475), .A2(new_n478), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n577), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n571), .A2(new_n573), .A3(new_n575), .ZN(new_n591));
  INV_X1    g405(.A(new_n566), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n286), .B1(new_n592), .B2(new_n558), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n590), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n567), .A2(new_n576), .A3(new_n577), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT95), .B1(new_n596), .B2(new_n535), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n598));
  INV_X1    g412(.A(new_n535), .ZN(new_n599));
  AOI211_X1 g413(.A(new_n598), .B(new_n599), .C1(new_n594), .C2(new_n595), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n589), .B(new_n532), .C1(new_n597), .C2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT96), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n580), .A2(new_n598), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n596), .A2(KEYINPUT95), .A3(new_n535), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT96), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n605), .A2(new_n606), .A3(new_n532), .A4(new_n589), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n420), .A2(new_n360), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n294), .B2(new_n298), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n251), .B1(new_n250), .B2(new_n265), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n292), .A2(new_n293), .B1(new_n611), .B2(new_n273), .ZN(new_n612));
  OAI22_X1  g426(.A1(new_n610), .A2(new_n300), .B1(new_n612), .B2(new_n306), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT97), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT34), .B(G104), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  INV_X1    g432(.A(new_n605), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n619), .A2(new_n531), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n522), .A2(new_n533), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n465), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n466), .B(new_n421), .C1(new_n455), .C2(new_n463), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n478), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n614), .A2(new_n620), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(new_n371), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT98), .B(KEYINPUT35), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  INV_X1    g445(.A(new_n359), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n343), .A2(new_n344), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n342), .A2(KEYINPUT36), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n633), .B(new_n634), .Z(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n350), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n420), .A2(new_n581), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n613), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT37), .B(G110), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G12));
  INV_X1    g456(.A(G900), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n527), .B1(new_n529), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n478), .B(new_n645), .C1(new_n623), .C2(new_n625), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n622), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n637), .A2(new_n605), .A3(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n308), .A2(new_n420), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT99), .ZN(new_n651));
  INV_X1    g465(.A(new_n420), .ZN(new_n652));
  OAI21_X1  g466(.A(KEYINPUT32), .B1(new_n612), .B2(new_n306), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n299), .A2(new_n289), .A3(new_n304), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n652), .B1(new_n655), .B2(new_n288), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n657), .A3(new_n649), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  XNOR2_X1  g474(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n644), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n420), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n663), .B(KEYINPUT40), .Z(new_n664));
  NAND2_X1  g478(.A1(new_n272), .A2(new_n256), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n665), .B(new_n286), .C1(new_n256), .C2(new_n282), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(G472), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n655), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n479), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n622), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n359), .B1(new_n350), .B2(new_n635), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n670), .A2(new_n671), .A3(new_n535), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n596), .B(KEYINPUT38), .Z(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n664), .A2(new_n668), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT101), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n209), .ZN(G45));
  NAND2_X1  g491(.A1(new_n584), .A2(new_n588), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n479), .A2(new_n678), .A3(new_n645), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n619), .A2(new_n671), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n656), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G146), .ZN(G48));
  OAI21_X1  g496(.A(new_n286), .B1(new_n417), .B2(new_n418), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(G469), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n419), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n363), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n608), .A2(new_n308), .A3(new_n360), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT41), .B(G113), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  NOR3_X1   g503(.A1(new_n619), .A2(new_n685), .A3(new_n363), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n632), .A2(new_n352), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n531), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n308), .A2(new_n690), .A3(new_n627), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G116), .ZN(G18));
  NOR3_X1   g508(.A1(new_n671), .A2(new_n479), .A3(new_n534), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n308), .A2(new_n690), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT102), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT102), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n308), .A2(new_n690), .A3(new_n698), .A4(new_n695), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G119), .ZN(G21));
  NAND3_X1  g515(.A1(new_n620), .A2(new_n670), .A3(new_n686), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT104), .B(G472), .Z(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n705), .B1(new_n612), .B2(G902), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n304), .B(KEYINPUT103), .Z(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n250), .B1(new_n267), .B2(new_n281), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n273), .B1(new_n709), .B2(new_n297), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n708), .B1(new_n294), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n706), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n703), .B1(new_n713), .B2(new_n691), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n706), .A2(KEYINPUT105), .A3(new_n360), .A4(new_n712), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n702), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n482), .ZN(G24));
  AOI21_X1  g531(.A(new_n704), .B1(new_n299), .B2(new_n286), .ZN(new_n718));
  NOR4_X1   g532(.A1(new_n718), .A2(new_n671), .A3(new_n679), .A4(new_n711), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n719), .A2(new_n690), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n426), .ZN(G27));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n413), .B2(G469), .ZN(new_n723));
  INV_X1    g537(.A(new_n386), .ZN(new_n724));
  INV_X1    g538(.A(new_n390), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n387), .A2(KEYINPUT80), .A3(new_n388), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n411), .B1(new_n727), .B2(new_n406), .ZN(new_n728));
  INV_X1    g542(.A(new_n412), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n722), .A2(new_n286), .A3(G469), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n419), .B1(new_n723), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n596), .A2(new_n599), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n733), .A2(new_n362), .A3(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n679), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n735), .A2(new_n308), .A3(new_n360), .A4(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI22_X1  g553(.A1(new_n653), .A2(new_n654), .B1(new_n287), .B2(G472), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n691), .ZN(new_n741));
  INV_X1    g555(.A(new_n738), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(new_n736), .A3(new_n735), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  NAND4_X1  g559(.A1(new_n735), .A2(new_n308), .A3(new_n360), .A4(new_n647), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G134), .ZN(G36));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n730), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n728), .A2(new_n729), .A3(KEYINPUT45), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n750), .A3(G469), .ZN(new_n751));
  NAND2_X1  g565(.A1(G469), .A2(G902), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT46), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n751), .A2(KEYINPUT46), .A3(new_n752), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n419), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n362), .A3(new_n662), .ZN(new_n758));
  XOR2_X1   g572(.A(new_n758), .B(KEYINPUT108), .Z(new_n759));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT43), .B1(new_n669), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n669), .A2(new_n678), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n613), .A3(new_n637), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n734), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n766), .B1(new_n765), .B2(new_n764), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n759), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  NAND2_X1  g583(.A1(new_n757), .A2(new_n362), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(KEYINPUT47), .Z(new_n771));
  INV_X1    g585(.A(new_n734), .ZN(new_n772));
  NOR4_X1   g586(.A1(new_n308), .A2(new_n360), .A3(new_n679), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n321), .ZN(G42));
  AND2_X1   g591(.A1(new_n763), .A2(new_n527), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n686), .A3(new_n734), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT120), .Z(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n741), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT48), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n686), .A2(new_n360), .A3(new_n527), .A4(new_n734), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n783), .A2(new_n668), .ZN(new_n784));
  INV_X1    g598(.A(new_n589), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n524), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n714), .A2(new_n715), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n778), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n786), .B1(new_n789), .B2(new_n690), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n789), .A2(new_n599), .A3(new_n673), .A4(new_n686), .ZN(new_n791));
  XOR2_X1   g605(.A(new_n791), .B(KEYINPUT50), .Z(new_n792));
  NOR3_X1   g606(.A1(new_n784), .A2(new_n479), .A3(new_n678), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n713), .A2(new_n671), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n793), .B1(new_n780), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n788), .A2(new_n772), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n685), .A2(new_n362), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n797), .B1(new_n771), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT51), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n782), .B(new_n790), .C1(new_n796), .C2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n796), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n798), .B(KEYINPUT119), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n797), .B1(new_n771), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT51), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g620(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n656), .A2(new_n680), .B1(new_n719), .B2(new_n690), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n733), .A2(new_n362), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n670), .A2(new_n605), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n637), .A2(new_n644), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n668), .A2(new_n810), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n657), .B1(new_n656), .B2(new_n649), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n740), .A2(KEYINPUT99), .A3(new_n652), .A4(new_n648), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n809), .B(new_n813), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT52), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n659), .A2(new_n818), .A3(new_n809), .A4(new_n813), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n817), .A2(KEYINPUT114), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT114), .B1(new_n817), .B2(new_n819), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n687), .A2(new_n693), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(new_n716), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n824), .A2(new_n744), .A3(KEYINPUT53), .A4(new_n700), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n596), .A2(new_n535), .A3(new_n532), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT112), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n621), .A2(new_n475), .A3(new_n478), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n589), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n669), .A2(KEYINPUT112), .A3(new_n621), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n826), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n614), .A2(new_n831), .B1(new_n638), .B2(new_n639), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n671), .A2(new_n772), .A3(new_n621), .A4(new_n646), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n308), .A2(new_n420), .A3(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n832), .A2(new_n746), .A3(new_n582), .A4(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT113), .B1(new_n719), .B2(new_n735), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n733), .A2(new_n362), .A3(new_n734), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n706), .A2(new_n736), .A3(new_n712), .A4(new_n637), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n835), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT117), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(new_n835), .B2(new_n841), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n825), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n842), .A2(new_n700), .A3(new_n744), .A4(new_n824), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n817), .A2(new_n819), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT116), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n852), .B(new_n847), .C1(new_n848), .C2(new_n849), .ZN(new_n853));
  AOI221_X4 g667(.A(new_n808), .B1(new_n822), .B2(new_n846), .C1(new_n851), .C2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n820), .A2(new_n821), .A3(new_n848), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n824), .A2(new_n744), .A3(new_n700), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(new_n842), .A3(new_n819), .A4(new_n817), .ZN(new_n857));
  OAI22_X1  g671(.A1(new_n855), .A2(KEYINPUT53), .B1(new_n857), .B2(new_n847), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n854), .B1(new_n858), .B2(KEYINPUT54), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n806), .A2(new_n859), .B1(new_n523), .B2(new_n333), .ZN(new_n860));
  NOR4_X1   g674(.A1(new_n762), .A2(new_n691), .A3(new_n363), .A4(new_n599), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n685), .A2(KEYINPUT49), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n673), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n685), .A2(KEYINPUT49), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n863), .A2(new_n668), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT111), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n860), .A2(new_n866), .ZN(G75));
  NOR2_X1   g681(.A1(new_n333), .A2(G952), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n822), .A2(new_n846), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n852), .B1(new_n857), .B2(new_n847), .ZN(new_n871));
  INV_X1    g685(.A(new_n853), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n286), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT56), .B1(new_n875), .B2(G210), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n571), .A2(new_n575), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(new_n573), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT55), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n869), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n876), .B2(new_n880), .ZN(G51));
  NAND2_X1  g696(.A1(new_n873), .A2(new_n808), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n851), .A2(new_n853), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(new_n807), .A3(new_n870), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n752), .B(KEYINPUT57), .ZN(new_n888));
  OAI22_X1  g702(.A1(new_n887), .A2(new_n888), .B1(new_n418), .B2(new_n417), .ZN(new_n889));
  OR3_X1    g703(.A1(new_n874), .A2(new_n286), .A3(new_n751), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n868), .B1(new_n889), .B2(new_n890), .ZN(G54));
  OR2_X1    g705(.A1(new_n455), .A2(new_n463), .ZN(new_n892));
  AND2_X1   g706(.A1(KEYINPUT58), .A2(G475), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n875), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n892), .B1(new_n875), .B2(new_n893), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n895), .A3(new_n868), .ZN(G60));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n585), .A2(new_n587), .ZN(new_n899));
  NAND2_X1  g713(.A1(G478), .A2(G902), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT59), .Z(new_n901));
  NOR2_X1   g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n807), .B1(new_n884), .B2(new_n870), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n898), .B(new_n902), .C1(new_n854), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n869), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n898), .B1(new_n886), .B2(new_n902), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n897), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n902), .B1(new_n854), .B2(new_n903), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT121), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(KEYINPUT122), .A3(new_n869), .A4(new_n904), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n899), .B1(new_n859), .B2(new_n901), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n907), .A2(new_n910), .A3(new_n911), .ZN(G63));
  NAND2_X1  g726(.A1(G217), .A2(G902), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT123), .Z(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT60), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n874), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n635), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n341), .A2(new_n345), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n874), .B2(new_n915), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n869), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(G66));
  INV_X1    g736(.A(new_n530), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n333), .B1(new_n923), .B2(G224), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n824), .A2(new_n700), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n832), .A2(new_n582), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n924), .B1(new_n927), .B2(new_n333), .ZN(new_n928));
  INV_X1    g742(.A(G898), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n877), .B1(new_n929), .B2(G953), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n928), .B(new_n930), .ZN(G69));
  AOI21_X1  g745(.A(new_n772), .B1(new_n829), .B2(new_n830), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n741), .A2(new_n420), .A3(new_n662), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n768), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n776), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n659), .A2(new_n809), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n676), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT62), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n333), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n269), .B1(new_n270), .B2(new_n268), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT124), .Z(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(new_n433), .Z(new_n943));
  NAND3_X1  g757(.A1(new_n940), .A2(KEYINPUT125), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT125), .ZN(new_n945));
  AOI21_X1  g759(.A(G953), .B1(new_n935), .B2(new_n938), .ZN(new_n946));
  INV_X1    g760(.A(new_n943), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n741), .A2(new_n811), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n759), .B1(new_n767), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n659), .A2(new_n809), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n950), .A2(new_n744), .A3(new_n746), .A4(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n333), .B1(new_n776), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n643), .A2(G953), .ZN(new_n954));
  AOI21_X1  g768(.A(KEYINPUT126), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n953), .A2(KEYINPUT126), .A3(new_n954), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n947), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n944), .B(new_n948), .C1(new_n955), .C2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n333), .B1(G227), .B2(G900), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(G72));
  XNOR2_X1  g774(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n300), .A2(new_n286), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n272), .A2(new_n273), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n290), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n858), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n869), .B1(new_n965), .B2(new_n963), .ZN(new_n967));
  OR4_X1    g781(.A1(new_n256), .A2(new_n776), .A3(new_n952), .A4(new_n272), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n665), .B2(new_n939), .ZN(new_n969));
  INV_X1    g783(.A(new_n927), .ZN(new_n970));
  AOI211_X1 g784(.A(new_n966), .B(new_n967), .C1(new_n969), .C2(new_n970), .ZN(G57));
endmodule


