//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n547, new_n548, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n562, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT67), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(KEYINPUT3), .A3(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n464), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n469), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND3_X1  g054(.A1(new_n464), .A2(G2105), .A3(new_n467), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT68), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(new_n465), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n468), .A2(G136), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n482), .A2(new_n486), .ZN(G162));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n464), .A2(new_n467), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n472), .ZN(new_n491));
  NOR3_X1   g066(.A1(new_n488), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n490), .A2(KEYINPUT4), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n464), .A2(G126), .A3(G2105), .A4(new_n467), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  XNOR2_X1  g070(.A(KEYINPUT69), .B(G114), .ZN(new_n496));
  OAI211_X1 g071(.A(G2104), .B(new_n495), .C1(new_n496), .C2(new_n465), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n493), .A2(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT71), .B1(new_n500), .B2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n502), .A2(new_n503), .A3(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(KEYINPUT70), .ZN(new_n511));
  XNOR2_X1  g086(.A(new_n511), .B(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n510), .A2(new_n517), .ZN(G166));
  INV_X1    g093(.A(new_n513), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G89), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n524), .B2(new_n515), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n520), .B(new_n522), .C1(new_n525), .C2(KEYINPUT72), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n525), .A2(KEYINPUT72), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(G168));
  AOI22_X1  g103(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n509), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n513), .A2(new_n531), .B1(new_n515), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(G171));
  AOI22_X1  g109(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n509), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n507), .A2(G81), .A3(new_n512), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n512), .A2(G43), .A3(G543), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(KEYINPUT73), .A3(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(KEYINPUT73), .B1(new_n537), .B2(new_n538), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n536), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n545));
  XOR2_X1   g120(.A(new_n545), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  INV_X1    g124(.A(G53), .ZN(new_n550));
  OR3_X1    g125(.A1(new_n515), .A2(KEYINPUT9), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(KEYINPUT9), .B1(new_n515), .B2(new_n550), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n551), .A2(new_n552), .B1(G91), .B2(new_n519), .ZN(new_n553));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(new_n507), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n553), .B1(new_n509), .B2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(G168), .ZN(G286));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  XNOR2_X1  g137(.A(G166), .B(new_n562), .ZN(G303));
  INV_X1    g138(.A(G87), .ZN(new_n564));
  OR3_X1    g139(.A1(new_n513), .A2(KEYINPUT76), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT76), .B1(new_n513), .B2(new_n564), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n507), .A2(G74), .ZN(new_n568));
  INV_X1    g143(.A(new_n515), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n568), .A2(G651), .B1(new_n569), .B2(G49), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(G288));
  AOI22_X1  g146(.A1(new_n519), .A2(G86), .B1(new_n569), .B2(G48), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n505), .A2(G61), .A3(new_n506), .ZN(new_n573));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT77), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT78), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n578), .B(G651), .C1(new_n573), .C2(new_n575), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n572), .A2(new_n577), .A3(new_n579), .ZN(G305));
  INV_X1    g155(.A(G85), .ZN(new_n581));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n513), .A2(new_n581), .B1(new_n515), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n583), .A2(new_n584), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n585), .A2(new_n586), .B1(new_n509), .B2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n519), .A2(G92), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n555), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G54), .B2(new_n569), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n589), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n589), .B1(new_n598), .B2(G868), .ZN(G321));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  OR3_X1    g176(.A1(G168), .A2(KEYINPUT80), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(KEYINPUT80), .B1(G168), .B2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(G299), .A2(new_n601), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(G297));
  NAND3_X1  g180(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n598), .B1(new_n607), .B2(G860), .ZN(G148));
  NOR2_X1   g183(.A1(new_n543), .A2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n598), .A2(new_n607), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT81), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n491), .A2(new_n476), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT13), .Z(new_n616));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G2100), .ZN(new_n618));
  INV_X1    g193(.A(G2100), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(KEYINPUT82), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n481), .A2(G123), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n465), .A2(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n468), .A2(G135), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G2096), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n616), .A2(new_n617), .A3(G2100), .ZN(new_n628));
  INV_X1    g203(.A(G2096), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n621), .A2(new_n629), .A3(new_n625), .ZN(new_n630));
  NAND4_X1  g205(.A1(new_n620), .A2(new_n627), .A3(new_n628), .A4(new_n630), .ZN(G156));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT83), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT14), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n640), .B2(new_n639), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n636), .B(new_n642), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(G14), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n644), .ZN(G401));
  INV_X1    g223(.A(KEYINPUT18), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(new_n619), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n652), .B2(KEYINPUT18), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(new_n629), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1956), .B(G2474), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n662), .A2(new_n667), .A3(new_n665), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n662), .A2(new_n667), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n670));
  AOI211_X1 g245(.A(new_n666), .B(new_n668), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(new_n669), .B2(new_n670), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT85), .ZN(new_n673));
  XOR2_X1   g248(.A(G1991), .B(G1996), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT86), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n675), .B(new_n679), .ZN(G229));
  INV_X1    g255(.A(G288), .ZN(new_n681));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n682), .B2(G23), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT33), .B(G1976), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n686), .ZN(new_n688));
  NOR2_X1   g263(.A1(G166), .A2(new_n682), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n682), .B2(G22), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n691), .A2(G1971), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(G1971), .ZN(new_n693));
  NAND4_X1  g268(.A1(new_n687), .A2(new_n688), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G6), .B(G305), .S(G16), .Z(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT32), .B(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  OR3_X1    g272(.A1(new_n694), .A2(KEYINPUT34), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(KEYINPUT34), .B1(new_n694), .B2(new_n697), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n481), .A2(G119), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n468), .A2(G131), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n465), .A2(G107), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n700), .B(new_n701), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT87), .Z(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G29), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G25), .B2(G29), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT35), .B(G1991), .Z(new_n708));
  AND2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  MUX2_X1   g285(.A(G24), .B(G290), .S(G16), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G1986), .ZN(new_n712));
  NOR3_X1   g287(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n698), .A2(new_n699), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT36), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n682), .A2(G20), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT23), .Z(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G299), .B2(G16), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(G1956), .Z(new_n719));
  NOR2_X1   g294(.A1(G29), .A2(G35), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G162), .B2(G29), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n719), .B1(new_n723), .B2(G2090), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT95), .Z(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G33), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n468), .A2(G139), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT90), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT89), .B(KEYINPUT25), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  NAND2_X1  g309(.A1(G115), .A2(G2104), .ZN(new_n735));
  INV_X1    g310(.A(G127), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n472), .B2(new_n736), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n733), .A2(new_n734), .B1(G2105), .B2(new_n737), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n729), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n727), .B1(new_n739), .B2(new_n726), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(G2072), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n682), .A2(G21), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G168), .B2(new_n682), .ZN(new_n743));
  INV_X1    g318(.A(G1966), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n481), .A2(G129), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n468), .A2(G141), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT26), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n476), .A2(G105), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n747), .A2(new_n748), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  MUX2_X1   g327(.A(G32), .B(new_n752), .S(G29), .Z(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT27), .Z(new_n754));
  OAI22_X1  g329(.A1(new_n754), .A2(G1996), .B1(G2090), .B2(new_n723), .ZN(new_n755));
  AOI211_X1 g330(.A(new_n746), .B(new_n755), .C1(G1996), .C2(new_n754), .ZN(new_n756));
  NOR2_X1   g331(.A1(G171), .A2(new_n682), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G5), .B2(new_n682), .ZN(new_n758));
  INV_X1    g333(.A(G1961), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT93), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n543), .A2(G16), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G16), .B2(G19), .ZN(new_n763));
  INV_X1    g338(.A(G1341), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n726), .A2(G26), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT28), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n481), .A2(G128), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n465), .A2(G116), .ZN(new_n769));
  OAI21_X1  g344(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n468), .A2(G140), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n767), .B1(new_n773), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2067), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n761), .A2(new_n765), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G4), .A2(G16), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n598), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT88), .B(G1348), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n764), .B2(new_n763), .ZN(new_n781));
  INV_X1    g356(.A(G2078), .ZN(new_n782));
  NOR2_X1   g357(.A1(G164), .A2(new_n726), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G27), .B2(new_n726), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n758), .A2(new_n759), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G34), .ZN(new_n786));
  AOI21_X1  g361(.A(G29), .B1(new_n786), .B2(KEYINPUT24), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(KEYINPUT24), .B2(new_n786), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n478), .B2(new_n726), .ZN(new_n789));
  INV_X1    g364(.A(G2084), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(KEYINPUT91), .ZN(new_n793));
  INV_X1    g368(.A(new_n784), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n794), .A2(G2078), .B1(new_n792), .B2(KEYINPUT91), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT31), .B(G11), .Z(new_n796));
  INV_X1    g371(.A(KEYINPUT30), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n726), .B1(new_n797), .B2(G28), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n799), .A2(KEYINPUT92), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n799), .A2(KEYINPUT92), .B1(new_n797), .B2(G28), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n796), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n626), .B2(new_n726), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n790), .B2(new_n789), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n785), .A2(new_n793), .A3(new_n795), .A4(new_n804), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n776), .A2(new_n781), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n715), .A2(new_n725), .A3(new_n756), .A4(new_n806), .ZN(G150));
  INV_X1    g382(.A(G150), .ZN(G311));
  AOI22_X1  g383(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n809), .A2(new_n509), .ZN(new_n810));
  INV_X1    g385(.A(G93), .ZN(new_n811));
  INV_X1    g386(.A(G55), .ZN(new_n812));
  OAI22_X1  g387(.A1(new_n513), .A2(new_n811), .B1(new_n515), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G860), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT97), .B(KEYINPUT37), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n597), .A2(new_n607), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  INV_X1    g395(.A(new_n814), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT96), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n536), .B(new_n822), .C1(new_n540), .C2(new_n541), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n537), .A2(new_n538), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT73), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(new_n539), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n822), .B1(new_n828), .B2(new_n536), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n821), .B1(new_n824), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n542), .A2(KEYINPUT96), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n831), .A2(new_n814), .A3(new_n823), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n820), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n815), .B1(new_n835), .B2(KEYINPUT39), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n818), .B1(new_n836), .B2(new_n837), .ZN(G145));
  INV_X1    g413(.A(KEYINPUT100), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n739), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n752), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n773), .ZN(new_n842));
  INV_X1    g417(.A(new_n498), .ZN(new_n843));
  AOI221_X4 g418(.A(KEYINPUT98), .B1(new_n491), .B2(new_n492), .C1(new_n490), .C2(KEYINPUT4), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n491), .A2(new_n492), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n843), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT99), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g426(.A(KEYINPUT99), .B(new_n843), .C1(new_n844), .C2(new_n848), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n842), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n842), .A2(new_n853), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n468), .A2(G142), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n465), .A2(G118), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(G130), .B2(new_n481), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(new_n615), .Z(new_n861));
  XOR2_X1   g436(.A(new_n705), .B(new_n861), .Z(new_n862));
  NAND3_X1  g437(.A1(new_n854), .A2(new_n855), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n854), .A2(new_n855), .ZN(new_n866));
  INV_X1    g441(.A(new_n862), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n868), .A2(KEYINPUT101), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(KEYINPUT101), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n865), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n626), .B(new_n478), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(G162), .Z(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n873), .B1(new_n866), .B2(new_n867), .ZN(new_n875));
  AOI21_X1  g450(.A(G37), .B1(new_n875), .B2(new_n863), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n874), .A2(KEYINPUT40), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT40), .B1(new_n874), .B2(new_n876), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(G395));
  XOR2_X1   g454(.A(new_n833), .B(new_n610), .Z(new_n880));
  NAND2_X1  g455(.A1(new_n597), .A2(G299), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n597), .A2(G299), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(new_n882), .B2(new_n883), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n597), .A2(G299), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n889), .A2(KEYINPUT41), .A3(new_n881), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n880), .A2(new_n891), .ZN(new_n892));
  OR3_X1    g467(.A1(new_n886), .A2(new_n892), .A3(KEYINPUT104), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT104), .B1(new_n886), .B2(new_n892), .ZN(new_n894));
  XNOR2_X1  g469(.A(G290), .B(G166), .ZN(new_n895));
  XOR2_X1   g470(.A(G288), .B(G305), .Z(new_n896));
  OR2_X1    g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n896), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n899), .A2(KEYINPUT42), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT103), .B1(new_n897), .B2(new_n898), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n897), .A2(KEYINPUT103), .A3(new_n898), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n900), .B1(new_n904), .B2(KEYINPUT42), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n893), .A2(new_n894), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n905), .B1(new_n893), .B2(new_n894), .ZN(new_n907));
  OAI21_X1  g482(.A(G868), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n821), .A2(new_n601), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(G295));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n911));
  XNOR2_X1  g486(.A(G295), .B(new_n911), .ZN(G331));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n831), .A2(new_n814), .A3(new_n823), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n814), .B1(new_n831), .B2(new_n823), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n915), .A2(new_n916), .A3(G171), .ZN(new_n917));
  AOI21_X1  g492(.A(G301), .B1(new_n830), .B2(new_n832), .ZN(new_n918));
  OAI21_X1  g493(.A(G286), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(G171), .B1(new_n915), .B2(new_n916), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n830), .A2(G301), .A3(new_n832), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n921), .A3(G168), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n919), .A2(new_n884), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n888), .A2(new_n890), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n924), .B1(new_n919), .B2(new_n922), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n914), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n919), .A2(new_n884), .A3(new_n922), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT106), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n904), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n903), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n930), .A2(new_n901), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n917), .A2(new_n918), .A3(G286), .ZN(new_n932));
  AOI21_X1  g507(.A(G168), .B1(new_n920), .B2(new_n921), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n891), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n927), .ZN(new_n935));
  AOI21_X1  g510(.A(G37), .B1(new_n931), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n929), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n913), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n938), .B2(new_n937), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n930), .A2(new_n901), .A3(KEYINPUT107), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT106), .B1(new_n934), .B2(new_n927), .ZN(new_n942));
  INV_X1    g517(.A(new_n928), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n902), .A2(new_n945), .A3(new_n903), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n926), .A2(new_n928), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G37), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n944), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n940), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n929), .A2(new_n936), .A3(new_n913), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT108), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n929), .A2(new_n936), .A3(new_n954), .A4(new_n913), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n951), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n957), .B1(new_n956), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n950), .B1(new_n959), .B2(new_n960), .ZN(G397));
  INV_X1    g536(.A(new_n853), .ZN(new_n962));
  XOR2_X1   g537(.A(KEYINPUT111), .B(G1384), .Z(new_n963));
  AOI21_X1  g538(.A(KEYINPUT45), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n469), .A2(G40), .A3(new_n475), .A4(new_n477), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n773), .B(G2067), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT114), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n752), .B(G1996), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n971), .A2(new_n705), .A3(new_n708), .A4(new_n973), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n773), .A2(G2067), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n967), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OR3_X1    g551(.A1(new_n967), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT46), .B1(new_n967), .B2(G1996), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n969), .A2(new_n752), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n977), .A2(new_n978), .B1(new_n968), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT47), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n705), .B(new_n708), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n968), .ZN(new_n983));
  OR2_X1    g558(.A1(G290), .A2(G1986), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n967), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT48), .Z(new_n986));
  AND4_X1   g561(.A1(new_n983), .A2(new_n986), .A3(new_n971), .A4(new_n973), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n976), .A2(new_n981), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n989));
  INV_X1    g564(.A(G1384), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n989), .B(new_n990), .C1(new_n493), .C2(new_n498), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n966), .A2(new_n991), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n849), .A2(new_n990), .ZN(new_n993));
  OAI211_X1 g568(.A(KEYINPUT118), .B(new_n992), .C1(new_n993), .C2(new_n989), .ZN(new_n994));
  INV_X1    g569(.A(G2090), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT118), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n989), .B1(new_n849), .B2(new_n990), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n966), .A2(new_n991), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n996), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n994), .A2(new_n995), .A3(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n990), .B1(new_n493), .B2(new_n498), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n966), .B1(new_n1002), .B2(KEYINPUT45), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n963), .A2(KEYINPUT45), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n851), .A2(new_n852), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT115), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n851), .A2(new_n1007), .A3(new_n852), .A4(new_n1004), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1003), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1000), .B1(new_n1009), .B2(G1971), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g587(.A(KEYINPUT119), .B(new_n1000), .C1(new_n1009), .C2(G1971), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(G8), .A3(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(G303), .B(G8), .C1(KEYINPUT116), .C2(KEYINPUT55), .ZN(new_n1015));
  AND2_X1   g590(.A1(G303), .A2(G8), .ZN(new_n1016));
  XOR2_X1   g591(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n1017));
  OAI21_X1  g592(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1014), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1009), .A2(G1971), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n849), .A2(new_n989), .A3(new_n990), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n965), .B1(new_n1001), .B2(KEYINPUT50), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(G2090), .ZN(new_n1026));
  OAI211_X1 g601(.A(G8), .B(new_n1018), .C1(new_n1021), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT49), .ZN(new_n1028));
  NAND2_X1  g603(.A1(G305), .A2(G1981), .ZN(new_n1029));
  INV_X1    g604(.A(G1981), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n572), .A2(new_n577), .A3(new_n1030), .A4(new_n579), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1028), .B1(new_n1032), .B2(KEYINPUT117), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n1034));
  AOI211_X1 g609(.A(new_n1034), .B(KEYINPUT49), .C1(new_n1029), .C2(new_n1031), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n993), .A2(new_n966), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G8), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1033), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1976), .ZN(new_n1039));
  NOR2_X1   g614(.A1(G288), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT52), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1040), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(G288), .B2(new_n1039), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1042), .A2(new_n1043), .A3(G8), .A4(new_n1036), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1038), .A2(new_n1045), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1027), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1020), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n997), .A2(new_n998), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(G1956), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT56), .B(G2072), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n1009), .B2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g627(.A(G299), .B(KEYINPUT57), .Z(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT123), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1053), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1009), .A2(new_n1051), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1055), .B(new_n1056), .C1(new_n1057), .C2(new_n1050), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT123), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OAI22_X1  g635(.A1(new_n1024), .A2(G1348), .B1(new_n1036), .B2(G2067), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1061), .A2(new_n598), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1054), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  OAI221_X1 g638(.A(KEYINPUT60), .B1(new_n1036), .B2(G2067), .C1(G1348), .C2(new_n1024), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1064), .A2(KEYINPUT126), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1064), .A2(KEYINPUT126), .A3(new_n597), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n597), .B1(new_n1064), .B2(KEYINPUT126), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1065), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT60), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1061), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT61), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1054), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT125), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1054), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1052), .A2(KEYINPUT125), .A3(new_n1053), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(KEYINPUT61), .A3(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1071), .B(new_n1075), .C1(new_n1079), .C2(new_n1060), .ZN(new_n1080));
  INV_X1    g655(.A(G1996), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1009), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT124), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1009), .A2(KEYINPUT124), .A3(new_n1081), .ZN(new_n1085));
  XOR2_X1   g660(.A(KEYINPUT58), .B(G1341), .Z(new_n1086));
  NAND2_X1  g661(.A1(new_n1036), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n543), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(new_n1088), .B2(new_n543), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1063), .B1(new_n1080), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT127), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1024), .A2(new_n790), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1024), .A2(KEYINPUT120), .A3(new_n790), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n965), .B1(new_n1002), .B2(KEYINPUT45), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n993), .B2(KEYINPUT45), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n744), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1097), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1094), .B1(new_n1102), .B2(G8), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT51), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1102), .A2(G286), .ZN(new_n1106));
  OAI21_X1  g681(.A(G8), .B1(new_n1102), .B2(G286), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI221_X1 g683(.A(G8), .B1(G286), .B2(new_n1102), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT53), .B1(new_n1009), .B2(new_n782), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(new_n759), .B2(new_n1025), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n782), .A2(KEYINPUT53), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1112), .B1(new_n1100), .B2(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(G171), .B(KEYINPUT54), .Z(new_n1115));
  NOR3_X1   g690(.A1(new_n964), .A2(new_n965), .A3(new_n1113), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1114), .A2(new_n1115), .B1(new_n1112), .B2(new_n1118), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1110), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1093), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1110), .A2(KEYINPUT62), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1108), .A2(new_n1123), .A3(new_n1109), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1122), .A2(G171), .A3(new_n1124), .A4(new_n1114), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1048), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n1127));
  INV_X1    g702(.A(G8), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1128), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1018), .B1(new_n1129), .B2(new_n1013), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1027), .A2(new_n1046), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1102), .A2(G8), .A3(G168), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1127), .B1(new_n1133), .B2(KEYINPUT63), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT63), .ZN(new_n1135));
  OAI211_X1 g710(.A(KEYINPUT121), .B(new_n1135), .C1(new_n1048), .C2(new_n1132), .ZN(new_n1136));
  OAI21_X1  g711(.A(G8), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1137));
  AOI211_X1 g712(.A(new_n1135), .B(new_n1132), .C1(new_n1019), .C2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1047), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1134), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1140));
  OR3_X1    g715(.A1(new_n1038), .A2(G1976), .A3(G288), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1037), .B1(new_n1141), .B2(new_n1031), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1027), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1143), .B2(new_n1046), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1140), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT122), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1140), .A2(new_n1147), .A3(new_n1144), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1126), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n984), .A2(KEYINPUT112), .ZN(new_n1150));
  NAND2_X1  g725(.A1(G290), .A2(G1986), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n1150), .B(new_n1151), .Z(new_n1152));
  NOR2_X1   g727(.A1(new_n1152), .A2(new_n967), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n1153), .B(KEYINPUT113), .Z(new_n1154));
  NAND4_X1  g729(.A1(new_n1154), .A2(new_n983), .A3(new_n973), .A4(new_n971), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n988), .B1(new_n1149), .B2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g731(.A1(new_n874), .A2(new_n876), .ZN(new_n1158));
  NOR4_X1   g732(.A1(G229), .A2(new_n458), .A3(G401), .A4(G227), .ZN(new_n1159));
  NAND3_X1  g733(.A1(new_n1158), .A2(new_n956), .A3(new_n1159), .ZN(G225));
  INV_X1    g734(.A(G225), .ZN(G308));
endmodule


