//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT73), .ZN(new_n203));
  AND2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G155gat), .ZN(new_n207));
  INV_X1    g006(.A(G162gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(KEYINPUT73), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(KEYINPUT2), .ZN(new_n213));
  INV_X1    g012(.A(G141gat), .ZN(new_n214));
  INV_X1    g013(.A(G148gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n213), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n212), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT74), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT74), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n212), .A2(new_n221), .A3(new_n218), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT75), .B(G162gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G155gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT2), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n216), .A2(new_n217), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n210), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n220), .A2(new_n222), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n230));
  INV_X1    g029(.A(G113gat), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n231), .A2(G120gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(G120gat), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT1), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G127gat), .B(G134gat), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n230), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n234), .A2(new_n230), .A3(new_n235), .ZN(new_n238));
  NOR2_X1   g037(.A1(G127gat), .A2(G134gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(KEYINPUT66), .B(G127gat), .Z(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G134gat), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n237), .A2(new_n238), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT79), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n229), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n225), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n212), .A2(new_n221), .A3(new_n218), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n221), .B1(new_n212), .B2(new_n218), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OR2_X1    g048(.A1(G127gat), .A2(G134gat), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n232), .A2(new_n233), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n242), .B(new_n250), .C1(new_n251), .C2(KEYINPUT1), .ZN(new_n252));
  INV_X1    g051(.A(new_n238), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(new_n253), .B2(new_n236), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT79), .B1(new_n249), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n245), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT76), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n249), .A2(new_n257), .ZN(new_n258));
  OAI211_X1 g057(.A(KEYINPUT76), .B(new_n246), .C1(new_n247), .C2(new_n248), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n259), .A3(new_n254), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT80), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT80), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n258), .A2(new_n259), .A3(new_n262), .A4(new_n254), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n256), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G225gat), .A2(G233gat), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT5), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT81), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT81), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n268), .B(KEYINPUT5), .C1(new_n264), .C2(new_n265), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n256), .A2(KEYINPUT4), .ZN(new_n271));
  INV_X1    g070(.A(new_n265), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n229), .A2(new_n243), .A3(KEYINPUT4), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n259), .A3(KEYINPUT3), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT77), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n258), .A2(new_n259), .A3(KEYINPUT77), .A4(KEYINPUT3), .ZN(new_n278));
  XOR2_X1   g077(.A(KEYINPUT78), .B(KEYINPUT3), .Z(new_n279));
  AOI21_X1  g078(.A(new_n243), .B1(new_n229), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n274), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n270), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT4), .B1(new_n229), .B2(new_n243), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n284), .B1(new_n256), .B2(KEYINPUT4), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n272), .A2(KEYINPUT5), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT82), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G1gat), .B(G29gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT0), .ZN(new_n291));
  XNOR2_X1  g090(.A(G57gat), .B(G85gat), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n291), .B(new_n292), .Z(new_n293));
  NAND3_X1  g092(.A1(new_n283), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n293), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n267), .A2(new_n269), .B1(new_n281), .B2(new_n274), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n295), .B1(new_n296), .B2(new_n288), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n294), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n289), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n300), .A2(KEYINPUT88), .A3(KEYINPUT6), .A4(new_n295), .ZN(new_n301));
  INV_X1    g100(.A(G226gat), .ZN(new_n302));
  INV_X1    g101(.A(G233gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT23), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(G169gat), .B2(G176gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT24), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(G183gat), .A3(G190gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT24), .ZN(new_n311));
  NOR2_X1   g110(.A1(G183gat), .A2(G190gat), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n307), .B(new_n309), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT64), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT25), .ZN(new_n316));
  NAND2_X1  g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(G169gat), .A2(G176gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n317), .B1(new_n319), .B2(new_n306), .ZN(new_n320));
  OAI22_X1  g119(.A1(new_n315), .A2(new_n316), .B1(new_n313), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n313), .ZN(new_n322));
  INV_X1    g121(.A(new_n320), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n322), .A2(new_n323), .A3(new_n314), .A4(KEYINPUT25), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT28), .ZN(new_n325));
  INV_X1    g124(.A(G183gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT27), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT65), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G190gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT27), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G183gat), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n328), .B1(new_n327), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n325), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n327), .A2(new_n333), .A3(KEYINPUT28), .A4(new_n330), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT26), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n310), .B1(new_n319), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n318), .A2(KEYINPUT26), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n339), .B1(new_n317), .B2(new_n340), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n321), .A2(new_n324), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n305), .B1(new_n342), .B2(KEYINPUT29), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n333), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT65), .ZN(new_n345));
  AOI21_X1  g144(.A(G190gat), .B1(new_n327), .B2(new_n328), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT28), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n336), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n341), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n326), .A2(new_n330), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n350), .A2(KEYINPUT24), .A3(new_n310), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n351), .A2(KEYINPUT64), .A3(new_n307), .A4(new_n309), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n322), .A2(new_n323), .B1(new_n352), .B2(KEYINPUT25), .ZN(new_n353));
  NOR4_X1   g152(.A1(new_n313), .A2(new_n320), .A3(KEYINPUT64), .A4(new_n316), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n349), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n304), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n343), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT71), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n359));
  OR2_X1    g158(.A1(new_n359), .A2(KEYINPUT69), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(KEYINPUT69), .ZN(new_n361));
  INV_X1    g160(.A(G197gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G204gat), .ZN(new_n363));
  INV_X1    g162(.A(G204gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G197gat), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n360), .A2(new_n361), .A3(new_n363), .A4(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT70), .ZN(new_n367));
  XNOR2_X1  g166(.A(G211gat), .B(G218gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n368), .B1(new_n366), .B2(new_n367), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n358), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n371), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(KEYINPUT71), .A3(new_n369), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n357), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT72), .ZN(new_n378));
  NOR3_X1   g177(.A1(new_n342), .A2(new_n378), .A3(new_n305), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT72), .B1(new_n355), .B2(new_n304), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n343), .B(new_n375), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G8gat), .B(G36gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G64gat), .B(G92gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n383), .B(new_n384), .Z(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT87), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT37), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n382), .B2(new_n386), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT38), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT29), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n304), .B1(new_n355), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n356), .A2(new_n378), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n355), .A2(KEYINPUT72), .A3(new_n304), .ZN(new_n396));
  AOI211_X1 g195(.A(new_n375), .B(new_n394), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n342), .A2(new_n305), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n375), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT37), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n392), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n388), .B1(new_n391), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n389), .B1(new_n357), .B2(new_n375), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n343), .B(new_n376), .C1(new_n379), .C2(new_n380), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT38), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n385), .B1(new_n377), .B2(new_n381), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n405), .B(KEYINPUT87), .C1(new_n406), .C2(new_n390), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n387), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT89), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n389), .B1(new_n377), .B2(new_n381), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n409), .B(KEYINPUT38), .C1(new_n391), .C2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT38), .B1(new_n391), .B2(new_n410), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT89), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n408), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(KEYINPUT6), .B(new_n295), .C1(new_n296), .C2(new_n288), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT88), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n299), .A2(new_n301), .A3(new_n414), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n281), .A2(new_n285), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT39), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n420), .A3(new_n272), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n264), .A2(new_n265), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT39), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n265), .B1(new_n281), .B2(new_n285), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n293), .B(new_n421), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT40), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n295), .B1(new_n424), .B2(new_n420), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT40), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n427), .B(new_n428), .C1(new_n424), .C2(new_n423), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT30), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n406), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(new_n387), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n297), .A3(new_n433), .ZN(new_n434));
  XOR2_X1   g233(.A(G78gat), .B(G106gat), .Z(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT31), .B(G50gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G22gat), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n373), .A2(new_n393), .A3(new_n369), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT84), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT3), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT84), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n373), .A2(new_n442), .A3(new_n393), .A4(new_n369), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n258), .A2(new_n259), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(G228gat), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n447), .A2(new_n303), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT29), .B1(new_n229), .B2(new_n279), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n375), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n446), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT83), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n368), .B(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n393), .B1(new_n453), .B2(new_n366), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n366), .A2(new_n452), .A3(new_n368), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n279), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n249), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n457), .B1(new_n375), .B2(new_n449), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n458), .B1(new_n447), .B2(new_n303), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n438), .B1(new_n451), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n437), .B1(new_n460), .B2(KEYINPUT85), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n448), .B1(new_n375), .B2(new_n449), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n462), .B1(new_n445), .B2(new_n444), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n448), .B1(new_n450), .B2(new_n457), .ZN(new_n464));
  OAI21_X1  g263(.A(G22gat), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n451), .A2(new_n438), .A3(new_n459), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n465), .A2(KEYINPUT85), .A3(new_n466), .A4(new_n437), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n434), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n418), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT36), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n355), .A2(new_n243), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n254), .B(new_n349), .C1(new_n353), .C2(new_n354), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(G227gat), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n478), .A2(new_n303), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT34), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n475), .A2(new_n476), .A3(new_n479), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n484), .A2(KEYINPUT68), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(KEYINPUT68), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT33), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  XOR2_X1   g286(.A(G15gat), .B(G43gat), .Z(new_n488));
  XNOR2_X1  g287(.A(G71gat), .B(G99gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n483), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n481), .B(KEYINPUT34), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT33), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n484), .A2(KEYINPUT68), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n484), .A2(KEYINPUT68), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n493), .A2(new_n497), .A3(new_n490), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n485), .A2(new_n486), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT32), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n492), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n501), .B1(new_n492), .B2(new_n498), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n474), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n492), .A2(new_n498), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n500), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n492), .A2(new_n498), .A3(new_n501), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n506), .A2(KEYINPUT36), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n433), .B1(new_n299), .B2(new_n415), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT86), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n470), .B(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n509), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n473), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n506), .A2(new_n469), .A3(new_n468), .A4(new_n507), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n299), .A2(new_n301), .A3(new_n417), .ZN(new_n518));
  INV_X1    g317(.A(new_n433), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT35), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n468), .A2(new_n520), .A3(new_n469), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n506), .A2(KEYINPUT90), .A3(new_n507), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT90), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(new_n502), .B2(new_n503), .ZN(new_n524));
  AND4_X1   g323(.A1(new_n519), .A2(new_n521), .A3(new_n522), .A4(new_n524), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n517), .A2(KEYINPUT35), .B1(new_n518), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n202), .B1(new_n514), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n470), .B(KEYINPUT86), .ZN(new_n528));
  INV_X1    g327(.A(new_n415), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT6), .B1(new_n300), .B2(new_n295), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(new_n294), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n528), .B1(new_n531), .B2(new_n433), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n418), .A2(new_n472), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n533), .A3(new_n509), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n525), .A2(new_n518), .ZN(new_n535));
  AOI211_X1 g334(.A(new_n433), .B(new_n515), .C1(new_n299), .C2(new_n415), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(new_n520), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n537), .A3(KEYINPUT91), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n527), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT97), .ZN(new_n540));
  XNOR2_X1  g339(.A(G15gat), .B(G22gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT16), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n541), .B1(new_n542), .B2(G1gat), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(G1gat), .B2(new_n541), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(G8gat), .ZN(new_n545));
  INV_X1    g344(.A(G50gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(G43gat), .ZN(new_n547));
  INV_X1    g346(.A(G43gat), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n548), .A2(G50gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT15), .ZN(new_n550));
  NOR3_X1   g349(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n551), .B1(G29gat), .B2(G36gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(KEYINPUT93), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT93), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n554), .B1(new_n548), .B2(G50gat), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n553), .B(new_n555), .C1(G43gat), .C2(new_n546), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(new_n550), .ZN(new_n557));
  INV_X1    g356(.A(G29gat), .ZN(new_n558));
  INV_X1    g357(.A(G36gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n559), .A3(KEYINPUT14), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT14), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(G29gat), .B2(G36gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n552), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(KEYINPUT92), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT92), .ZN(new_n567));
  OAI22_X1  g366(.A1(new_n563), .A2(new_n567), .B1(new_n558), .B2(new_n559), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n551), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n545), .A2(new_n570), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n571), .A2(KEYINPUT94), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(KEYINPUT94), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n570), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n575), .A2(KEYINPUT17), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n544), .B(G8gat), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(KEYINPUT17), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n574), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT18), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n574), .A2(new_n579), .A3(KEYINPUT18), .A4(new_n580), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT95), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n574), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n572), .A2(KEYINPUT95), .A3(new_n573), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n586), .A2(new_n587), .B1(new_n575), .B2(new_n577), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n580), .B(KEYINPUT13), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n583), .B(new_n584), .C1(new_n588), .C2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G113gat), .B(G141gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(new_n362), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT11), .B(G169gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT12), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT96), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n596), .B1(new_n583), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n591), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n591), .A2(new_n598), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n540), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n591), .A2(new_n598), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n591), .A2(new_n598), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(KEYINPUT97), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n606));
  INV_X1    g405(.A(G57gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(G64gat), .ZN(new_n608));
  INV_X1    g407(.A(G64gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(G57gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n606), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n613), .B1(new_n612), .B2(new_n611), .ZN(new_n614));
  XOR2_X1   g413(.A(G71gat), .B(G78gat), .Z(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n606), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n608), .A2(KEYINPUT99), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n608), .A2(KEYINPUT99), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n610), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n617), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n623), .A2(KEYINPUT21), .ZN(new_n624));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G127gat), .B(G155gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT20), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n626), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G183gat), .B(G211gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n545), .B1(new_n623), .B2(KEYINPUT21), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G85gat), .A2(G92gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  NAND2_X1  g439(.A1(G99gat), .A2(G106gat), .ZN(new_n641));
  INV_X1    g440(.A(G85gat), .ZN(new_n642));
  INV_X1    g441(.A(G92gat), .ZN(new_n643));
  AOI22_X1  g442(.A1(KEYINPUT8), .A2(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(G99gat), .B(G106gat), .Z(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n646), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n640), .A2(new_n648), .A3(new_n644), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n576), .A2(new_n578), .A3(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(G232gat), .A2(G233gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(KEYINPUT41), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n651), .B(new_n653), .C1(new_n575), .C2(new_n650), .ZN(new_n654));
  XNOR2_X1  g453(.A(G190gat), .B(G218gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT102), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n654), .B(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n652), .A2(KEYINPUT41), .ZN(new_n658));
  XNOR2_X1  g457(.A(G134gat), .B(G162gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n657), .A2(new_n660), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n637), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G120gat), .B(G148gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(G176gat), .B(G204gat), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n665), .B(new_n666), .Z(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(G230gat), .A2(G233gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT104), .Z(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n622), .A2(new_n650), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n616), .A2(new_n647), .A3(new_n621), .A4(new_n649), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n672), .A2(KEYINPUT103), .A3(new_n673), .ZN(new_n674));
  OR3_X1    g473(.A1(new_n622), .A2(new_n650), .A3(KEYINPUT103), .ZN(new_n675));
  AOI21_X1  g474(.A(KEYINPUT10), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT10), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n671), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT105), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n681), .B(new_n671), .C1(new_n676), .C2(new_n678), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n674), .A2(new_n675), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n671), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n668), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n679), .B(new_n667), .C1(new_n671), .C2(new_n684), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n664), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n539), .A2(new_n605), .A3(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n531), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g492(.A(KEYINPUT16), .B(G8gat), .Z(new_n694));
  NAND3_X1  g493(.A1(new_n691), .A2(new_n433), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT42), .ZN(new_n696));
  OAI21_X1  g495(.A(G8gat), .B1(new_n690), .B2(new_n519), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n697), .A2(KEYINPUT106), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(KEYINPUT106), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n696), .A2(new_n698), .A3(new_n699), .ZN(G1325gat));
  OAI21_X1  g499(.A(G15gat), .B1(new_n690), .B2(new_n509), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n524), .A2(new_n522), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n702), .A2(G15gat), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(new_n690), .B2(new_n703), .ZN(G1326gat));
  NAND3_X1  g503(.A1(new_n691), .A2(KEYINPUT107), .A3(new_n528), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n690), .B2(new_n512), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT43), .B(G22gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n663), .A2(new_n711), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n534), .A2(KEYINPUT91), .A3(new_n537), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT91), .B1(new_n534), .B2(new_n537), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n534), .A2(new_n537), .ZN(new_n716));
  INV_X1    g515(.A(new_n663), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n711), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n602), .A2(new_n603), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n637), .A2(new_n721), .A3(new_n688), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n715), .A2(new_n531), .A3(new_n719), .A4(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT44), .B1(new_n716), .B2(new_n717), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n726), .B1(new_n539), .B2(new_n712), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n727), .A2(KEYINPUT108), .A3(new_n531), .A4(new_n722), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n725), .A2(new_n728), .A3(G29gat), .ZN(new_n729));
  INV_X1    g528(.A(new_n637), .ZN(new_n730));
  INV_X1    g529(.A(new_n688), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(new_n717), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n605), .B(new_n733), .C1(new_n713), .C2(new_n714), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n531), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(G29gat), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT45), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n739));
  NOR4_X1   g538(.A1(new_n734), .A2(new_n739), .A3(G29gat), .A4(new_n736), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n729), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n741), .A3(KEYINPUT109), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(G1328gat));
  NAND2_X1  g545(.A1(new_n433), .A2(new_n559), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT46), .B1(new_n734), .B2(new_n747), .ZN(new_n748));
  OR3_X1    g547(.A1(new_n734), .A2(KEYINPUT46), .A3(new_n747), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n727), .A2(new_n433), .A3(new_n722), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n748), .B(new_n749), .C1(new_n750), .C2(new_n559), .ZN(G1329gat));
  INV_X1    g550(.A(new_n702), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n735), .A2(new_n548), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n509), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n727), .A2(new_n754), .A3(new_n722), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G43gat), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n755), .A2(new_n756), .ZN(new_n759));
  OAI211_X1 g558(.A(KEYINPUT47), .B(new_n753), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n755), .A2(G43gat), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n753), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT47), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n760), .A2(new_n764), .ZN(G1330gat));
  INV_X1    g564(.A(KEYINPUT48), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n715), .A2(new_n470), .A3(new_n719), .A4(new_n722), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G50gat), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n512), .A2(G50gat), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n735), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n766), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n769), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n766), .B1(new_n734), .B2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n715), .A2(new_n528), .A3(new_n719), .A4(new_n722), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(G50gat), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT111), .B1(new_n771), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(G50gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n767), .A2(G50gat), .B1(new_n735), .B2(new_n769), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n779), .B(new_n780), .C1(new_n766), .C2(new_n781), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n776), .A2(new_n782), .ZN(G1331gat));
  NOR3_X1   g582(.A1(new_n664), .A2(new_n720), .A3(new_n731), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n716), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n531), .ZN(new_n786));
  XNOR2_X1  g585(.A(KEYINPUT112), .B(G57gat), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n786), .B(new_n787), .ZN(G1332gat));
  AND2_X1   g587(.A1(new_n785), .A2(new_n433), .ZN(new_n789));
  NOR2_X1   g588(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n790));
  AND2_X1   g589(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n789), .B2(new_n790), .ZN(G1333gat));
  NAND2_X1  g592(.A1(new_n785), .A2(new_n754), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n702), .A2(G71gat), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n794), .A2(G71gat), .B1(new_n785), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g596(.A1(new_n785), .A2(new_n528), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g598(.A1(new_n637), .A2(new_n720), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n716), .A2(new_n717), .A3(new_n800), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n801), .B(KEYINPUT51), .Z(new_n802));
  NAND4_X1  g601(.A1(new_n802), .A2(new_n642), .A3(new_n531), .A4(new_n688), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n715), .A2(new_n719), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n800), .A2(new_n688), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n804), .A2(new_n736), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n803), .B1(new_n806), .B2(new_n642), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT113), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n803), .B(new_n809), .C1(new_n642), .C2(new_n806), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(G1336gat));
  NAND4_X1  g610(.A1(new_n802), .A2(new_n643), .A3(new_n433), .A4(new_n688), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n804), .A2(new_n519), .A3(new_n805), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n813), .B2(new_n643), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT52), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n812), .B(new_n816), .C1(new_n643), .C2(new_n813), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(G1337gat));
  NOR3_X1   g617(.A1(new_n702), .A2(G99gat), .A3(new_n731), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n805), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n727), .A2(new_n754), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT114), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G99gat), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n822), .A2(KEYINPUT114), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n820), .B1(new_n824), .B2(new_n825), .ZN(G1338gat));
  NOR3_X1   g625(.A1(new_n731), .A2(new_n471), .A3(G106gat), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n802), .A2(new_n827), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n804), .A2(new_n512), .A3(new_n805), .ZN(new_n829));
  INV_X1    g628(.A(G106gat), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT53), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT53), .B1(new_n802), .B2(new_n827), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n727), .A2(new_n470), .A3(new_n821), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(G106gat), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n834), .B1(new_n833), .B2(new_n836), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n832), .B1(new_n837), .B2(new_n838), .ZN(G1339gat));
  NOR2_X1   g638(.A1(new_n676), .A2(new_n678), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n840), .A2(KEYINPUT116), .A3(new_n670), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT116), .B1(new_n840), .B2(new_n670), .ZN(new_n842));
  OAI211_X1 g641(.A(KEYINPUT54), .B(new_n679), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n680), .A2(new_n844), .A3(new_n682), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n845), .A2(KEYINPUT117), .A3(new_n668), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT117), .B1(new_n845), .B2(new_n668), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n843), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT55), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n843), .B(KEYINPUT55), .C1(new_n846), .C2(new_n847), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n850), .A2(new_n720), .A3(new_n687), .A4(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n596), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n580), .B1(new_n574), .B2(new_n579), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(new_n590), .B2(new_n588), .ZN(new_n855));
  INV_X1    g654(.A(new_n595), .ZN(new_n856));
  OAI22_X1  g655(.A1(new_n591), .A2(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n731), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n717), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n850), .A2(new_n687), .A3(new_n851), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n860), .A2(new_n663), .A3(new_n857), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n730), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n689), .A2(new_n721), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n736), .A2(new_n433), .A3(new_n702), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n862), .A2(KEYINPUT118), .A3(new_n863), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n866), .A2(new_n867), .A3(new_n512), .A4(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n605), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n872), .A3(G113gat), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n872), .B1(new_n871), .B2(G113gat), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n862), .A2(KEYINPUT118), .A3(new_n863), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT118), .B1(new_n862), .B2(new_n863), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n736), .A2(new_n433), .A3(new_n515), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n720), .A2(new_n231), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT120), .ZN(new_n882));
  OAI22_X1  g681(.A1(new_n874), .A2(new_n875), .B1(new_n880), .B2(new_n882), .ZN(G1340gat));
  OAI21_X1  g682(.A(G120gat), .B1(new_n869), .B2(new_n731), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n731), .A2(G120gat), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT121), .Z(G1341gat));
  OAI21_X1  g686(.A(new_n241), .B1(new_n869), .B2(new_n730), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n730), .A2(new_n241), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n880), .B2(new_n889), .ZN(G1342gat));
  OAI21_X1  g689(.A(G134gat), .B1(new_n869), .B2(new_n663), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n663), .A2(G134gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n878), .A2(new_n879), .A3(new_n892), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n893), .A2(KEYINPUT122), .A3(KEYINPUT56), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT122), .B1(new_n893), .B2(KEYINPUT56), .ZN(new_n895));
  OAI221_X1 g694(.A(new_n891), .B1(KEYINPUT56), .B2(new_n893), .C1(new_n894), .C2(new_n895), .ZN(G1343gat));
  NOR3_X1   g695(.A1(new_n736), .A2(new_n433), .A3(new_n754), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n878), .A2(new_n470), .A3(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n870), .A2(G141gat), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT58), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n866), .A2(new_n470), .A3(new_n868), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n605), .A2(new_n850), .A3(new_n687), .A4(new_n851), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n717), .B1(new_n904), .B2(new_n858), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n730), .B1(new_n905), .B2(new_n861), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n863), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n512), .A2(new_n903), .ZN(new_n908));
  AOI22_X1  g707(.A1(new_n902), .A2(new_n903), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n897), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n909), .A2(new_n870), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n901), .B1(new_n911), .B2(new_n214), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT57), .B1(new_n878), .B2(new_n470), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n907), .A2(new_n908), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n720), .B(new_n897), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n915), .A2(G141gat), .B1(new_n899), .B2(new_n900), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT58), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n912), .B1(new_n916), .B2(new_n917), .ZN(G1344gat));
  NAND2_X1  g717(.A1(new_n897), .A2(new_n688), .ZN(new_n919));
  OR3_X1    g718(.A1(new_n902), .A2(G148gat), .A3(new_n919), .ZN(new_n920));
  XNOR2_X1  g719(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n689), .A2(new_n870), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n528), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n903), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n471), .A2(new_n903), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n866), .A2(new_n868), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n919), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n215), .B1(new_n928), .B2(KEYINPUT124), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n878), .A2(new_n926), .B1(new_n903), .B2(new_n924), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(new_n919), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n921), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n215), .A2(KEYINPUT59), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n909), .A2(new_n910), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n935), .B2(new_n688), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n920), .B1(new_n933), .B2(new_n936), .ZN(G1345gat));
  AOI21_X1  g736(.A(G155gat), .B1(new_n899), .B2(new_n637), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n730), .A2(new_n207), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n935), .B2(new_n939), .ZN(G1346gat));
  INV_X1    g739(.A(new_n223), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n899), .A2(new_n941), .A3(new_n717), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n909), .A2(new_n663), .A3(new_n910), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(new_n941), .ZN(G1347gat));
  NOR3_X1   g743(.A1(new_n876), .A2(new_n877), .A3(new_n531), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n433), .A3(new_n516), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n721), .A2(G169gat), .ZN(new_n947));
  OR3_X1    g746(.A1(new_n946), .A2(KEYINPUT125), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(KEYINPUT125), .B1(new_n946), .B2(new_n947), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n531), .A2(new_n519), .A3(new_n702), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n878), .A2(new_n512), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(G169gat), .B1(new_n952), .B2(new_n870), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n953), .A2(KEYINPUT126), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(KEYINPUT126), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n950), .A2(new_n954), .A3(new_n955), .ZN(G1348gat));
  OAI21_X1  g755(.A(G176gat), .B1(new_n952), .B2(new_n731), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n731), .A2(G176gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n957), .B1(new_n946), .B2(new_n958), .ZN(G1349gat));
  OAI21_X1  g758(.A(G183gat), .B1(new_n952), .B2(new_n730), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n730), .A2(new_n344), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n960), .B1(new_n946), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT60), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT60), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n960), .B(new_n965), .C1(new_n946), .C2(new_n962), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1350gat));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n952), .A2(new_n663), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(G190gat), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n968), .B(G190gat), .C1(new_n952), .C2(new_n663), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n717), .A2(new_n330), .ZN(new_n973));
  OAI22_X1  g772(.A1(new_n970), .A2(new_n972), .B1(new_n946), .B2(new_n973), .ZN(G1351gat));
  NOR3_X1   g773(.A1(new_n754), .A2(new_n519), .A3(new_n471), .ZN(new_n975));
  AND4_X1   g774(.A1(new_n362), .A2(new_n945), .A3(new_n720), .A4(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT127), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n925), .A2(new_n927), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n531), .A2(new_n754), .A3(new_n519), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(G197gat), .B1(new_n981), .B2(new_n870), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n978), .A2(new_n982), .ZN(G1352gat));
  OAI21_X1  g782(.A(G204gat), .B1(new_n981), .B2(new_n731), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n945), .A2(new_n975), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n688), .A2(new_n364), .ZN(new_n986));
  OR3_X1    g785(.A1(new_n985), .A2(KEYINPUT62), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g786(.A(KEYINPUT62), .B1(new_n985), .B2(new_n986), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n984), .A2(new_n987), .A3(new_n988), .ZN(G1353gat));
  OR3_X1    g788(.A1(new_n985), .A2(G211gat), .A3(new_n730), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n979), .A2(new_n637), .A3(new_n980), .ZN(new_n991));
  AND3_X1   g790(.A1(new_n991), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n992));
  AOI21_X1  g791(.A(KEYINPUT63), .B1(new_n991), .B2(G211gat), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(G1354gat));
  OAI21_X1  g793(.A(G218gat), .B1(new_n981), .B2(new_n663), .ZN(new_n995));
  OR3_X1    g794(.A1(new_n985), .A2(G218gat), .A3(new_n663), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(G1355gat));
endmodule


