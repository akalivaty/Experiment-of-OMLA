

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X2 U321 ( .A(n385), .B(KEYINPUT41), .ZN(n578) );
  XNOR2_X2 U322 ( .A(n493), .B(KEYINPUT64), .ZN(n385) );
  NOR2_X1 U323 ( .A1(n408), .A2(n582), .ZN(n410) );
  XNOR2_X1 U324 ( .A(n366), .B(G64GAT), .ZN(n428) );
  XNOR2_X1 U325 ( .A(n434), .B(KEYINPUT54), .ZN(n436) );
  XNOR2_X1 U326 ( .A(n334), .B(n424), .ZN(n336) );
  NOR2_X1 U327 ( .A1(n544), .A2(n465), .ZN(n579) );
  XNOR2_X1 U328 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U329 ( .A(KEYINPUT79), .B(n569), .Z(n554) );
  NAND2_X1 U330 ( .A1(n493), .A2(n415), .ZN(n289) );
  AND2_X1 U331 ( .A1(G232GAT), .A2(G233GAT), .ZN(n290) );
  INV_X1 U332 ( .A(KEYINPUT106), .ZN(n409) );
  XNOR2_X1 U333 ( .A(n410), .B(n409), .ZN(n411) );
  NOR2_X1 U334 ( .A1(n416), .A2(n289), .ZN(n417) );
  INV_X1 U335 ( .A(G92GAT), .ZN(n367) );
  XNOR2_X1 U336 ( .A(n328), .B(n290), .ZN(n334) );
  XNOR2_X1 U337 ( .A(n428), .B(n367), .ZN(n369) );
  INV_X2 U338 ( .A(G204GAT), .ZN(n366) );
  XNOR2_X1 U339 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U340 ( .A(n378), .B(n377), .ZN(n379) );
  NOR2_X1 U341 ( .A1(n560), .A2(n463), .ZN(n472) );
  XOR2_X1 U342 ( .A(KEYINPUT36), .B(n554), .Z(n506) );
  XNOR2_X1 U343 ( .A(n460), .B(G218GAT), .ZN(n461) );
  XNOR2_X1 U344 ( .A(n469), .B(n366), .ZN(n470) );
  XNOR2_X1 U345 ( .A(n462), .B(n461), .ZN(G1355GAT) );
  XNOR2_X1 U346 ( .A(n471), .B(n470), .ZN(G1353GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT91), .B(G204GAT), .Z(n292) );
  XNOR2_X1 U348 ( .A(KEYINPUT22), .B(KEYINPUT89), .ZN(n291) );
  XNOR2_X1 U349 ( .A(n292), .B(n291), .ZN(n309) );
  XOR2_X1 U350 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n294) );
  XNOR2_X1 U351 ( .A(KEYINPUT23), .B(KEYINPUT88), .ZN(n293) );
  XNOR2_X1 U352 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U353 ( .A(n295), .B(G106GAT), .Z(n297) );
  XOR2_X1 U354 ( .A(G22GAT), .B(G155GAT), .Z(n400) );
  XNOR2_X1 U355 ( .A(n400), .B(G218GAT), .ZN(n296) );
  XNOR2_X1 U356 ( .A(n297), .B(n296), .ZN(n302) );
  XOR2_X1 U357 ( .A(G50GAT), .B(G162GAT), .Z(n339) );
  XNOR2_X1 U358 ( .A(G78GAT), .B(KEYINPUT74), .ZN(n298) );
  XNOR2_X1 U359 ( .A(n298), .B(G148GAT), .ZN(n382) );
  XOR2_X1 U360 ( .A(n339), .B(n382), .Z(n300) );
  NAND2_X1 U361 ( .A1(G228GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U362 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U363 ( .A(n302), .B(n301), .Z(n307) );
  XNOR2_X1 U364 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n303) );
  XNOR2_X1 U365 ( .A(n303), .B(G211GAT), .ZN(n422) );
  XOR2_X1 U366 ( .A(KEYINPUT90), .B(KEYINPUT3), .Z(n305) );
  XNOR2_X1 U367 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n304) );
  XNOR2_X1 U368 ( .A(n305), .B(n304), .ZN(n451) );
  XNOR2_X1 U369 ( .A(n422), .B(n451), .ZN(n306) );
  XNOR2_X1 U370 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U371 ( .A(n309), .B(n308), .ZN(n484) );
  XOR2_X1 U372 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n315) );
  XOR2_X1 U373 ( .A(KEYINPUT65), .B(KEYINPUT20), .Z(n311) );
  XNOR2_X1 U374 ( .A(G99GAT), .B(G190GAT), .ZN(n310) );
  XNOR2_X1 U375 ( .A(n311), .B(n310), .ZN(n313) );
  XNOR2_X1 U376 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n312) );
  XNOR2_X1 U377 ( .A(n312), .B(KEYINPUT83), .ZN(n452) );
  XNOR2_X1 U378 ( .A(n313), .B(n452), .ZN(n314) );
  XNOR2_X1 U379 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U380 ( .A(G120GAT), .B(G71GAT), .Z(n374) );
  XOR2_X1 U381 ( .A(G15GAT), .B(G127GAT), .Z(n399) );
  XOR2_X1 U382 ( .A(n374), .B(n399), .Z(n317) );
  NAND2_X1 U383 ( .A1(G227GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U384 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U385 ( .A(n319), .B(n318), .Z(n326) );
  XOR2_X1 U386 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n321) );
  XNOR2_X1 U387 ( .A(KEYINPUT19), .B(KEYINPUT86), .ZN(n320) );
  XNOR2_X1 U388 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U389 ( .A(n322), .B(G183GAT), .Z(n324) );
  XNOR2_X1 U390 ( .A(G169GAT), .B(G176GAT), .ZN(n323) );
  XNOR2_X1 U391 ( .A(n324), .B(n323), .ZN(n423) );
  XOR2_X1 U392 ( .A(G43GAT), .B(G134GAT), .Z(n328) );
  XNOR2_X1 U393 ( .A(n423), .B(n328), .ZN(n325) );
  XNOR2_X1 U394 ( .A(n326), .B(n325), .ZN(n544) );
  NAND2_X1 U395 ( .A1(n484), .A2(n544), .ZN(n327) );
  XNOR2_X1 U396 ( .A(n327), .B(KEYINPUT26), .ZN(n560) );
  INV_X1 U397 ( .A(G218GAT), .ZN(n329) );
  NAND2_X1 U398 ( .A1(G92GAT), .A2(n329), .ZN(n331) );
  NAND2_X1 U399 ( .A1(n367), .A2(G218GAT), .ZN(n330) );
  NAND2_X1 U400 ( .A1(n331), .A2(n330), .ZN(n333) );
  XNOR2_X1 U401 ( .A(G36GAT), .B(G190GAT), .ZN(n332) );
  XNOR2_X1 U402 ( .A(n333), .B(n332), .ZN(n424) );
  INV_X1 U403 ( .A(KEYINPUT66), .ZN(n335) );
  XNOR2_X1 U404 ( .A(n336), .B(n335), .ZN(n343) );
  XOR2_X1 U405 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n338) );
  XNOR2_X1 U406 ( .A(KEYINPUT78), .B(KEYINPUT77), .ZN(n337) );
  XOR2_X1 U407 ( .A(n338), .B(n337), .Z(n341) );
  XNOR2_X1 U408 ( .A(n339), .B(KEYINPUT10), .ZN(n340) );
  XNOR2_X1 U409 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n344) );
  XNOR2_X1 U410 ( .A(n344), .B(KEYINPUT7), .ZN(n361) );
  XNOR2_X1 U411 ( .A(G99GAT), .B(G106GAT), .ZN(n345) );
  XNOR2_X1 U412 ( .A(n345), .B(G85GAT), .ZN(n381) );
  XNOR2_X1 U413 ( .A(n361), .B(n381), .ZN(n346) );
  XNOR2_X1 U414 ( .A(n347), .B(n346), .ZN(n569) );
  XOR2_X1 U415 ( .A(KEYINPUT105), .B(KEYINPUT46), .Z(n387) );
  XOR2_X1 U416 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n349) );
  XNOR2_X1 U417 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n348) );
  XNOR2_X1 U418 ( .A(n349), .B(n348), .ZN(n357) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n355) );
  XOR2_X1 U420 ( .A(G141GAT), .B(G197GAT), .Z(n351) );
  XNOR2_X1 U421 ( .A(G50GAT), .B(G22GAT), .ZN(n350) );
  XNOR2_X1 U422 ( .A(n351), .B(n350), .ZN(n353) );
  XOR2_X1 U423 ( .A(G36GAT), .B(G43GAT), .Z(n352) );
  XNOR2_X1 U424 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U425 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U426 ( .A(n357), .B(n356), .ZN(n365) );
  XOR2_X1 U427 ( .A(KEYINPUT69), .B(G15GAT), .Z(n359) );
  XNOR2_X1 U428 ( .A(G169GAT), .B(G113GAT), .ZN(n358) );
  XNOR2_X1 U429 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U430 ( .A(n361), .B(n360), .ZN(n363) );
  XOR2_X1 U431 ( .A(G1GAT), .B(KEYINPUT70), .Z(n362) );
  XNOR2_X1 U432 ( .A(G8GAT), .B(n362), .ZN(n394) );
  XNOR2_X1 U433 ( .A(n363), .B(n394), .ZN(n364) );
  XNOR2_X1 U434 ( .A(n365), .B(n364), .ZN(n573) );
  XOR2_X2 U435 ( .A(G57GAT), .B(KEYINPUT13), .Z(n401) );
  XNOR2_X1 U436 ( .A(G176GAT), .B(n401), .ZN(n368) );
  XNOR2_X1 U437 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U438 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n371) );
  NAND2_X1 U439 ( .A1(G230GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U440 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n373), .B(n372), .ZN(n380) );
  XOR2_X1 U442 ( .A(n374), .B(KEYINPUT33), .Z(n378) );
  XOR2_X1 U443 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n376) );
  XNOR2_X1 U444 ( .A(KEYINPUT75), .B(KEYINPUT31), .ZN(n375) );
  XOR2_X1 U445 ( .A(n376), .B(n375), .Z(n377) );
  XNOR2_X1 U446 ( .A(n380), .B(n379), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X2 U448 ( .A(n384), .B(n383), .ZN(n493) );
  NAND2_X1 U449 ( .A1(n573), .A2(n578), .ZN(n386) );
  XOR2_X1 U450 ( .A(n387), .B(n386), .Z(n408) );
  XOR2_X1 U451 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n389) );
  XNOR2_X1 U452 ( .A(G183GAT), .B(G71GAT), .ZN(n388) );
  XNOR2_X1 U453 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U454 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n391) );
  XNOR2_X1 U455 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n390) );
  XNOR2_X1 U456 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n407) );
  INV_X1 U458 ( .A(n394), .ZN(n395) );
  XOR2_X1 U459 ( .A(n395), .B(KEYINPUT14), .Z(n397) );
  NAND2_X1 U460 ( .A1(G231GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U461 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U462 ( .A(n399), .B(n398), .ZN(n405) );
  XOR2_X1 U463 ( .A(n401), .B(n400), .Z(n403) );
  XNOR2_X1 U464 ( .A(G211GAT), .B(G78GAT), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U466 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n407), .B(n406), .ZN(n503) );
  INV_X1 U468 ( .A(n503), .ZN(n582) );
  NOR2_X1 U469 ( .A1(n569), .A2(n411), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n412), .B(KEYINPUT47), .ZN(n419) );
  INV_X1 U471 ( .A(KEYINPUT45), .ZN(n414) );
  NOR2_X1 U472 ( .A1(n506), .A2(n503), .ZN(n413) );
  XNOR2_X1 U473 ( .A(n414), .B(n413), .ZN(n416) );
  INV_X1 U474 ( .A(n573), .ZN(n415) );
  XNOR2_X1 U475 ( .A(KEYINPUT107), .B(n417), .ZN(n418) );
  NAND2_X1 U476 ( .A1(n419), .A2(n418), .ZN(n421) );
  XNOR2_X1 U477 ( .A(KEYINPUT108), .B(KEYINPUT48), .ZN(n420) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n542) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n432) );
  XOR2_X1 U480 ( .A(n424), .B(KEYINPUT98), .Z(n426) );
  NAND2_X1 U481 ( .A1(G226GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U482 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U483 ( .A(n427), .B(KEYINPUT97), .Z(n430) );
  XNOR2_X1 U484 ( .A(G8GAT), .B(n428), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n533) );
  XNOR2_X1 U487 ( .A(KEYINPUT117), .B(n533), .ZN(n433) );
  NAND2_X1 U488 ( .A1(n542), .A2(n433), .ZN(n434) );
  XNOR2_X1 U489 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n459) );
  NAND2_X1 U491 ( .A1(G225GAT), .A2(G233GAT), .ZN(n442) );
  XOR2_X1 U492 ( .A(G155GAT), .B(G148GAT), .Z(n438) );
  XNOR2_X1 U493 ( .A(G134GAT), .B(G162GAT), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n440) );
  XOR2_X1 U495 ( .A(G29GAT), .B(G85GAT), .Z(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n458) );
  XOR2_X1 U498 ( .A(KEYINPUT6), .B(KEYINPUT93), .Z(n444) );
  XNOR2_X1 U499 ( .A(KEYINPUT96), .B(KEYINPUT4), .ZN(n443) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n456) );
  XOR2_X1 U501 ( .A(KEYINPUT5), .B(G120GAT), .Z(n446) );
  XNOR2_X1 U502 ( .A(G1GAT), .B(G127GAT), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U504 ( .A(KEYINPUT95), .B(G57GAT), .Z(n448) );
  XNOR2_X1 U505 ( .A(KEYINPUT1), .B(KEYINPUT94), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U507 ( .A(n450), .B(n449), .Z(n454) );
  XNOR2_X1 U508 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U509 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U510 ( .A(n456), .B(n455), .Z(n457) );
  XNOR2_X1 U511 ( .A(n458), .B(n457), .ZN(n531) );
  NAND2_X1 U512 ( .A1(n459), .A2(n531), .ZN(n463) );
  XOR2_X1 U513 ( .A(n472), .B(KEYINPUT124), .Z(n468) );
  NOR2_X1 U514 ( .A1(n468), .A2(n506), .ZN(n462) );
  XNOR2_X1 U515 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n460) );
  NOR2_X1 U516 ( .A1(n463), .A2(n484), .ZN(n464) );
  XNOR2_X1 U517 ( .A(n464), .B(KEYINPUT55), .ZN(n465) );
  NAND2_X1 U518 ( .A1(n582), .A2(n579), .ZN(n467) );
  XNOR2_X1 U519 ( .A(G183GAT), .B(KEYINPUT122), .ZN(n466) );
  XNOR2_X1 U520 ( .A(n467), .B(n466), .ZN(G1350GAT) );
  NOR2_X1 U521 ( .A1(n468), .A2(n493), .ZN(n471) );
  XNOR2_X1 U522 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n469) );
  XNOR2_X1 U523 ( .A(n472), .B(KEYINPUT124), .ZN(n583) );
  NAND2_X1 U524 ( .A1(n573), .A2(n583), .ZN(n475) );
  XOR2_X1 U525 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n473) );
  XNOR2_X1 U526 ( .A(n473), .B(G197GAT), .ZN(n474) );
  XNOR2_X1 U527 ( .A(n475), .B(n474), .ZN(G1352GAT) );
  NAND2_X1 U528 ( .A1(n579), .A2(n554), .ZN(n478) );
  XOR2_X1 U529 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n476) );
  XNOR2_X1 U530 ( .A(n476), .B(G190GAT), .ZN(n477) );
  XNOR2_X1 U531 ( .A(n478), .B(n477), .ZN(G1351GAT) );
  XNOR2_X1 U532 ( .A(n533), .B(KEYINPUT27), .ZN(n481) );
  NOR2_X1 U533 ( .A1(n531), .A2(n481), .ZN(n541) );
  XNOR2_X1 U534 ( .A(KEYINPUT28), .B(n484), .ZN(n547) );
  XNOR2_X1 U535 ( .A(KEYINPUT87), .B(n544), .ZN(n479) );
  NOR2_X1 U536 ( .A1(n547), .A2(n479), .ZN(n480) );
  NAND2_X1 U537 ( .A1(n541), .A2(n480), .ZN(n490) );
  NOR2_X1 U538 ( .A1(n560), .A2(n481), .ZN(n482) );
  XNOR2_X1 U539 ( .A(KEYINPUT99), .B(n482), .ZN(n487) );
  NOR2_X1 U540 ( .A1(n544), .A2(n533), .ZN(n483) );
  NOR2_X1 U541 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U542 ( .A(KEYINPUT25), .B(n485), .ZN(n486) );
  NAND2_X1 U543 ( .A1(n487), .A2(n486), .ZN(n488) );
  NAND2_X1 U544 ( .A1(n531), .A2(n488), .ZN(n489) );
  NAND2_X1 U545 ( .A1(n490), .A2(n489), .ZN(n502) );
  OR2_X1 U546 ( .A1(n554), .A2(n503), .ZN(n491) );
  XOR2_X1 U547 ( .A(KEYINPUT16), .B(n491), .Z(n492) );
  AND2_X1 U548 ( .A1(n502), .A2(n492), .ZN(n521) );
  NAND2_X1 U549 ( .A1(n493), .A2(n573), .ZN(n494) );
  XOR2_X1 U550 ( .A(KEYINPUT76), .B(n494), .Z(n508) );
  NAND2_X1 U551 ( .A1(n521), .A2(n508), .ZN(n500) );
  NOR2_X1 U552 ( .A1(n531), .A2(n500), .ZN(n495) );
  XOR2_X1 U553 ( .A(KEYINPUT34), .B(n495), .Z(n496) );
  XNOR2_X1 U554 ( .A(G1GAT), .B(n496), .ZN(G1324GAT) );
  NOR2_X1 U555 ( .A1(n533), .A2(n500), .ZN(n497) );
  XOR2_X1 U556 ( .A(G8GAT), .B(n497), .Z(G1325GAT) );
  NOR2_X1 U557 ( .A1(n544), .A2(n500), .ZN(n499) );
  XNOR2_X1 U558 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(G1326GAT) );
  INV_X1 U560 ( .A(n547), .ZN(n538) );
  NOR2_X1 U561 ( .A1(n538), .A2(n500), .ZN(n501) );
  XOR2_X1 U562 ( .A(G22GAT), .B(n501), .Z(G1327GAT) );
  XNOR2_X1 U563 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n511) );
  NAND2_X1 U564 ( .A1(n503), .A2(n502), .ZN(n504) );
  XNOR2_X1 U565 ( .A(KEYINPUT100), .B(n504), .ZN(n505) );
  NOR2_X1 U566 ( .A1(n506), .A2(n505), .ZN(n507) );
  XOR2_X1 U567 ( .A(KEYINPUT37), .B(n507), .Z(n530) );
  NAND2_X1 U568 ( .A1(n530), .A2(n508), .ZN(n509) );
  XNOR2_X1 U569 ( .A(KEYINPUT38), .B(n509), .ZN(n516) );
  NOR2_X1 U570 ( .A1(n531), .A2(n516), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n511), .B(n510), .ZN(G1328GAT) );
  NOR2_X1 U572 ( .A1(n533), .A2(n516), .ZN(n512) );
  XOR2_X1 U573 ( .A(G36GAT), .B(n512), .Z(G1329GAT) );
  XNOR2_X1 U574 ( .A(KEYINPUT40), .B(KEYINPUT101), .ZN(n514) );
  NOR2_X1 U575 ( .A1(n544), .A2(n516), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U577 ( .A(G43GAT), .B(n515), .ZN(G1330GAT) );
  NOR2_X1 U578 ( .A1(n516), .A2(n538), .ZN(n517) );
  XOR2_X1 U579 ( .A(G50GAT), .B(n517), .Z(G1331GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n519) );
  XNOR2_X1 U581 ( .A(G57GAT), .B(KEYINPUT102), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n519), .B(n518), .ZN(n523) );
  INV_X1 U583 ( .A(n578), .ZN(n520) );
  NOR2_X1 U584 ( .A1(n573), .A2(n520), .ZN(n529) );
  NAND2_X1 U585 ( .A1(n529), .A2(n521), .ZN(n526) );
  NOR2_X1 U586 ( .A1(n531), .A2(n526), .ZN(n522) );
  XOR2_X1 U587 ( .A(n523), .B(n522), .Z(G1332GAT) );
  NOR2_X1 U588 ( .A1(n533), .A2(n526), .ZN(n524) );
  XOR2_X1 U589 ( .A(G64GAT), .B(n524), .Z(G1333GAT) );
  NOR2_X1 U590 ( .A1(n544), .A2(n526), .ZN(n525) );
  XOR2_X1 U591 ( .A(G71GAT), .B(n525), .Z(G1334GAT) );
  NOR2_X1 U592 ( .A1(n538), .A2(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(G1335GAT) );
  NAND2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n537) );
  NOR2_X1 U596 ( .A1(n531), .A2(n537), .ZN(n532) );
  XOR2_X1 U597 ( .A(G85GAT), .B(n532), .Z(G1336GAT) );
  NOR2_X1 U598 ( .A1(n533), .A2(n537), .ZN(n534) );
  XOR2_X1 U599 ( .A(G92GAT), .B(n534), .Z(G1337GAT) );
  NOR2_X1 U600 ( .A1(n544), .A2(n537), .ZN(n535) );
  XOR2_X1 U601 ( .A(KEYINPUT104), .B(n535), .Z(n536) );
  XNOR2_X1 U602 ( .A(G99GAT), .B(n536), .ZN(G1338GAT) );
  NOR2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U604 ( .A(KEYINPUT44), .B(n539), .Z(n540) );
  XNOR2_X1 U605 ( .A(G106GAT), .B(n540), .ZN(G1339GAT) );
  XOR2_X1 U606 ( .A(G113GAT), .B(KEYINPUT111), .Z(n549) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U608 ( .A(KEYINPUT109), .B(n543), .Z(n559) );
  NOR2_X1 U609 ( .A1(n544), .A2(n559), .ZN(n545) );
  XOR2_X1 U610 ( .A(KEYINPUT110), .B(n545), .Z(n546) );
  NOR2_X1 U611 ( .A1(n547), .A2(n546), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n555), .A2(n573), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n549), .B(n548), .ZN(G1340GAT) );
  XOR2_X1 U614 ( .A(G120GAT), .B(KEYINPUT49), .Z(n551) );
  NAND2_X1 U615 ( .A1(n555), .A2(n578), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(G1341GAT) );
  NAND2_X1 U617 ( .A1(n582), .A2(n555), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n552), .B(KEYINPUT50), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G127GAT), .B(n553), .ZN(G1342GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT112), .B(KEYINPUT51), .Z(n557) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G134GAT), .B(n558), .ZN(G1343GAT) );
  XOR2_X1 U624 ( .A(G141GAT), .B(KEYINPUT113), .Z(n562) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n570) );
  NAND2_X1 U626 ( .A1(n570), .A2(n573), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1344GAT) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT114), .ZN(n566) );
  XOR2_X1 U629 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n564) );
  NAND2_X1 U630 ( .A1(n570), .A2(n578), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1345GAT) );
  XOR2_X1 U633 ( .A(G155GAT), .B(KEYINPUT115), .Z(n568) );
  NAND2_X1 U634 ( .A1(n570), .A2(n582), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(G1346GAT) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT116), .ZN(n572) );
  XNOR2_X1 U638 ( .A(G162GAT), .B(n572), .ZN(G1347GAT) );
  NAND2_X1 U639 ( .A1(n573), .A2(n579), .ZN(n574) );
  XNOR2_X1 U640 ( .A(G169GAT), .B(n574), .ZN(G1348GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n576) );
  XNOR2_X1 U642 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U644 ( .A(KEYINPUT56), .B(n577), .Z(n581) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1349GAT) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(KEYINPUT126), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G211GAT), .B(n585), .ZN(G1354GAT) );
endmodule

