//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  AND2_X1   g001(.A1(KEYINPUT68), .A2(G237), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT68), .A2(G237), .ZN(new_n189));
  OAI211_X1 g003(.A(G214), .B(new_n187), .C1(new_n188), .C2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT68), .B(G237), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n193), .A2(G143), .A3(G214), .A4(new_n187), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT18), .A3(G131), .ZN(new_n196));
  INV_X1    g010(.A(G140), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G125), .ZN(new_n198));
  INV_X1    g012(.A(G125), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  XNOR2_X1  g016(.A(G125), .B(G140), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT18), .A2(G131), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n192), .A2(new_n194), .A3(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n196), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT73), .B1(new_n198), .B2(KEYINPUT16), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n198), .A2(new_n200), .A3(KEYINPUT16), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT73), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n212), .A2(new_n213), .A3(new_n197), .A4(G125), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n210), .A2(new_n211), .A3(G146), .A4(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n201), .A2(KEYINPUT19), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT19), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n203), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n218), .A3(new_n204), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT90), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT64), .B(G131), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n192), .A2(new_n194), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n222), .B1(new_n192), .B2(new_n194), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n215), .B(new_n221), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n219), .A2(new_n220), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n209), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G113), .B(G122), .ZN(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n228), .B(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n222), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n195), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT17), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n192), .A2(new_n194), .A3(new_n222), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n210), .A2(new_n211), .A3(new_n214), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n204), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n215), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n224), .A2(KEYINPUT17), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n237), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(new_n230), .A3(new_n209), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n232), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(G475), .A2(G902), .ZN(new_n246));
  XOR2_X1   g060(.A(new_n246), .B(KEYINPUT91), .Z(new_n247));
  AOI21_X1  g061(.A(KEYINPUT20), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT20), .ZN(new_n249));
  INV_X1    g063(.A(new_n247), .ZN(new_n250));
  AOI211_X1 g064(.A(new_n249), .B(new_n250), .C1(new_n232), .C2(new_n244), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n243), .A2(new_n209), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(new_n230), .ZN(new_n254));
  OAI21_X1  g068(.A(G475), .B1(new_n254), .B2(G902), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT92), .ZN(new_n258));
  INV_X1    g072(.A(G122), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G116), .ZN(new_n260));
  INV_X1    g074(.A(G116), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G122), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n258), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n260), .A2(new_n262), .A3(new_n258), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(G107), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G107), .ZN(new_n267));
  INV_X1    g081(.A(new_n265), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n267), .B1(new_n268), .B2(new_n263), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G128), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(G143), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(G143), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT13), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n278), .B1(new_n271), .B2(G143), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT93), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n272), .A2(KEYINPUT13), .ZN(new_n282));
  OAI211_X1 g096(.A(KEYINPUT93), .B(new_n278), .C1(new_n271), .C2(G143), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n281), .A2(new_n282), .A3(new_n274), .A4(new_n283), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n284), .A2(KEYINPUT94), .A3(G134), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT94), .B1(new_n284), .B2(G134), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n270), .B(new_n277), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT95), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n284), .A2(G134), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT94), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n284), .A2(KEYINPUT94), .A3(G134), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n294), .A2(KEYINPUT95), .A3(new_n277), .A4(new_n270), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n275), .B(new_n276), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n262), .A2(KEYINPUT14), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n260), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n262), .A2(KEYINPUT14), .ZN(new_n299));
  OAI21_X1  g113(.A(G107), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n296), .A2(new_n269), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n289), .A2(new_n295), .A3(new_n301), .ZN(new_n302));
  XOR2_X1   g116(.A(KEYINPUT9), .B(G234), .Z(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G217), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n304), .A2(new_n305), .A3(G953), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n289), .A2(new_n295), .A3(new_n301), .A4(new_n306), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(KEYINPUT96), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G902), .ZN(new_n311));
  INV_X1    g125(.A(new_n302), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT96), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(new_n306), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G478), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(KEYINPUT15), .ZN(new_n317));
  OR2_X1    g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G234), .ZN(new_n319));
  INV_X1    g133(.A(G237), .ZN(new_n320));
  OAI211_X1 g134(.A(G902), .B(G953), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(KEYINPUT97), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT21), .B(G898), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n187), .A2(G952), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n319), .B2(new_n320), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n315), .A2(new_n317), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n257), .A2(new_n318), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(G214), .B1(G237), .B2(G902), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G119), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G116), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n261), .A2(G119), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT2), .B(G113), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(KEYINPUT5), .ZN(new_n339));
  OAI21_X1  g153(.A(G113), .B1(new_n333), .B2(KEYINPUT5), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n338), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n267), .A2(G104), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT79), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n267), .A2(G104), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n344), .B(G101), .C1(new_n347), .C2(new_n343), .ZN(new_n348));
  INV_X1    g162(.A(new_n343), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n350));
  OAI22_X1  g164(.A1(new_n350), .A2(KEYINPUT3), .B1(new_n229), .B2(G107), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n349), .B(new_n351), .C1(new_n352), .C2(new_n345), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n348), .B1(new_n353), .B2(G101), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT8), .ZN(new_n355));
  XOR2_X1   g169(.A(G110), .B(G122), .Z(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n342), .A2(new_n354), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n339), .B(KEYINPUT88), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n338), .B1(new_n359), .B2(new_n341), .ZN(new_n360));
  OAI221_X1 g174(.A(new_n358), .B1(new_n355), .B2(new_n357), .C1(new_n360), .C2(new_n354), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(KEYINPUT89), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n229), .A2(G107), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n350), .A2(KEYINPUT3), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT3), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(KEYINPUT78), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n363), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G101), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n367), .A2(new_n368), .A3(new_n349), .A4(new_n351), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n369), .A2(new_n370), .A3(new_n348), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n370), .B1(new_n369), .B2(new_n348), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n342), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n353), .A2(G101), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT4), .A3(new_n369), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n335), .B(new_n337), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n353), .A2(new_n378), .A3(G101), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n375), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n373), .A2(new_n380), .A3(new_n357), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT85), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n373), .A2(KEYINPUT85), .A3(new_n380), .A4(new_n357), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n204), .A2(G143), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n191), .A2(G146), .ZN(new_n387));
  AND2_X1   g201(.A1(KEYINPUT0), .A2(G128), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G143), .B(G146), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT0), .B(G128), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G125), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n271), .A2(KEYINPUT1), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n386), .A3(new_n387), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n191), .B(G146), .C1(new_n271), .C2(KEYINPUT1), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n271), .A2(new_n204), .A3(G143), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n393), .B1(G125), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G224), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(G953), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(KEYINPUT86), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT7), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n399), .B(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n362), .A2(new_n385), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n357), .B1(new_n373), .B2(new_n380), .ZN(new_n407));
  OR2_X1    g221(.A1(new_n407), .A2(KEYINPUT6), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n407), .B1(new_n383), .B2(new_n384), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n399), .B(new_n402), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n411), .A2(KEYINPUT87), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT87), .B1(new_n411), .B2(new_n412), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n311), .B(new_n406), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(G210), .B1(G237), .B2(G902), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n411), .A2(new_n412), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n411), .A2(KEYINPUT87), .A3(new_n412), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n423), .A2(new_n311), .A3(new_n416), .A4(new_n406), .ZN(new_n424));
  AOI211_X1 g238(.A(new_n329), .B(new_n331), .C1(new_n418), .C2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT74), .ZN(new_n426));
  XOR2_X1   g240(.A(KEYINPUT24), .B(G110), .Z(new_n427));
  INV_X1    g241(.A(KEYINPUT72), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n428), .B1(new_n271), .B2(G119), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n332), .A2(KEYINPUT72), .A3(G128), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n429), .A2(new_n430), .B1(G119), .B2(new_n271), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n239), .A2(new_n215), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT23), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(G119), .B2(new_n271), .ZN(new_n434));
  NOR3_X1   g248(.A1(new_n332), .A2(KEYINPUT23), .A3(G128), .ZN(new_n435));
  OAI22_X1  g249(.A1(new_n434), .A2(new_n435), .B1(G119), .B2(new_n271), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G110), .ZN(new_n437));
  OAI22_X1  g251(.A1(new_n436), .A2(G110), .B1(new_n431), .B2(new_n427), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n215), .A2(new_n205), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n432), .A2(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(KEYINPUT22), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(G137), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n426), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n431), .A2(new_n427), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n240), .A2(new_n437), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n439), .A2(new_n438), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n443), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(KEYINPUT74), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT75), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(new_n448), .B2(new_n449), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n440), .A2(KEYINPUT75), .A3(new_n443), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n455), .A3(new_n311), .ZN(new_n456));
  AND2_X1   g270(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n305), .B1(G234), .B2(new_n311), .ZN(new_n459));
  NOR2_X1   g273(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n451), .A2(new_n455), .A3(new_n311), .A4(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n458), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT77), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n458), .A2(KEYINPUT77), .A3(new_n459), .A4(new_n462), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n451), .A2(new_n455), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n459), .A2(G902), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n465), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(G221), .B1(new_n304), .B2(G902), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(G110), .B(G140), .ZN(new_n473));
  INV_X1    g287(.A(G227), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(G953), .ZN(new_n475));
  XOR2_X1   g289(.A(new_n473), .B(new_n475), .Z(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT66), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n392), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n389), .B(KEYINPUT66), .C1(new_n390), .C2(new_n391), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n375), .A2(new_n379), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT80), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n395), .A2(new_n482), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n396), .A2(new_n397), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n390), .A2(KEYINPUT80), .A3(new_n394), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n369), .A3(new_n348), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT10), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n481), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT11), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n491), .B1(new_n276), .B2(G137), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n276), .A2(G137), .ZN(new_n493));
  INV_X1    g307(.A(G137), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(KEYINPUT11), .A3(G134), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G131), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n222), .A2(new_n493), .A3(new_n492), .A4(new_n495), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g313(.A(KEYINPUT10), .B(new_n398), .C1(new_n371), .C2(new_n372), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n490), .A2(KEYINPUT82), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n500), .A2(new_n499), .A3(new_n489), .A4(new_n481), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT82), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n477), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n490), .A2(new_n500), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n497), .A2(new_n498), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n398), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n354), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n487), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT12), .B1(new_n512), .B2(new_n507), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT12), .ZN(new_n514));
  AOI211_X1 g328(.A(new_n514), .B(new_n499), .C1(new_n511), .C2(new_n487), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n516), .B1(new_n501), .B2(new_n504), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n509), .B(G469), .C1(new_n476), .C2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT83), .ZN(new_n519));
  NAND2_X1  g333(.A1(G469), .A2(G902), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n501), .A2(new_n504), .ZN(new_n522));
  INV_X1    g336(.A(new_n516), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n524), .A2(new_n477), .B1(new_n505), .B2(new_n508), .ZN(new_n525));
  OAI211_X1 g339(.A(KEYINPUT83), .B(G469), .C1(new_n525), .C2(G902), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G469), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n476), .B1(new_n522), .B2(new_n508), .ZN(new_n529));
  AOI211_X1 g343(.A(new_n477), .B(new_n516), .C1(new_n501), .C2(new_n504), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n528), .B(new_n311), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT84), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n502), .A2(new_n503), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n502), .A2(new_n503), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n508), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n477), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n505), .A2(new_n523), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT84), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n538), .A2(new_n539), .A3(new_n528), .A4(new_n311), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n532), .A2(new_n540), .ZN(new_n541));
  AOI211_X1 g355(.A(new_n470), .B(new_n472), .C1(new_n527), .C2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(G472), .A2(G902), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n479), .A2(new_n507), .A3(new_n480), .ZN(new_n544));
  INV_X1    g358(.A(new_n493), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n276), .A2(G137), .ZN(new_n546));
  OAI21_X1  g360(.A(G131), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n398), .A2(new_n498), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n544), .A2(KEYINPUT30), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT65), .ZN(new_n550));
  INV_X1    g364(.A(new_n392), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n507), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n507), .B2(new_n551), .ZN(new_n553));
  INV_X1    g367(.A(new_n548), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n377), .B(new_n549), .C1(new_n555), .C2(KEYINPUT30), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT67), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n193), .A2(G210), .A3(new_n187), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(KEYINPUT27), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT26), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n558), .A2(KEYINPUT27), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT26), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n558), .A2(KEYINPUT27), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n368), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n560), .A2(new_n564), .A3(G101), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n544), .A2(new_n376), .A3(new_n548), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT65), .B1(new_n499), .B2(new_n392), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n507), .A2(new_n550), .A3(new_n551), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n548), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT30), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT67), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n575), .A2(new_n576), .A3(new_n377), .A4(new_n549), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n557), .A2(new_n569), .A3(new_n570), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT31), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n544), .A2(KEYINPUT69), .A3(new_n548), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT69), .B1(new_n544), .B2(new_n548), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n581), .A2(new_n582), .A3(new_n377), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(KEYINPUT28), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT28), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n573), .A2(new_n377), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n585), .B1(new_n586), .B2(new_n570), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n568), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n578), .B2(KEYINPUT31), .ZN(new_n589));
  OAI211_X1 g403(.A(KEYINPUT32), .B(new_n543), .C1(new_n580), .C2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT71), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n557), .A2(new_n570), .A3(new_n577), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT31), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n594), .A3(new_n569), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(new_n579), .A3(new_n588), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n596), .A2(KEYINPUT71), .A3(KEYINPUT32), .A4(new_n543), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n593), .A2(new_n568), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n584), .A2(new_n587), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n569), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT29), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n569), .A2(KEYINPUT29), .ZN(new_n603));
  INV_X1    g417(.A(new_n570), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n376), .B1(new_n544), .B2(new_n548), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT28), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(new_n583), .B2(KEYINPUT28), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n311), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(G472), .B1(new_n602), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n543), .B1(new_n580), .B2(new_n589), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT70), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT32), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n611), .B1(new_n610), .B2(new_n612), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n598), .B(new_n609), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n425), .A2(new_n542), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT98), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n418), .A2(new_n424), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n310), .A2(new_n622), .A3(new_n314), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n308), .A2(KEYINPUT33), .A3(new_n309), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n316), .A2(G902), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n315), .A2(new_n316), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n256), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n415), .A2(KEYINPUT99), .A3(new_n417), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n621), .A2(new_n330), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n327), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n527), .A2(new_n541), .ZN(new_n635));
  INV_X1    g449(.A(new_n470), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n311), .B1(new_n580), .B2(new_n589), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(G472), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n638), .A2(new_n610), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n635), .A2(new_n636), .A3(new_n639), .A4(new_n471), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  AND3_X1   g458(.A1(new_n621), .A2(new_n330), .A3(new_n631), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n327), .B(KEYINPUT100), .Z(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n256), .B1(new_n318), .B2(new_n328), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n645), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n640), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT35), .B(G107), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  AOI21_X1  g466(.A(G902), .B1(new_n536), .B2(new_n537), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n539), .B1(new_n653), .B2(new_n528), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n531), .A2(KEYINPUT84), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n521), .A2(new_n526), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n471), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n449), .A2(KEYINPUT36), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(new_n448), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n468), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n465), .A2(new_n466), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n465), .A2(KEYINPUT101), .A3(new_n466), .A4(new_n661), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n658), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n425), .A3(new_n639), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT37), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n669), .B(G110), .Z(G12));
  INV_X1    g484(.A(new_n326), .ZN(new_n671));
  INV_X1    g485(.A(G900), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n671), .B1(new_n322), .B2(new_n672), .ZN(new_n673));
  AOI211_X1 g487(.A(new_n673), .B(new_n256), .C1(new_n318), .C2(new_n328), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n645), .A2(new_n667), .A3(new_n616), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  XOR2_X1   g490(.A(new_n673), .B(KEYINPUT39), .Z(new_n677));
  NAND3_X1  g491(.A1(new_n635), .A2(new_n471), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n678), .B(KEYINPUT40), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n418), .A2(new_n424), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n257), .B1(new_n328), .B2(new_n318), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n666), .A2(new_n330), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT103), .ZN(new_n685));
  INV_X1    g499(.A(new_n593), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n569), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n604), .A2(new_n605), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n311), .B1(new_n569), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n598), .B(new_n691), .C1(new_n614), .C2(new_n615), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n679), .A2(new_n682), .A3(new_n685), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G143), .ZN(G45));
  AOI221_X4 g508(.A(new_n673), .B1(new_n255), .B2(new_n252), .C1(new_n626), .C2(new_n627), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n645), .A2(new_n667), .A3(new_n616), .A4(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT104), .B(G146), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G48));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n645), .A2(new_n327), .A3(new_n630), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n653), .A2(new_n528), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n541), .A2(new_n471), .A3(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n616), .A2(new_n636), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n699), .B1(new_n700), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n610), .A2(new_n612), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT70), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n707), .A2(new_n613), .B1(new_n597), .B2(new_n592), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n470), .B1(new_n708), .B2(new_n609), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n634), .A2(KEYINPUT105), .A3(new_n709), .A4(new_n703), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n705), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT41), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G113), .ZN(G15));
  NOR2_X1   g527(.A1(new_n649), .A2(new_n704), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n261), .ZN(G18));
  INV_X1    g529(.A(new_n666), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n702), .A2(new_n329), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n645), .A2(new_n616), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n470), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n607), .A2(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n606), .B(KEYINPUT106), .C1(new_n583), .C2(KEYINPUT28), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n723), .A2(new_n568), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n595), .A2(new_n579), .A3(new_n725), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n637), .A2(G472), .B1(new_n726), .B2(new_n543), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n465), .A2(KEYINPUT107), .A3(new_n466), .A4(new_n469), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n721), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n729), .A2(new_n702), .A3(new_n646), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n645), .A2(new_n683), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  AND4_X1   g546(.A1(new_n664), .A2(new_n727), .A3(new_n665), .A4(new_n695), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n645), .A2(new_n703), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G125), .ZN(G27));
  NAND2_X1  g549(.A1(new_n518), .A2(new_n520), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n737), .B1(new_n654), .B2(new_n655), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(KEYINPUT108), .A3(new_n471), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n736), .B1(new_n532), .B2(new_n540), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n740), .B1(new_n741), .B2(new_n472), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n418), .A2(new_n424), .A3(new_n330), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n743), .A2(new_n709), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n695), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(KEYINPUT42), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n721), .A2(new_n728), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n609), .A2(new_n706), .A3(new_n590), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n743), .A2(new_n751), .A3(new_n695), .A4(new_n744), .ZN(new_n752));
  AOI22_X1  g566(.A1(new_n745), .A2(new_n747), .B1(new_n752), .B2(KEYINPUT42), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  NAND4_X1  g568(.A1(new_n743), .A2(new_n709), .A3(new_n674), .A4(new_n744), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  NAND2_X1  g570(.A1(new_n628), .A2(new_n257), .ZN(new_n757));
  XOR2_X1   g571(.A(new_n757), .B(KEYINPUT43), .Z(new_n758));
  NAND2_X1  g572(.A1(new_n638), .A2(new_n610), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n759), .A3(new_n716), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT44), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n744), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n509), .B1(new_n476), .B2(new_n517), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n528), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n525), .A2(KEYINPUT45), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n767), .A2(new_n768), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n520), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n520), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n541), .A3(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n777), .A2(new_n471), .A3(new_n677), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n761), .A2(KEYINPUT110), .A3(new_n744), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n764), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G137), .ZN(G39));
  NAND2_X1  g595(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n777), .B2(new_n471), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n520), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT46), .B1(new_n772), .B2(new_n520), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n784), .A2(new_n785), .A3(new_n656), .ZN(new_n786));
  OAI22_X1  g600(.A1(new_n786), .A2(new_n472), .B1(KEYINPUT111), .B2(KEYINPUT47), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n783), .B1(new_n787), .B2(new_n782), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n744), .A2(new_n695), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n789), .A2(new_n616), .A3(new_n636), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT112), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  NAND2_X1  g607(.A1(new_n758), .A2(new_n671), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n729), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n541), .A2(new_n701), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n471), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n744), .B(new_n795), .C1(new_n788), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n744), .A2(new_n703), .ZN(new_n799));
  OR4_X1    g613(.A1(new_n326), .A2(new_n799), .A3(new_n470), .A4(new_n692), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n800), .A2(new_n256), .A3(new_n628), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n716), .A2(new_n727), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n794), .A2(new_n799), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n794), .A2(new_n702), .A3(new_n729), .ZN(new_n805));
  INV_X1    g619(.A(new_n682), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n331), .A3(new_n806), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT50), .Z(new_n808));
  NAND3_X1  g622(.A1(new_n798), .A2(new_n804), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n811), .B1(new_n809), .B2(new_n810), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n803), .A2(new_n751), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT48), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n815), .B(new_n325), .C1(new_n629), .C2(new_n800), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n812), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n621), .A2(new_n330), .A3(new_n631), .A4(new_n683), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n738), .A2(new_n471), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n662), .A2(new_n673), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n692), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n818), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n823), .A2(new_n819), .A3(KEYINPUT119), .A4(new_n820), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n675), .A2(new_n696), .A3(new_n734), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n827), .A2(KEYINPUT52), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n825), .ZN(new_n830));
  INV_X1    g644(.A(new_n826), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n675), .A2(new_n734), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(KEYINPUT118), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n675), .B2(new_n734), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n832), .B(new_n696), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n829), .B1(new_n837), .B2(KEYINPUT52), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n743), .A2(new_n839), .A3(new_n733), .A4(new_n744), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n257), .A2(new_n318), .A3(new_n328), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n673), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n667), .A2(new_n616), .A3(new_n744), .A4(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n733), .A2(new_n744), .A3(new_n739), .A4(new_n742), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT115), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n755), .A2(new_n840), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT116), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n714), .B1(new_n705), .B2(new_n710), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n680), .A2(new_n330), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n640), .A2(new_n849), .A3(new_n629), .A4(new_n646), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n425), .A2(new_n542), .A3(new_n616), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT114), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n853));
  INV_X1    g667(.A(new_n849), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(new_n542), .A3(new_n639), .A4(new_n647), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n617), .B(new_n853), .C1(new_n855), .C2(new_n629), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n641), .A2(new_n854), .A3(new_n647), .A4(new_n648), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n858), .A2(new_n718), .A3(new_n731), .A4(new_n668), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n848), .A2(new_n857), .A3(new_n860), .A4(new_n753), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n847), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n838), .A2(new_n862), .A3(KEYINPUT53), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n844), .B(new_n839), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n865), .A2(KEYINPUT116), .A3(new_n755), .A4(new_n843), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n846), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n859), .B1(new_n852), .B2(new_n856), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n869), .A2(new_n753), .A3(new_n870), .A4(new_n848), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT52), .ZN(new_n872));
  INV_X1    g686(.A(new_n828), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n832), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT52), .B1(new_n827), .B2(new_n828), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n864), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n863), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n871), .A2(new_n876), .A3(new_n864), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n862), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n871), .A2(KEYINPUT117), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n882), .A2(new_n838), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n880), .B1(new_n884), .B2(new_n864), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n817), .B(new_n879), .C1(new_n878), .C2(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n805), .A2(new_n645), .ZN(new_n887));
  OAI22_X1  g701(.A1(new_n886), .A2(new_n887), .B1(G952), .B2(G953), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n796), .A2(KEYINPUT49), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n757), .A2(new_n472), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n748), .A3(new_n330), .A4(new_n890), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT113), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n806), .B1(KEYINPUT49), .B2(new_n796), .ZN(new_n893));
  OR3_X1    g707(.A1(new_n892), .A2(new_n893), .A3(new_n692), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n888), .A2(new_n894), .ZN(G75));
  XNOR2_X1  g709(.A(new_n411), .B(new_n412), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT55), .ZN(new_n897));
  INV_X1    g711(.A(G210), .ZN(new_n898));
  AOI211_X1 g712(.A(new_n898), .B(new_n311), .C1(new_n863), .C2(new_n877), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n897), .B1(new_n899), .B2(KEYINPUT56), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n187), .A2(G952), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n863), .A2(new_n877), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(G210), .A3(G902), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  INV_X1    g719(.A(new_n897), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n900), .A2(new_n902), .A3(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n900), .A2(KEYINPUT121), .A3(new_n907), .A4(new_n902), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(G51));
  XOR2_X1   g726(.A(new_n520), .B(KEYINPUT57), .Z(new_n913));
  AND3_X1   g727(.A1(new_n863), .A2(new_n877), .A3(new_n878), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n878), .B1(new_n863), .B2(new_n877), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g732(.A(KEYINPUT122), .B(new_n913), .C1(new_n914), .C2(new_n915), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n538), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n903), .A2(G902), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n921), .A2(new_n772), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n901), .B1(new_n920), .B2(new_n922), .ZN(G54));
  NAND4_X1  g737(.A1(new_n903), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n924));
  INV_X1    g738(.A(new_n245), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n901), .ZN(G60));
  OAI21_X1  g742(.A(new_n879), .B1(new_n885), .B2(new_n878), .ZN(new_n929));
  NAND2_X1  g743(.A1(G478), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT59), .Z(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AOI22_X1  g746(.A1(new_n929), .A2(new_n932), .B1(new_n623), .B2(new_n624), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n914), .A2(new_n915), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n623), .A2(new_n624), .A3(new_n932), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n933), .A2(new_n901), .A3(new_n936), .ZN(G63));
  NAND2_X1  g751(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n938));
  OR2_X1    g752(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n939));
  NAND2_X1  g753(.A1(G217), .A2(G902), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT60), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n863), .B2(new_n877), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n942), .A2(new_n660), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n902), .B1(new_n942), .B2(new_n467), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n938), .B(new_n939), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NOR4_X1   g760(.A1(new_n943), .A2(new_n944), .A3(KEYINPUT123), .A4(KEYINPUT61), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(G66));
  NAND2_X1  g762(.A1(new_n870), .A2(new_n848), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n187), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT124), .ZN(new_n951));
  OAI21_X1  g765(.A(G953), .B1(new_n323), .B2(new_n400), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT125), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n411), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(G898), .B2(new_n187), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n954), .B(new_n956), .ZN(G69));
  XNOR2_X1  g771(.A(new_n833), .B(KEYINPUT118), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n958), .A2(new_n693), .A3(new_n696), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n648), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n678), .B1(new_n962), .B2(new_n629), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n963), .A2(new_n709), .A3(new_n744), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n780), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n961), .A2(new_n792), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(KEYINPUT127), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n961), .A2(new_n968), .A3(new_n792), .A4(new_n965), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n575), .A2(new_n549), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT126), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n216), .A2(new_n218), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n970), .A2(new_n187), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n672), .B1(new_n974), .B2(new_n474), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n958), .A2(new_n696), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n792), .A2(new_n753), .A3(new_n755), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n764), .A2(new_n779), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(new_n819), .B2(new_n750), .ZN(new_n980));
  AOI211_X1 g794(.A(new_n977), .B(new_n978), .C1(new_n778), .C2(new_n980), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n981), .A2(G953), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n982), .A2(new_n974), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n187), .A2(G227), .ZN(new_n984));
  OAI221_X1 g798(.A(new_n975), .B1(new_n187), .B2(new_n976), .C1(new_n983), .C2(new_n984), .ZN(G72));
  NAND3_X1  g799(.A1(new_n967), .A2(new_n688), .A3(new_n969), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n981), .A2(new_n568), .A3(new_n593), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n949), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n687), .A2(new_n599), .ZN(new_n989));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT63), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n902), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n885), .A2(new_n991), .A3(new_n989), .ZN(new_n994));
  NOR3_X1   g808(.A1(new_n988), .A2(new_n993), .A3(new_n994), .ZN(G57));
endmodule


