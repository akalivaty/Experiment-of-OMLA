

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U547 ( .A(n751), .B(KEYINPUT93), .Z(n511) );
  INV_X1 U548 ( .A(KEYINPUT31), .ZN(n720) );
  XNOR2_X1 U549 ( .A(n720), .B(KEYINPUT94), .ZN(n721) );
  XNOR2_X1 U550 ( .A(n722), .B(n721), .ZN(n752) );
  NAND2_X1 U551 ( .A1(n710), .A2(n709), .ZN(n725) );
  NOR2_X2 U552 ( .A1(G2105), .A2(n522), .ZN(n861) );
  NOR2_X1 U553 ( .A1(G651), .A2(n631), .ZN(n625) );
  NOR2_X1 U554 ( .A1(G651), .A2(G543), .ZN(n617) );
  NAND2_X1 U555 ( .A1(G91), .A2(n617), .ZN(n514) );
  INV_X1 U556 ( .A(G651), .ZN(n516) );
  XOR2_X1 U557 ( .A(KEYINPUT0), .B(G543), .Z(n631) );
  OR2_X1 U558 ( .A1(n516), .A2(n631), .ZN(n512) );
  XNOR2_X1 U559 ( .A(KEYINPUT67), .B(n512), .ZN(n622) );
  NAND2_X1 U560 ( .A1(G78), .A2(n622), .ZN(n513) );
  NAND2_X1 U561 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U562 ( .A(KEYINPUT69), .B(n515), .ZN(n521) );
  NOR2_X1 U563 ( .A1(G543), .A2(n516), .ZN(n517) );
  XOR2_X1 U564 ( .A(KEYINPUT1), .B(n517), .Z(n630) );
  NAND2_X1 U565 ( .A1(G65), .A2(n630), .ZN(n519) );
  NAND2_X1 U566 ( .A1(G53), .A2(n625), .ZN(n518) );
  AND2_X1 U567 ( .A1(n519), .A2(n518), .ZN(n520) );
  NAND2_X1 U568 ( .A1(n521), .A2(n520), .ZN(G299) );
  INV_X1 U569 ( .A(G2104), .ZN(n522) );
  NAND2_X1 U570 ( .A1(G101), .A2(n861), .ZN(n524) );
  XOR2_X1 U571 ( .A(KEYINPUT64), .B(KEYINPUT23), .Z(n523) );
  XNOR2_X1 U572 ( .A(n524), .B(n523), .ZN(n526) );
  AND2_X1 U573 ( .A1(n522), .A2(G2105), .ZN(n857) );
  NAND2_X1 U574 ( .A1(n857), .A2(G125), .ZN(n525) );
  NAND2_X1 U575 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U576 ( .A(n527), .B(KEYINPUT65), .ZN(n677) );
  NOR2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  XOR2_X2 U578 ( .A(KEYINPUT17), .B(n528), .Z(n862) );
  NAND2_X1 U579 ( .A1(G137), .A2(n862), .ZN(n675) );
  AND2_X1 U580 ( .A1(n677), .A2(n675), .ZN(n530) );
  AND2_X1 U581 ( .A1(G2104), .A2(G2105), .ZN(n858) );
  NAND2_X1 U582 ( .A1(G113), .A2(n858), .ZN(n529) );
  XNOR2_X1 U583 ( .A(KEYINPUT66), .B(n529), .ZN(n673) );
  AND2_X1 U584 ( .A1(n530), .A2(n673), .ZN(G160) );
  NAND2_X1 U585 ( .A1(G90), .A2(n617), .ZN(n532) );
  NAND2_X1 U586 ( .A1(G77), .A2(n622), .ZN(n531) );
  NAND2_X1 U587 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U588 ( .A(n533), .B(KEYINPUT9), .ZN(n535) );
  NAND2_X1 U589 ( .A1(G64), .A2(n630), .ZN(n534) );
  NAND2_X1 U590 ( .A1(n535), .A2(n534), .ZN(n538) );
  NAND2_X1 U591 ( .A1(n625), .A2(G52), .ZN(n536) );
  XOR2_X1 U592 ( .A(KEYINPUT68), .B(n536), .Z(n537) );
  NOR2_X1 U593 ( .A1(n538), .A2(n537), .ZN(G171) );
  AND2_X1 U594 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U595 ( .A1(G99), .A2(n861), .ZN(n540) );
  NAND2_X1 U596 ( .A1(G111), .A2(n858), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U598 ( .A(KEYINPUT78), .B(n541), .ZN(n547) );
  NAND2_X1 U599 ( .A1(G123), .A2(n857), .ZN(n542) );
  XOR2_X1 U600 ( .A(KEYINPUT77), .B(n542), .Z(n543) );
  XNOR2_X1 U601 ( .A(n543), .B(KEYINPUT18), .ZN(n545) );
  NAND2_X1 U602 ( .A1(G135), .A2(n862), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U604 ( .A1(n547), .A2(n546), .ZN(n968) );
  XNOR2_X1 U605 ( .A(n968), .B(G2096), .ZN(n548) );
  XNOR2_X1 U606 ( .A(n548), .B(KEYINPUT79), .ZN(n549) );
  OR2_X1 U607 ( .A1(G2100), .A2(n549), .ZN(G156) );
  INV_X1 U608 ( .A(G57), .ZN(G237) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  NAND2_X1 U611 ( .A1(n625), .A2(G51), .ZN(n550) );
  XOR2_X1 U612 ( .A(KEYINPUT75), .B(n550), .Z(n552) );
  NAND2_X1 U613 ( .A1(n630), .A2(G63), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U615 ( .A(KEYINPUT6), .B(n553), .ZN(n560) );
  NAND2_X1 U616 ( .A1(G89), .A2(n617), .ZN(n554) );
  XNOR2_X1 U617 ( .A(n554), .B(KEYINPUT74), .ZN(n555) );
  XNOR2_X1 U618 ( .A(n555), .B(KEYINPUT4), .ZN(n557) );
  NAND2_X1 U619 ( .A1(G76), .A2(n622), .ZN(n556) );
  NAND2_X1 U620 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U621 ( .A(n558), .B(KEYINPUT5), .Z(n559) );
  NOR2_X1 U622 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U623 ( .A(KEYINPUT7), .B(n561), .Z(n562) );
  XNOR2_X1 U624 ( .A(KEYINPUT76), .B(n562), .ZN(G168) );
  XOR2_X1 U625 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U626 ( .A1(G7), .A2(G661), .ZN(n563) );
  XNOR2_X1 U627 ( .A(n563), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U628 ( .A(G223), .ZN(n812) );
  NAND2_X1 U629 ( .A1(n812), .A2(G567), .ZN(n564) );
  XOR2_X1 U630 ( .A(KEYINPUT11), .B(n564), .Z(G234) );
  NAND2_X1 U631 ( .A1(G56), .A2(n630), .ZN(n565) );
  XOR2_X1 U632 ( .A(KEYINPUT14), .B(n565), .Z(n571) );
  NAND2_X1 U633 ( .A1(n617), .A2(G81), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n566), .B(KEYINPUT12), .ZN(n568) );
  NAND2_X1 U635 ( .A1(G68), .A2(n622), .ZN(n567) );
  NAND2_X1 U636 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U637 ( .A(KEYINPUT13), .B(n569), .Z(n570) );
  NOR2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n625), .A2(G43), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n940) );
  XOR2_X1 U641 ( .A(G860), .B(KEYINPUT70), .Z(n587) );
  NOR2_X1 U642 ( .A1(n940), .A2(n587), .ZN(n574) );
  XNOR2_X1 U643 ( .A(n574), .B(KEYINPUT71), .ZN(G153) );
  XOR2_X1 U644 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U645 ( .A1(G868), .A2(G301), .ZN(n584) );
  NAND2_X1 U646 ( .A1(n622), .A2(G79), .ZN(n581) );
  NAND2_X1 U647 ( .A1(G66), .A2(n630), .ZN(n576) );
  NAND2_X1 U648 ( .A1(G92), .A2(n617), .ZN(n575) );
  NAND2_X1 U649 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U650 ( .A1(G54), .A2(n625), .ZN(n577) );
  XNOR2_X1 U651 ( .A(KEYINPUT73), .B(n577), .ZN(n578) );
  NOR2_X1 U652 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U653 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U654 ( .A(KEYINPUT15), .B(n582), .Z(n947) );
  INV_X1 U655 ( .A(G868), .ZN(n634) );
  NAND2_X1 U656 ( .A1(n947), .A2(n634), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n584), .A2(n583), .ZN(G284) );
  NAND2_X1 U658 ( .A1(G868), .A2(G286), .ZN(n586) );
  NAND2_X1 U659 ( .A1(G299), .A2(n634), .ZN(n585) );
  NAND2_X1 U660 ( .A1(n586), .A2(n585), .ZN(G297) );
  NAND2_X1 U661 ( .A1(n587), .A2(G559), .ZN(n588) );
  INV_X1 U662 ( .A(n947), .ZN(n884) );
  NAND2_X1 U663 ( .A1(n588), .A2(n884), .ZN(n589) );
  XNOR2_X1 U664 ( .A(n589), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U665 ( .A1(G868), .A2(n940), .ZN(n592) );
  NAND2_X1 U666 ( .A1(G868), .A2(n884), .ZN(n590) );
  NOR2_X1 U667 ( .A1(G559), .A2(n590), .ZN(n591) );
  NOR2_X1 U668 ( .A1(n592), .A2(n591), .ZN(G282) );
  NAND2_X1 U669 ( .A1(G93), .A2(n617), .ZN(n594) );
  NAND2_X1 U670 ( .A1(G55), .A2(n625), .ZN(n593) );
  NAND2_X1 U671 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U672 ( .A1(n622), .A2(G80), .ZN(n595) );
  XOR2_X1 U673 ( .A(KEYINPUT80), .B(n595), .Z(n596) );
  NOR2_X1 U674 ( .A1(n597), .A2(n596), .ZN(n599) );
  NAND2_X1 U675 ( .A1(n630), .A2(G67), .ZN(n598) );
  NAND2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n635) );
  NAND2_X1 U677 ( .A1(n884), .A2(G559), .ZN(n642) );
  XNOR2_X1 U678 ( .A(n940), .B(n642), .ZN(n600) );
  NOR2_X1 U679 ( .A1(G860), .A2(n600), .ZN(n601) );
  XOR2_X1 U680 ( .A(KEYINPUT81), .B(n601), .Z(n602) );
  XOR2_X1 U681 ( .A(n635), .B(n602), .Z(G145) );
  NAND2_X1 U682 ( .A1(G61), .A2(n630), .ZN(n604) );
  NAND2_X1 U683 ( .A1(G86), .A2(n617), .ZN(n603) );
  NAND2_X1 U684 ( .A1(n604), .A2(n603), .ZN(n607) );
  NAND2_X1 U685 ( .A1(n622), .A2(G73), .ZN(n605) );
  XOR2_X1 U686 ( .A(KEYINPUT2), .B(n605), .Z(n606) );
  NOR2_X1 U687 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U688 ( .A(KEYINPUT83), .B(n608), .Z(n610) );
  NAND2_X1 U689 ( .A1(n625), .A2(G48), .ZN(n609) );
  NAND2_X1 U690 ( .A1(n610), .A2(n609), .ZN(G305) );
  NAND2_X1 U691 ( .A1(G88), .A2(n617), .ZN(n612) );
  NAND2_X1 U692 ( .A1(G75), .A2(n622), .ZN(n611) );
  NAND2_X1 U693 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U694 ( .A1(G62), .A2(n630), .ZN(n614) );
  NAND2_X1 U695 ( .A1(G50), .A2(n625), .ZN(n613) );
  NAND2_X1 U696 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U697 ( .A1(n616), .A2(n615), .ZN(G166) );
  AND2_X1 U698 ( .A1(n617), .A2(G85), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G60), .A2(n630), .ZN(n619) );
  NAND2_X1 U700 ( .A1(G47), .A2(n625), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n622), .A2(G72), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n624), .A2(n623), .ZN(G290) );
  NAND2_X1 U705 ( .A1(G49), .A2(n625), .ZN(n627) );
  NAND2_X1 U706 ( .A1(G74), .A2(G651), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U708 ( .A(KEYINPUT82), .B(n628), .ZN(n629) );
  NOR2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n631), .A2(G87), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(G288) );
  NAND2_X1 U712 ( .A1(n635), .A2(n634), .ZN(n645) );
  INV_X1 U713 ( .A(G299), .ZN(n938) );
  XNOR2_X1 U714 ( .A(n938), .B(n940), .ZN(n638) );
  XOR2_X1 U715 ( .A(KEYINPUT19), .B(n635), .Z(n636) );
  XNOR2_X1 U716 ( .A(n636), .B(G290), .ZN(n637) );
  XNOR2_X1 U717 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U718 ( .A(G166), .B(n639), .ZN(n640) );
  XNOR2_X1 U719 ( .A(n640), .B(G288), .ZN(n641) );
  XNOR2_X1 U720 ( .A(G305), .B(n641), .ZN(n883) );
  XNOR2_X1 U721 ( .A(n883), .B(n642), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n643), .A2(G868), .ZN(n644) );
  NAND2_X1 U723 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U724 ( .A(n646), .B(KEYINPUT84), .ZN(G295) );
  NAND2_X1 U725 ( .A1(G2084), .A2(G2078), .ZN(n647) );
  XOR2_X1 U726 ( .A(KEYINPUT20), .B(n647), .Z(n648) );
  NAND2_X1 U727 ( .A1(G2090), .A2(n648), .ZN(n649) );
  XNOR2_X1 U728 ( .A(KEYINPUT21), .B(n649), .ZN(n650) );
  NAND2_X1 U729 ( .A1(n650), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U730 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U731 ( .A1(G220), .A2(G219), .ZN(n651) );
  XOR2_X1 U732 ( .A(KEYINPUT22), .B(n651), .Z(n652) );
  NOR2_X1 U733 ( .A1(G218), .A2(n652), .ZN(n653) );
  NAND2_X1 U734 ( .A1(G96), .A2(n653), .ZN(n904) );
  NAND2_X1 U735 ( .A1(n904), .A2(G2106), .ZN(n657) );
  NAND2_X1 U736 ( .A1(G69), .A2(G120), .ZN(n654) );
  NOR2_X1 U737 ( .A1(G237), .A2(n654), .ZN(n655) );
  NAND2_X1 U738 ( .A1(G108), .A2(n655), .ZN(n903) );
  NAND2_X1 U739 ( .A1(n903), .A2(G567), .ZN(n656) );
  NAND2_X1 U740 ( .A1(n657), .A2(n656), .ZN(n818) );
  NAND2_X1 U741 ( .A1(G483), .A2(G661), .ZN(n658) );
  NOR2_X1 U742 ( .A1(n818), .A2(n658), .ZN(n817) );
  NAND2_X1 U743 ( .A1(n817), .A2(G36), .ZN(G176) );
  NAND2_X1 U744 ( .A1(n861), .A2(G102), .ZN(n661) );
  NAND2_X1 U745 ( .A1(G126), .A2(n857), .ZN(n659) );
  XOR2_X1 U746 ( .A(KEYINPUT85), .B(n659), .Z(n660) );
  NAND2_X1 U747 ( .A1(n661), .A2(n660), .ZN(n665) );
  NAND2_X1 U748 ( .A1(G114), .A2(n858), .ZN(n663) );
  NAND2_X1 U749 ( .A1(G138), .A2(n862), .ZN(n662) );
  NAND2_X1 U750 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U751 ( .A1(n665), .A2(n664), .ZN(G164) );
  INV_X1 U752 ( .A(G166), .ZN(G303) );
  NAND2_X1 U753 ( .A1(G129), .A2(n857), .ZN(n667) );
  NAND2_X1 U754 ( .A1(G117), .A2(n858), .ZN(n666) );
  NAND2_X1 U755 ( .A1(n667), .A2(n666), .ZN(n670) );
  NAND2_X1 U756 ( .A1(n861), .A2(G105), .ZN(n668) );
  XOR2_X1 U757 ( .A(KEYINPUT38), .B(n668), .Z(n669) );
  NOR2_X1 U758 ( .A1(n670), .A2(n669), .ZN(n672) );
  NAND2_X1 U759 ( .A1(n862), .A2(G141), .ZN(n671) );
  NAND2_X1 U760 ( .A1(n672), .A2(n671), .ZN(n871) );
  NOR2_X1 U761 ( .A1(G1996), .A2(n871), .ZN(n960) );
  NOR2_X1 U762 ( .A1(G164), .A2(G1384), .ZN(n709) );
  AND2_X1 U763 ( .A1(G40), .A2(n673), .ZN(n674) );
  AND2_X1 U764 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U765 ( .A1(n677), .A2(n676), .ZN(n708) );
  NOR2_X1 U766 ( .A1(n709), .A2(n708), .ZN(n799) );
  NAND2_X1 U767 ( .A1(G1996), .A2(n871), .ZN(n685) );
  NAND2_X1 U768 ( .A1(G95), .A2(n861), .ZN(n679) );
  NAND2_X1 U769 ( .A1(G107), .A2(n858), .ZN(n678) );
  NAND2_X1 U770 ( .A1(n679), .A2(n678), .ZN(n683) );
  NAND2_X1 U771 ( .A1(G119), .A2(n857), .ZN(n681) );
  NAND2_X1 U772 ( .A1(G131), .A2(n862), .ZN(n680) );
  NAND2_X1 U773 ( .A1(n681), .A2(n680), .ZN(n682) );
  OR2_X1 U774 ( .A1(n683), .A2(n682), .ZN(n876) );
  NAND2_X1 U775 ( .A1(G1991), .A2(n876), .ZN(n684) );
  NAND2_X1 U776 ( .A1(n685), .A2(n684), .ZN(n971) );
  NAND2_X1 U777 ( .A1(n799), .A2(n971), .ZN(n802) );
  INV_X1 U778 ( .A(n802), .ZN(n688) );
  NOR2_X1 U779 ( .A1(G1991), .A2(n876), .ZN(n969) );
  NOR2_X1 U780 ( .A1(G1986), .A2(G290), .ZN(n686) );
  NOR2_X1 U781 ( .A1(n969), .A2(n686), .ZN(n687) );
  NOR2_X1 U782 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U783 ( .A1(n960), .A2(n689), .ZN(n690) );
  XNOR2_X1 U784 ( .A(KEYINPUT39), .B(n690), .ZN(n691) );
  XNOR2_X1 U785 ( .A(n691), .B(KEYINPUT100), .ZN(n701) );
  NAND2_X1 U786 ( .A1(G104), .A2(n861), .ZN(n693) );
  NAND2_X1 U787 ( .A1(G140), .A2(n862), .ZN(n692) );
  NAND2_X1 U788 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U789 ( .A(KEYINPUT34), .B(n694), .ZN(n699) );
  NAND2_X1 U790 ( .A1(G128), .A2(n857), .ZN(n696) );
  NAND2_X1 U791 ( .A1(G116), .A2(n858), .ZN(n695) );
  NAND2_X1 U792 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U793 ( .A(KEYINPUT35), .B(n697), .Z(n698) );
  NOR2_X1 U794 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U795 ( .A(KEYINPUT36), .B(n700), .Z(n880) );
  XOR2_X1 U796 ( .A(KEYINPUT37), .B(G2067), .Z(n703) );
  AND2_X1 U797 ( .A1(n880), .A2(n703), .ZN(n975) );
  NAND2_X1 U798 ( .A1(n799), .A2(n975), .ZN(n804) );
  NAND2_X1 U799 ( .A1(n701), .A2(n804), .ZN(n702) );
  XOR2_X1 U800 ( .A(KEYINPUT101), .B(n702), .Z(n705) );
  NOR2_X1 U801 ( .A1(n880), .A2(n703), .ZN(n704) );
  XOR2_X1 U802 ( .A(KEYINPUT102), .B(n704), .Z(n978) );
  NAND2_X1 U803 ( .A1(n705), .A2(n978), .ZN(n706) );
  NAND2_X1 U804 ( .A1(n706), .A2(n799), .ZN(n809) );
  INV_X1 U805 ( .A(KEYINPUT88), .ZN(n707) );
  XNOR2_X1 U806 ( .A(n708), .B(n707), .ZN(n710) );
  BUF_X2 U807 ( .A(n725), .Z(n754) );
  NAND2_X1 U808 ( .A1(G8), .A2(n754), .ZN(n781) );
  NOR2_X1 U809 ( .A1(G2084), .A2(n754), .ZN(n766) );
  NOR2_X1 U810 ( .A1(n781), .A2(G1966), .ZN(n711) );
  XNOR2_X1 U811 ( .A(n711), .B(KEYINPUT89), .ZN(n768) );
  NAND2_X1 U812 ( .A1(G8), .A2(n768), .ZN(n712) );
  NOR2_X1 U813 ( .A1(n766), .A2(n712), .ZN(n713) );
  XOR2_X1 U814 ( .A(KEYINPUT30), .B(n713), .Z(n714) );
  NOR2_X1 U815 ( .A1(G168), .A2(n714), .ZN(n719) );
  XOR2_X1 U816 ( .A(G2078), .B(KEYINPUT25), .Z(n910) );
  NOR2_X1 U817 ( .A1(n910), .A2(n754), .ZN(n715) );
  XOR2_X1 U818 ( .A(KEYINPUT90), .B(n715), .Z(n717) );
  INV_X1 U819 ( .A(G1961), .ZN(n1003) );
  NAND2_X1 U820 ( .A1(n754), .A2(n1003), .ZN(n716) );
  NAND2_X1 U821 ( .A1(n717), .A2(n716), .ZN(n748) );
  NOR2_X1 U822 ( .A1(G171), .A2(n748), .ZN(n718) );
  NOR2_X1 U823 ( .A1(n719), .A2(n718), .ZN(n722) );
  XOR2_X1 U824 ( .A(KEYINPUT27), .B(KEYINPUT91), .Z(n724) );
  INV_X1 U825 ( .A(n725), .ZN(n734) );
  NAND2_X1 U826 ( .A1(G2072), .A2(n734), .ZN(n723) );
  XNOR2_X1 U827 ( .A(n724), .B(n723), .ZN(n728) );
  NAND2_X1 U828 ( .A1(G1956), .A2(n725), .ZN(n726) );
  XOR2_X1 U829 ( .A(KEYINPUT92), .B(n726), .Z(n727) );
  NOR2_X1 U830 ( .A1(n728), .A2(n727), .ZN(n742) );
  NOR2_X1 U831 ( .A1(n938), .A2(n742), .ZN(n729) );
  XOR2_X1 U832 ( .A(n729), .B(KEYINPUT28), .Z(n746) );
  AND2_X1 U833 ( .A1(n734), .A2(G1996), .ZN(n730) );
  XOR2_X1 U834 ( .A(n730), .B(KEYINPUT26), .Z(n732) );
  NAND2_X1 U835 ( .A1(n754), .A2(G1341), .ZN(n731) );
  NAND2_X1 U836 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U837 ( .A1(n940), .A2(n733), .ZN(n738) );
  NAND2_X1 U838 ( .A1(G1348), .A2(n754), .ZN(n736) );
  NAND2_X1 U839 ( .A1(G2067), .A2(n734), .ZN(n735) );
  NAND2_X1 U840 ( .A1(n736), .A2(n735), .ZN(n739) );
  NOR2_X1 U841 ( .A1(n947), .A2(n739), .ZN(n737) );
  OR2_X1 U842 ( .A1(n738), .A2(n737), .ZN(n741) );
  NAND2_X1 U843 ( .A1(n947), .A2(n739), .ZN(n740) );
  NAND2_X1 U844 ( .A1(n741), .A2(n740), .ZN(n744) );
  NAND2_X1 U845 ( .A1(n938), .A2(n742), .ZN(n743) );
  NAND2_X1 U846 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U847 ( .A1(n746), .A2(n745), .ZN(n747) );
  XOR2_X1 U848 ( .A(KEYINPUT29), .B(n747), .Z(n750) );
  NAND2_X1 U849 ( .A1(G171), .A2(n748), .ZN(n749) );
  NAND2_X1 U850 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U851 ( .A1(n752), .A2(n511), .ZN(n767) );
  AND2_X1 U852 ( .A1(G286), .A2(G8), .ZN(n753) );
  NAND2_X1 U853 ( .A1(n767), .A2(n753), .ZN(n763) );
  INV_X1 U854 ( .A(G8), .ZN(n761) );
  NOR2_X1 U855 ( .A1(G2090), .A2(n754), .ZN(n755) );
  XOR2_X1 U856 ( .A(KEYINPUT95), .B(n755), .Z(n757) );
  NOR2_X1 U857 ( .A1(G1971), .A2(n781), .ZN(n756) );
  NOR2_X1 U858 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U859 ( .A(n758), .B(KEYINPUT96), .ZN(n759) );
  NAND2_X1 U860 ( .A1(n759), .A2(G303), .ZN(n760) );
  OR2_X1 U861 ( .A1(n761), .A2(n760), .ZN(n762) );
  AND2_X1 U862 ( .A1(n763), .A2(n762), .ZN(n765) );
  XOR2_X1 U863 ( .A(KEYINPUT97), .B(KEYINPUT32), .Z(n764) );
  XNOR2_X1 U864 ( .A(n765), .B(n764), .ZN(n786) );
  NAND2_X1 U865 ( .A1(G8), .A2(n766), .ZN(n770) );
  AND2_X1 U866 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U867 ( .A1(n770), .A2(n769), .ZN(n784) );
  NAND2_X1 U868 ( .A1(n786), .A2(n784), .ZN(n773) );
  NOR2_X1 U869 ( .A1(G2090), .A2(G303), .ZN(n771) );
  NAND2_X1 U870 ( .A1(G8), .A2(n771), .ZN(n772) );
  NAND2_X1 U871 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U872 ( .A1(n781), .A2(n774), .ZN(n775) );
  XNOR2_X1 U873 ( .A(n775), .B(KEYINPUT98), .ZN(n779) );
  NOR2_X1 U874 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U875 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  OR2_X1 U876 ( .A1(n781), .A2(n777), .ZN(n778) );
  AND2_X1 U877 ( .A1(n779), .A2(n778), .ZN(n797) );
  XOR2_X1 U878 ( .A(G1981), .B(G305), .Z(n935) );
  NOR2_X1 U879 ( .A1(G1976), .A2(G288), .ZN(n788) );
  NAND2_X1 U880 ( .A1(n788), .A2(KEYINPUT33), .ZN(n780) );
  NOR2_X1 U881 ( .A1(n781), .A2(n780), .ZN(n794) );
  NAND2_X1 U882 ( .A1(G1976), .A2(G288), .ZN(n930) );
  INV_X1 U883 ( .A(n930), .ZN(n782) );
  OR2_X1 U884 ( .A1(n782), .A2(n781), .ZN(n789) );
  INV_X1 U885 ( .A(n789), .ZN(n783) );
  AND2_X1 U886 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U887 ( .A1(n786), .A2(n785), .ZN(n791) );
  NOR2_X1 U888 ( .A1(G1971), .A2(G303), .ZN(n787) );
  NOR2_X1 U889 ( .A1(n788), .A2(n787), .ZN(n931) );
  OR2_X1 U890 ( .A1(n789), .A2(n931), .ZN(n790) );
  NAND2_X1 U891 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U892 ( .A1(KEYINPUT33), .A2(n792), .ZN(n793) );
  NOR2_X1 U893 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U894 ( .A1(n935), .A2(n795), .ZN(n796) );
  NAND2_X1 U895 ( .A1(n797), .A2(n796), .ZN(n806) );
  XNOR2_X1 U896 ( .A(G1986), .B(KEYINPUT86), .ZN(n798) );
  XNOR2_X1 U897 ( .A(n798), .B(G290), .ZN(n953) );
  NAND2_X1 U898 ( .A1(n953), .A2(n799), .ZN(n800) );
  XOR2_X1 U899 ( .A(KEYINPUT87), .B(n800), .Z(n801) );
  AND2_X1 U900 ( .A1(n802), .A2(n801), .ZN(n803) );
  AND2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U903 ( .A(KEYINPUT99), .B(n807), .Z(n808) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n811) );
  XOR2_X1 U905 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n810) );
  XNOR2_X1 U906 ( .A(n811), .B(n810), .ZN(G329) );
  NAND2_X1 U907 ( .A1(G2106), .A2(n812), .ZN(G217) );
  INV_X1 U908 ( .A(G661), .ZN(n814) );
  NAND2_X1 U909 ( .A1(G2), .A2(G15), .ZN(n813) );
  NOR2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n815) );
  XOR2_X1 U911 ( .A(KEYINPUT104), .B(n815), .Z(G259) );
  NAND2_X1 U912 ( .A1(G3), .A2(G1), .ZN(n816) );
  NAND2_X1 U913 ( .A1(n817), .A2(n816), .ZN(G188) );
  INV_X1 U914 ( .A(n818), .ZN(G319) );
  XOR2_X1 U915 ( .A(G2096), .B(KEYINPUT43), .Z(n820) );
  XNOR2_X1 U916 ( .A(G2090), .B(G2678), .ZN(n819) );
  XNOR2_X1 U917 ( .A(n820), .B(n819), .ZN(n821) );
  XOR2_X1 U918 ( .A(n821), .B(KEYINPUT106), .Z(n823) );
  XNOR2_X1 U919 ( .A(G2067), .B(G2072), .ZN(n822) );
  XNOR2_X1 U920 ( .A(n823), .B(n822), .ZN(n827) );
  XOR2_X1 U921 ( .A(KEYINPUT42), .B(G2100), .Z(n825) );
  XNOR2_X1 U922 ( .A(G2084), .B(G2078), .ZN(n824) );
  XNOR2_X1 U923 ( .A(n825), .B(n824), .ZN(n826) );
  XNOR2_X1 U924 ( .A(n827), .B(n826), .ZN(G227) );
  XOR2_X1 U925 ( .A(G1966), .B(G1971), .Z(n829) );
  XNOR2_X1 U926 ( .A(G1986), .B(G1976), .ZN(n828) );
  XNOR2_X1 U927 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U928 ( .A(G1956), .B(G1981), .Z(n831) );
  XNOR2_X1 U929 ( .A(G1996), .B(G1991), .ZN(n830) );
  XNOR2_X1 U930 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U931 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U932 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n835), .B(n834), .ZN(n836) );
  XNOR2_X1 U934 ( .A(G2474), .B(n836), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n837), .B(n1003), .ZN(G229) );
  NAND2_X1 U936 ( .A1(G112), .A2(n858), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n838), .B(KEYINPUT110), .ZN(n841) );
  NAND2_X1 U938 ( .A1(G136), .A2(n862), .ZN(n839) );
  XOR2_X1 U939 ( .A(KEYINPUT109), .B(n839), .Z(n840) );
  NAND2_X1 U940 ( .A1(n841), .A2(n840), .ZN(n847) );
  NAND2_X1 U941 ( .A1(G124), .A2(n857), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n842), .B(KEYINPUT44), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n843), .B(KEYINPUT108), .ZN(n845) );
  NAND2_X1 U944 ( .A1(G100), .A2(n861), .ZN(n844) );
  NAND2_X1 U945 ( .A1(n845), .A2(n844), .ZN(n846) );
  NOR2_X1 U946 ( .A1(n847), .A2(n846), .ZN(G162) );
  XOR2_X1 U947 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n849) );
  XNOR2_X1 U948 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n875) );
  NAND2_X1 U950 ( .A1(G103), .A2(n861), .ZN(n851) );
  NAND2_X1 U951 ( .A1(G139), .A2(n862), .ZN(n850) );
  NAND2_X1 U952 ( .A1(n851), .A2(n850), .ZN(n856) );
  NAND2_X1 U953 ( .A1(G127), .A2(n857), .ZN(n853) );
  NAND2_X1 U954 ( .A1(G115), .A2(n858), .ZN(n852) );
  NAND2_X1 U955 ( .A1(n853), .A2(n852), .ZN(n854) );
  XOR2_X1 U956 ( .A(KEYINPUT47), .B(n854), .Z(n855) );
  NOR2_X1 U957 ( .A1(n856), .A2(n855), .ZN(n963) );
  XNOR2_X1 U958 ( .A(n963), .B(n968), .ZN(n869) );
  NAND2_X1 U959 ( .A1(G130), .A2(n857), .ZN(n860) );
  NAND2_X1 U960 ( .A1(G118), .A2(n858), .ZN(n859) );
  NAND2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n867) );
  NAND2_X1 U962 ( .A1(G106), .A2(n861), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G142), .A2(n862), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U965 ( .A(KEYINPUT45), .B(n865), .Z(n866) );
  NOR2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U968 ( .A(n871), .B(n870), .ZN(n873) );
  XNOR2_X1 U969 ( .A(G160), .B(G164), .ZN(n872) );
  XNOR2_X1 U970 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U971 ( .A(n875), .B(n874), .ZN(n878) );
  XNOR2_X1 U972 ( .A(n876), .B(G162), .ZN(n877) );
  XNOR2_X1 U973 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U974 ( .A(n880), .B(n879), .Z(n881) );
  NOR2_X1 U975 ( .A1(G37), .A2(n881), .ZN(n882) );
  XOR2_X1 U976 ( .A(KEYINPUT113), .B(n882), .Z(G395) );
  XNOR2_X1 U977 ( .A(n883), .B(KEYINPUT114), .ZN(n886) );
  XNOR2_X1 U978 ( .A(G171), .B(n884), .ZN(n885) );
  XNOR2_X1 U979 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U980 ( .A(n887), .B(G286), .Z(n888) );
  NOR2_X1 U981 ( .A1(G37), .A2(n888), .ZN(G397) );
  XOR2_X1 U982 ( .A(G2451), .B(G2430), .Z(n890) );
  XNOR2_X1 U983 ( .A(G2438), .B(G2443), .ZN(n889) );
  XNOR2_X1 U984 ( .A(n890), .B(n889), .ZN(n896) );
  XOR2_X1 U985 ( .A(G2435), .B(G2454), .Z(n892) );
  XNOR2_X1 U986 ( .A(G1341), .B(G1348), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n892), .B(n891), .ZN(n894) );
  XOR2_X1 U988 ( .A(G2446), .B(G2427), .Z(n893) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U990 ( .A(n896), .B(n895), .Z(n897) );
  NAND2_X1 U991 ( .A1(G14), .A2(n897), .ZN(n906) );
  NAND2_X1 U992 ( .A1(G319), .A2(n906), .ZN(n900) );
  NOR2_X1 U993 ( .A1(G227), .A2(G229), .ZN(n898) );
  XNOR2_X1 U994 ( .A(KEYINPUT49), .B(n898), .ZN(n899) );
  NOR2_X1 U995 ( .A1(n900), .A2(n899), .ZN(n902) );
  NOR2_X1 U996 ( .A1(G395), .A2(G397), .ZN(n901) );
  NAND2_X1 U997 ( .A1(n902), .A2(n901), .ZN(G225) );
  XNOR2_X1 U998 ( .A(KEYINPUT115), .B(G225), .ZN(G308) );
  INV_X1 U1000 ( .A(G120), .ZN(G236) );
  INV_X1 U1001 ( .A(G96), .ZN(G221) );
  INV_X1 U1002 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1003 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n905), .B(KEYINPUT105), .ZN(G261) );
  INV_X1 U1005 ( .A(G261), .ZN(G325) );
  INV_X1 U1006 ( .A(G108), .ZN(G238) );
  INV_X1 U1007 ( .A(n906), .ZN(G401) );
  XOR2_X1 U1008 ( .A(G1991), .B(G25), .Z(n907) );
  NAND2_X1 U1009 ( .A1(n907), .A2(G28), .ZN(n916) );
  XNOR2_X1 U1010 ( .A(G1996), .B(G32), .ZN(n909) );
  XNOR2_X1 U1011 ( .A(G33), .B(G2072), .ZN(n908) );
  NOR2_X1 U1012 ( .A1(n909), .A2(n908), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(G2067), .B(G26), .ZN(n912) );
  XNOR2_X1 U1014 ( .A(G27), .B(n910), .ZN(n911) );
  NOR2_X1 U1015 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1016 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1018 ( .A(KEYINPUT119), .B(n917), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(n918), .B(KEYINPUT53), .ZN(n922) );
  XOR2_X1 U1020 ( .A(G34), .B(KEYINPUT120), .Z(n920) );
  XNOR2_X1 U1021 ( .A(G2084), .B(KEYINPUT54), .ZN(n919) );
  XNOR2_X1 U1022 ( .A(n920), .B(n919), .ZN(n921) );
  NAND2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(G35), .B(G2090), .ZN(n923) );
  NOR2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1026 ( .A(KEYINPUT121), .B(n925), .Z(n926) );
  NOR2_X1 U1027 ( .A1(G29), .A2(n926), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(KEYINPUT55), .B(n927), .ZN(n928) );
  NAND2_X1 U1029 ( .A1(n928), .A2(G11), .ZN(n958) );
  XOR2_X1 U1030 ( .A(G16), .B(KEYINPUT122), .Z(n929) );
  XNOR2_X1 U1031 ( .A(KEYINPUT56), .B(n929), .ZN(n955) );
  AND2_X1 U1032 ( .A1(G303), .A2(G1971), .ZN(n933) );
  NAND2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1035 ( .A(KEYINPUT124), .B(n934), .Z(n946) );
  XNOR2_X1 U1036 ( .A(G1966), .B(G168), .ZN(n936) );
  NAND2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1038 ( .A(KEYINPUT57), .B(n937), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(n938), .B(G1956), .ZN(n939) );
  XNOR2_X1 U1040 ( .A(n939), .B(KEYINPUT123), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(G1341), .B(n940), .ZN(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n951) );
  XOR2_X1 U1045 ( .A(G171), .B(G1961), .Z(n949) );
  XNOR2_X1 U1046 ( .A(n947), .B(G1348), .ZN(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1051 ( .A(KEYINPUT125), .B(n956), .Z(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n986) );
  XOR2_X1 U1053 ( .A(G2090), .B(G162), .Z(n959) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(KEYINPUT117), .B(n961), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(n962), .B(KEYINPUT51), .ZN(n982) );
  XNOR2_X1 U1057 ( .A(G164), .B(G2078), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(G2072), .B(n963), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(n964), .B(KEYINPUT118), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(n967), .B(KEYINPUT50), .ZN(n980) );
  NOR2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n973) );
  XOR2_X1 U1063 ( .A(G160), .B(G2084), .Z(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(n976), .B(KEYINPUT116), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1070 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1071 ( .A(KEYINPUT52), .B(n983), .ZN(n984) );
  NAND2_X1 U1072 ( .A1(n984), .A2(G29), .ZN(n985) );
  NAND2_X1 U1073 ( .A1(n986), .A2(n985), .ZN(n1011) );
  XOR2_X1 U1074 ( .A(G1976), .B(G23), .Z(n990) );
  XNOR2_X1 U1075 ( .A(G1986), .B(G24), .ZN(n988) );
  XNOR2_X1 U1076 ( .A(G1971), .B(G22), .ZN(n987) );
  NOR2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(KEYINPUT58), .B(n991), .ZN(n1007) );
  XNOR2_X1 U1080 ( .A(G1348), .B(KEYINPUT59), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(n992), .B(G4), .ZN(n996) );
  XNOR2_X1 U1082 ( .A(G1981), .B(G6), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(G1341), .B(G19), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(G20), .B(G1956), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1088 ( .A(KEYINPUT60), .B(n999), .Z(n1001) );
  XNOR2_X1 U1089 ( .A(G1966), .B(G21), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(KEYINPUT126), .B(n1002), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(n1003), .B(G5), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1095 ( .A(KEYINPUT61), .B(n1008), .Z(n1009) );
  NOR2_X1 U1096 ( .A1(G16), .A2(n1009), .ZN(n1010) );
  NOR2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(n1012), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1099 ( .A(G311), .ZN(G150) );
endmodule

