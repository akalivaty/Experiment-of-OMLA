//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT99), .ZN(new_n203));
  NAND2_X1  g002(.A1(G71gat), .A2(G78gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT9), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n202), .A2(new_n203), .A3(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G71gat), .B(G78gat), .Z(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G231gat), .A2(G233gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G127gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT16), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n216), .B1(new_n217), .B2(G1gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(G1gat), .B2(new_n216), .ZN(new_n219));
  XOR2_X1   g018(.A(new_n219), .B(G8gat), .Z(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(new_n210), .B2(new_n209), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n215), .B(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n223));
  INV_X1    g022(.A(G155gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G183gat), .B(G211gat), .ZN(new_n226));
  XOR2_X1   g025(.A(new_n225), .B(new_n226), .Z(new_n227));
  OR2_X1    g026(.A1(new_n222), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n222), .A2(new_n227), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G232gat), .ZN(new_n231));
  INV_X1    g030(.A(G233gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(KEYINPUT41), .ZN(new_n234));
  XNOR2_X1  g033(.A(G134gat), .B(G162gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT100), .ZN(new_n238));
  INV_X1    g037(.A(G85gat), .ZN(new_n239));
  INV_X1    g038(.A(G92gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(KEYINPUT100), .A2(G85gat), .A3(G92gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(KEYINPUT7), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT7), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n238), .B(new_n244), .C1(new_n239), .C2(new_n240), .ZN(new_n245));
  NAND2_X1  g044(.A1(G99gat), .A2(G106gat), .ZN(new_n246));
  AOI22_X1  g045(.A1(KEYINPUT8), .A2(new_n246), .B1(new_n239), .B2(new_n240), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n243), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  OR2_X1    g047(.A1(G99gat), .A2(G106gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n246), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n243), .A2(new_n251), .A3(new_n245), .A4(new_n247), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G43gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(G50gat), .ZN(new_n255));
  INV_X1    g054(.A(G50gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(G43gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n258), .A2(KEYINPUT94), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT15), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT94), .ZN(new_n261));
  NOR3_X1   g060(.A1(new_n255), .A2(new_n257), .A3(new_n261), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G29gat), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n264), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT14), .B(G29gat), .ZN(new_n266));
  INV_X1    g065(.A(G36gat), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT95), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n256), .A2(G43gat), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n257), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(new_n271), .B2(new_n272), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n268), .B1(new_n274), .B2(new_n260), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n270), .B1(new_n263), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT17), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT96), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n277), .A2(KEYINPUT96), .ZN(new_n280));
  OAI221_X1 g079(.A(new_n253), .B1(KEYINPUT17), .B2(new_n276), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(G190gat), .B(G218gat), .Z(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n233), .A2(KEYINPUT41), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(new_n276), .B2(new_n253), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n283), .B1(new_n281), .B2(new_n286), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n237), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n289), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(new_n236), .A3(new_n287), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n230), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n253), .A2(new_n209), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n253), .A2(new_n209), .ZN(new_n297));
  OR3_X1    g096(.A1(new_n296), .A2(new_n297), .A3(KEYINPUT10), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G230gat), .A2(G233gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n301), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(new_n296), .B2(new_n297), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G120gat), .B(G148gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(G176gat), .B(G204gat), .ZN(new_n307));
  XOR2_X1   g106(.A(new_n306), .B(new_n307), .Z(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n302), .A2(new_n304), .A3(new_n308), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n295), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G228gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(new_n232), .ZN(new_n316));
  XOR2_X1   g115(.A(G197gat), .B(G204gat), .Z(new_n317));
  INV_X1    g116(.A(G218gat), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n318), .A2(KEYINPUT70), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(KEYINPUT70), .ZN(new_n320));
  OAI21_X1  g119(.A(G211gat), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT22), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n317), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G211gat), .B(G218gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT3), .ZN(new_n326));
  INV_X1    g125(.A(G162gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n224), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n331));
  XNOR2_X1  g130(.A(G141gat), .B(G148gat), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n330), .B(new_n331), .C1(KEYINPUT2), .C2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G148gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(G141gat), .ZN(new_n335));
  INV_X1    g134(.A(G141gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G148gat), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT2), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G155gat), .B(G162gat), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT75), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n335), .ZN(new_n342));
  AND2_X1   g141(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n342), .B1(new_n345), .B2(G148gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT2), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n328), .B1(new_n347), .B2(new_n329), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n349));
  NOR3_X1   g148(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT76), .B(G141gat), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n335), .B1(new_n351), .B2(new_n334), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n329), .A2(new_n347), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(new_n224), .B2(new_n327), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT77), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n326), .B(new_n341), .C1(new_n350), .C2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT29), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n325), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n349), .B1(new_n346), .B2(new_n348), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n352), .A2(KEYINPUT77), .A3(new_n354), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n359), .A2(new_n360), .B1(new_n340), .B2(new_n333), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT70), .B(G218gat), .ZN(new_n362));
  INV_X1    g161(.A(G211gat), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n322), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n317), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n324), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n324), .B1(new_n364), .B2(new_n365), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n357), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n361), .B1(new_n369), .B2(new_n326), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n316), .B1(new_n358), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT86), .B1(new_n323), .B2(new_n324), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT86), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT85), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n366), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n323), .A2(KEYINPUT85), .A3(new_n324), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n372), .A2(new_n374), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n357), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n361), .B1(new_n379), .B2(new_n326), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT29), .B1(new_n361), .B2(new_n326), .ZN(new_n381));
  OAI22_X1  g180(.A1(new_n381), .A2(new_n325), .B1(new_n315), .B2(new_n232), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n371), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(G22gat), .ZN(new_n384));
  INV_X1    g183(.A(G22gat), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n371), .B(new_n385), .C1(new_n380), .C2(new_n382), .ZN(new_n386));
  XNOR2_X1  g185(.A(G78gat), .B(G106gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT31), .B(G50gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n387), .B(new_n388), .Z(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n390), .A2(new_n391), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n384), .A2(new_n386), .ZN(new_n394));
  INV_X1    g193(.A(new_n389), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT88), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT88), .ZN(new_n397));
  AOI211_X1 g196(.A(new_n397), .B(new_n389), .C1(new_n384), .C2(new_n386), .ZN(new_n398));
  OAI22_X1  g197(.A1(new_n392), .A2(new_n393), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(G169gat), .A2(G176gat), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT26), .ZN(new_n403));
  INV_X1    g202(.A(G169gat), .ZN(new_n404));
  INV_X1    g203(.A(G176gat), .ZN(new_n405));
  AND4_X1   g204(.A1(KEYINPUT66), .A2(new_n403), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(G169gat), .A2(G176gat), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT66), .B1(new_n407), .B2(new_n403), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n402), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G183gat), .A2(G190gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT28), .ZN(new_n412));
  XOR2_X1   g211(.A(KEYINPUT27), .B(G183gat), .Z(new_n413));
  OAI21_X1  g212(.A(new_n412), .B1(new_n413), .B2(G190gat), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT65), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT27), .B(G183gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT65), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n412), .A2(G190gat), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n416), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n411), .B1(new_n414), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT64), .ZN(new_n422));
  AND2_X1   g221(.A1(G183gat), .A2(G190gat), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT24), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n423), .A2(new_n424), .B1(G169gat), .B2(G176gat), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT23), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n426), .A2(new_n404), .A3(new_n405), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G183gat), .B(G190gat), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n425), .B(new_n429), .C1(new_n424), .C2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT25), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n401), .B1(new_n410), .B2(KEYINPUT24), .ZN(new_n434));
  INV_X1    g233(.A(G183gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(G190gat), .ZN(new_n436));
  INV_X1    g235(.A(G190gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G183gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n434), .B1(new_n439), .B2(KEYINPUT24), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT25), .B1(new_n440), .B2(new_n429), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n422), .B1(new_n433), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n431), .A2(new_n432), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(KEYINPUT25), .A3(new_n429), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(KEYINPUT64), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n421), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(G113gat), .ZN(new_n447));
  INV_X1    g246(.A(G120gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(G113gat), .A2(G120gat), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT1), .ZN(new_n452));
  XOR2_X1   g251(.A(G127gat), .B(G134gat), .Z(new_n453));
  OAI211_X1 g252(.A(new_n451), .B(new_n452), .C1(new_n453), .C2(KEYINPUT67), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n449), .A2(new_n452), .A3(new_n450), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n449), .A2(KEYINPUT67), .A3(new_n450), .ZN(new_n456));
  XNOR2_X1  g255(.A(G127gat), .B(G134gat), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n446), .A2(new_n454), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n420), .A2(new_n414), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n460), .A2(new_n410), .A3(new_n409), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n443), .A2(KEYINPUT64), .A3(new_n444), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT64), .B1(new_n443), .B2(new_n444), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n454), .A2(new_n458), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(G227gat), .A2(G233gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n459), .A2(new_n466), .A3(G227gat), .A4(G233gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(KEYINPUT32), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT32), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n467), .A2(new_n472), .A3(new_n468), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT33), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  XOR2_X1   g275(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  XOR2_X1   g277(.A(G15gat), .B(G43gat), .Z(new_n479));
  XNOR2_X1  g278(.A(G71gat), .B(G99gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n476), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n478), .B1(new_n476), .B2(new_n481), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n474), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n476), .A2(new_n481), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n477), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n487), .A2(new_n473), .A3(new_n471), .A4(new_n482), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n399), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT35), .ZN(new_n491));
  INV_X1    g290(.A(new_n325), .ZN(new_n492));
  NAND2_X1  g291(.A1(G226gat), .A2(G233gat), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n446), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n443), .A2(new_n444), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n461), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(new_n357), .A3(new_n493), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n492), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n493), .B1(new_n446), .B2(KEYINPUT29), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT71), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT71), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n502), .B(new_n493), .C1(new_n446), .C2(KEYINPUT29), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n493), .B1(new_n461), .B2(new_n496), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n501), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n499), .B1(new_n506), .B2(new_n492), .ZN(new_n507));
  XOR2_X1   g306(.A(G8gat), .B(G36gat), .Z(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT72), .ZN(new_n509));
  XNOR2_X1  g308(.A(G64gat), .B(G92gat), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n509), .B(new_n510), .Z(new_n511));
  NAND3_X1  g310(.A1(new_n507), .A2(KEYINPUT30), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n511), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n504), .B1(new_n500), .B2(KEYINPUT71), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n325), .B1(new_n514), .B2(new_n503), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n513), .B1(new_n515), .B2(new_n499), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT73), .B1(new_n507), .B2(new_n511), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT73), .ZN(new_n519));
  NOR4_X1   g318(.A1(new_n515), .A2(new_n519), .A3(new_n499), .A4(new_n513), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(KEYINPUT74), .B(KEYINPUT30), .Z(new_n522));
  AOI21_X1  g321(.A(new_n517), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G1gat), .B(G29gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT0), .ZN(new_n525));
  XNOR2_X1  g324(.A(G57gat), .B(G85gat), .ZN(new_n526));
  XOR2_X1   g325(.A(new_n525), .B(new_n526), .Z(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT82), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n465), .B(new_n341), .C1(new_n350), .C2(new_n355), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(KEYINPUT4), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT4), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n361), .A2(KEYINPUT82), .A3(new_n532), .A4(new_n465), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n530), .A2(KEYINPUT83), .A3(KEYINPUT4), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT83), .B1(new_n530), .B2(KEYINPUT4), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT79), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT78), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n454), .A2(KEYINPUT78), .A3(new_n458), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n544), .B1(new_n361), .B2(new_n326), .ZN(new_n545));
  INV_X1    g344(.A(new_n356), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n538), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n341), .B1(new_n350), .B2(new_n355), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT3), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n549), .A2(KEYINPUT79), .A3(new_n356), .A4(new_n544), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n534), .A2(new_n537), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G225gat), .A2(G233gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(KEYINPUT5), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n528), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n553), .B1(new_n547), .B2(new_n550), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n530), .A2(KEYINPUT4), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT80), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT81), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(new_n530), .B2(KEYINPUT4), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n361), .A2(KEYINPUT81), .A3(new_n532), .A4(new_n465), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT80), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n530), .A2(new_n562), .A3(KEYINPUT4), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n558), .A2(new_n560), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n556), .A2(new_n564), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n542), .A2(new_n543), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n530), .B1(new_n566), .B2(new_n361), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n553), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT5), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT6), .B1(new_n555), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n569), .B1(new_n556), .B2(new_n564), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n547), .A2(new_n550), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT83), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n530), .A2(KEYINPUT83), .A3(KEYINPUT4), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n576), .A2(new_n531), .A3(new_n533), .A4(new_n577), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n574), .A2(new_n578), .A3(new_n554), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n528), .B1(new_n573), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n572), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT84), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT6), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n582), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n551), .A2(new_n554), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n571), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n586), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(new_n528), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n581), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n490), .A2(new_n491), .A3(new_n523), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n506), .A2(new_n492), .ZN(new_n590));
  INV_X1    g389(.A(new_n499), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n519), .B1(new_n592), .B2(new_n513), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n507), .A2(KEYINPUT73), .A3(new_n511), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n594), .A3(new_n522), .ZN(new_n595));
  INV_X1    g394(.A(new_n517), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n399), .A2(new_n595), .A3(new_n596), .A4(new_n489), .ZN(new_n597));
  INV_X1    g396(.A(new_n588), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT35), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n589), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT40), .ZN(new_n601));
  OAI21_X1  g400(.A(KEYINPUT39), .B1(new_n567), .B2(new_n553), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n602), .B(KEYINPUT89), .Z(new_n603));
  AOI21_X1  g402(.A(new_n552), .B1(new_n574), .B2(new_n578), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n528), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n601), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n607), .B(KEYINPUT40), .C1(new_n603), .C2(new_n604), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(new_n610), .A3(new_n580), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n399), .B1(new_n523), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n499), .A2(KEYINPUT37), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n511), .B1(new_n590), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT37), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n614), .B1(new_n615), .B2(new_n507), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT38), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n494), .B1(new_n464), .B2(new_n357), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n505), .B1(new_n619), .B2(new_n502), .ZN(new_n620));
  INV_X1    g419(.A(new_n503), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n325), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n495), .A2(new_n498), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n615), .B1(new_n623), .B2(new_n492), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT38), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n572), .A2(new_n580), .B1(new_n614), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n626), .A2(new_n521), .A3(new_n587), .A4(new_n584), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT90), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n618), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n584), .A2(new_n587), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n630), .A2(KEYINPUT90), .A3(new_n521), .A4(new_n626), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n612), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n523), .A2(new_n588), .ZN(new_n633));
  INV_X1    g432(.A(new_n399), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT69), .B(KEYINPUT36), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n489), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT69), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n489), .B1(new_n638), .B2(KEYINPUT36), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n600), .B1(new_n632), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n220), .ZN(new_n643));
  INV_X1    g442(.A(new_n276), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT17), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n279), .B2(new_n280), .ZN(new_n647));
  NAND2_X1  g446(.A1(G229gat), .A2(G233gat), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n276), .A2(new_n220), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT97), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT18), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n647), .A2(new_n650), .A3(KEYINPUT18), .A4(new_n648), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n276), .A2(new_n220), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n648), .B(KEYINPUT13), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n653), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G113gat), .B(G141gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT92), .ZN(new_n661));
  XNOR2_X1  g460(.A(G169gat), .B(G197gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT12), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n659), .A2(KEYINPUT93), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n666), .B1(new_n659), .B2(KEYINPUT93), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n642), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT98), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n642), .A2(KEYINPUT98), .A3(new_n669), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n314), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n598), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g475(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n677));
  NAND2_X1  g476(.A1(new_n595), .A2(new_n596), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT16), .B(G8gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT102), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n677), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(G8gat), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n682), .B(new_n683), .C1(new_n679), .C2(new_n685), .ZN(G1325gat));
  INV_X1    g485(.A(new_n640), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n674), .A2(G15gat), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(G15gat), .B1(new_n674), .B2(new_n489), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(KEYINPUT103), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691));
  AOI211_X1 g490(.A(new_n691), .B(G15gat), .C1(new_n674), .C2(new_n489), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n688), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g494(.A(KEYINPUT104), .B(new_n688), .C1(new_n690), .C2(new_n692), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(G1326gat));
  NAND2_X1  g496(.A1(new_n674), .A2(new_n634), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT43), .B(G22gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  NAND2_X1  g499(.A1(new_n672), .A2(new_n673), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n230), .A2(new_n313), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n293), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n264), .A3(new_n598), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT45), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n642), .A2(new_n294), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT44), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n709), .B1(new_n632), .B2(new_n641), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n614), .A2(new_n625), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n581), .A2(new_n593), .A3(new_n711), .A4(new_n594), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n584), .A2(new_n587), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n628), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(new_n631), .A3(new_n617), .ZN(new_n715));
  INV_X1    g514(.A(new_n611), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n634), .B1(new_n716), .B2(new_n678), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n633), .A2(new_n634), .B1(new_n637), .B2(new_n639), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n718), .A2(KEYINPUT105), .A3(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n589), .A2(new_n599), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n600), .A2(KEYINPUT106), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n710), .A2(new_n720), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n293), .A2(KEYINPUT44), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n725), .B1(new_n724), .B2(new_n726), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n708), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n659), .A2(KEYINPUT93), .ZN(new_n731));
  INV_X1    g530(.A(new_n666), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n659), .A2(KEYINPUT93), .A3(new_n666), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n702), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n730), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G29gat), .B1(new_n737), .B2(new_n588), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n706), .A2(new_n738), .ZN(G1328gat));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n523), .A2(G36gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n704), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n701), .A2(new_n703), .A3(new_n742), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT108), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n740), .B1(new_n746), .B2(KEYINPUT46), .ZN(new_n747));
  OAI21_X1  g546(.A(G36gat), .B1(new_n737), .B2(new_n523), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(KEYINPUT46), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT46), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n743), .A2(KEYINPUT109), .A3(new_n750), .A4(new_n745), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n747), .A2(new_n748), .A3(new_n749), .A4(new_n751), .ZN(G1329gat));
  NAND4_X1  g551(.A1(new_n730), .A2(G43gat), .A3(new_n687), .A4(new_n736), .ZN(new_n753));
  OR2_X1    g552(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n701), .A2(new_n489), .A3(new_n703), .ZN(new_n755));
  AOI22_X1  g554(.A1(new_n755), .A2(new_n254), .B1(KEYINPUT110), .B2(KEYINPUT47), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n754), .B1(new_n753), .B2(new_n756), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(G1330gat));
  NAND2_X1  g558(.A1(new_n704), .A2(new_n634), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n256), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n634), .A2(G50gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n737), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT48), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT48), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n761), .B(new_n765), .C1(new_n737), .C2(new_n762), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1331gat));
  NAND3_X1  g566(.A1(new_n295), .A2(new_n735), .A3(new_n312), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n724), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n598), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g572(.A(new_n523), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT111), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n776), .B(new_n777), .Z(G1333gat));
  OAI21_X1  g577(.A(G71gat), .B1(new_n770), .B2(new_n640), .ZN(new_n779));
  INV_X1    g578(.A(new_n489), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n780), .A2(G71gat), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n770), .B2(new_n781), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n782), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g582(.A1(new_n771), .A2(new_n634), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g584(.A1(new_n735), .A2(new_n230), .A3(new_n312), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n724), .A2(new_n726), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT107), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n727), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n786), .B1(new_n789), .B2(new_n708), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n790), .A2(new_n598), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n724), .A2(new_n735), .A3(new_n230), .A4(new_n294), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT51), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n598), .A2(new_n239), .A3(new_n312), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT112), .ZN(new_n795));
  OAI22_X1  g594(.A1(new_n791), .A2(new_n239), .B1(new_n793), .B2(new_n795), .ZN(G1336gat));
  AOI21_X1  g595(.A(new_n240), .B1(new_n790), .B2(new_n678), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n678), .A2(new_n240), .A3(new_n312), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT52), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n793), .A2(new_n798), .ZN(new_n801));
  INV_X1    g600(.A(new_n786), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n730), .A2(new_n678), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G92gat), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n801), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n800), .A2(new_n806), .ZN(G1337gat));
  NAND3_X1  g606(.A1(new_n730), .A2(new_n687), .A3(new_n802), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G99gat), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n808), .A2(new_n809), .ZN(new_n812));
  OR3_X1    g611(.A1(new_n780), .A2(G99gat), .A3(new_n313), .ZN(new_n813));
  OAI22_X1  g612(.A1(new_n811), .A2(new_n812), .B1(new_n793), .B2(new_n813), .ZN(G1338gat));
  INV_X1    g613(.A(G106gat), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n790), .B2(new_n634), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n634), .A2(new_n815), .A3(new_n312), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n793), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT53), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n793), .A2(new_n817), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n730), .A2(new_n634), .A3(new_n802), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G106gat), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n820), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n819), .A2(new_n824), .ZN(G1339gat));
  NAND3_X1  g624(.A1(new_n295), .A2(new_n735), .A3(new_n313), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n298), .A2(new_n299), .A3(new_n303), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n302), .A2(KEYINPUT54), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n303), .B1(new_n298), .B2(new_n299), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n308), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT55), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n828), .A2(KEYINPUT55), .A3(new_n831), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n311), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(KEYINPUT114), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(new_n836), .B2(new_n311), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n834), .B(new_n835), .C1(new_n838), .C2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n653), .A2(new_n654), .A3(new_n658), .A4(new_n666), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n656), .A2(new_n657), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n648), .B1(new_n647), .B2(new_n650), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n665), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n292), .A3(new_n290), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n841), .A2(new_n847), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n842), .A2(new_n312), .A3(new_n845), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(new_n841), .B2(new_n735), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n848), .B1(new_n851), .B2(new_n293), .ZN(new_n852));
  INV_X1    g651(.A(new_n230), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n826), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  OR3_X1    g654(.A1(new_n855), .A2(KEYINPUT116), .A3(new_n634), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT116), .B1(new_n855), .B2(new_n634), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n523), .A2(new_n598), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n859), .A2(new_n780), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(G113gat), .B1(new_n861), .B2(new_n735), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n855), .A2(new_n588), .A3(new_n597), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT117), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n447), .A3(new_n669), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n862), .A2(new_n865), .ZN(G1340gat));
  OAI21_X1  g665(.A(G120gat), .B1(new_n861), .B2(new_n313), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n864), .A2(new_n448), .A3(new_n312), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1341gat));
  NAND4_X1  g668(.A1(new_n858), .A2(G127gat), .A3(new_n853), .A4(new_n860), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n870), .A2(KEYINPUT118), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(KEYINPUT118), .ZN(new_n872));
  AOI21_X1  g671(.A(G127gat), .B1(new_n863), .B2(new_n853), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(G1342gat));
  NOR2_X1   g673(.A1(new_n293), .A2(G134gat), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT56), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n863), .B(new_n875), .C1(KEYINPUT120), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n863), .A2(new_n875), .ZN(new_n878));
  XOR2_X1   g677(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n858), .A2(new_n294), .A3(new_n860), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n881), .A2(new_n882), .A3(G134gat), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n881), .B2(G134gat), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n877), .B(new_n880), .C1(new_n883), .C2(new_n884), .ZN(G1343gat));
  NOR2_X1   g684(.A1(new_n687), .A2(new_n859), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT121), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n634), .A2(KEYINPUT57), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n838), .A2(new_n840), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n834), .A2(new_n835), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n889), .A2(new_n890), .A3(new_n294), .A4(new_n846), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n837), .A2(new_n832), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n733), .A2(new_n892), .A3(new_n734), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n294), .B1(new_n893), .B2(new_n850), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n849), .B1(new_n669), .B2(new_n892), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n897), .A2(KEYINPUT122), .A3(new_n294), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n230), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n888), .B1(new_n899), .B2(new_n826), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT57), .B1(new_n854), .B2(new_n634), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n887), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n351), .B1(new_n902), .B2(new_n735), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT58), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n855), .A2(new_n588), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n687), .A2(new_n399), .A3(new_n678), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n669), .A2(new_n336), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n903), .B(new_n904), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n902), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g711(.A(KEYINPUT123), .B(new_n887), .C1(new_n900), .C2(new_n901), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n669), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n910), .B1(new_n914), .B2(new_n351), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n909), .B1(new_n915), .B2(new_n904), .ZN(G1344gat));
  NOR3_X1   g715(.A1(new_n907), .A2(G148gat), .A3(new_n313), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n891), .B(KEYINPUT124), .C1(new_n897), .C2(new_n294), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n919), .B1(new_n894), .B2(new_n848), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n918), .A2(new_n920), .A3(new_n230), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n399), .B1(new_n921), .B2(new_n826), .ZN(new_n922));
  OAI22_X1  g721(.A1(new_n922), .A2(KEYINPUT57), .B1(new_n855), .B2(new_n888), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n312), .A3(new_n887), .ZN(new_n924));
  AND2_X1   g723(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n917), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n912), .A2(new_n913), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n334), .B1(new_n927), .B2(new_n312), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n926), .B1(new_n928), .B2(KEYINPUT59), .ZN(G1345gat));
  INV_X1    g728(.A(new_n907), .ZN(new_n930));
  AOI21_X1  g729(.A(G155gat), .B1(new_n930), .B2(new_n853), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n853), .A2(G155gat), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT125), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n931), .B1(new_n927), .B2(new_n933), .ZN(G1346gat));
  AOI21_X1  g733(.A(G162gat), .B1(new_n930), .B2(new_n294), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n293), .A2(new_n327), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n927), .B2(new_n936), .ZN(G1347gat));
  NOR2_X1   g736(.A1(new_n855), .A2(new_n598), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n634), .A2(new_n523), .A3(new_n780), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(G169gat), .B1(new_n941), .B2(new_n669), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n678), .A2(new_n588), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT126), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(new_n780), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n946), .B1(new_n856), .B2(new_n857), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n735), .A2(new_n404), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n942), .B1(new_n947), .B2(new_n948), .ZN(G1348gat));
  AOI21_X1  g748(.A(new_n405), .B1(new_n947), .B2(new_n312), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n940), .A2(G176gat), .A3(new_n313), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n950), .A2(new_n951), .ZN(G1349gat));
  AOI21_X1  g751(.A(new_n435), .B1(new_n947), .B2(new_n853), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n416), .A2(new_n418), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n940), .A2(new_n954), .A3(new_n230), .ZN(new_n955));
  OR3_X1    g754(.A1(new_n953), .A2(KEYINPUT60), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(KEYINPUT60), .B1(new_n953), .B2(new_n955), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1350gat));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n437), .A3(new_n294), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n947), .A2(new_n294), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n960), .B1(new_n961), .B2(G190gat), .ZN(new_n962));
  AOI211_X1 g761(.A(KEYINPUT61), .B(new_n437), .C1(new_n947), .C2(new_n294), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(G1351gat));
  AND4_X1   g763(.A1(new_n634), .A2(new_n938), .A3(new_n678), .A4(new_n640), .ZN(new_n965));
  AOI21_X1  g764(.A(G197gat), .B1(new_n965), .B2(new_n669), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n944), .A2(new_n687), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n923), .A2(new_n967), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n669), .A2(G197gat), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(G1352gat));
  INV_X1    g769(.A(G204gat), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n965), .A2(new_n971), .A3(new_n312), .ZN(new_n972));
  OR2_X1    g771(.A1(new_n972), .A2(KEYINPUT62), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(KEYINPUT62), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n968), .A2(new_n312), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n973), .B(new_n974), .C1(new_n971), .C2(new_n975), .ZN(G1353gat));
  NAND3_X1  g775(.A1(new_n965), .A2(new_n363), .A3(new_n853), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT127), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n923), .A2(new_n978), .A3(new_n853), .A4(new_n967), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n979), .A2(G211gat), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n923), .A2(new_n853), .A3(new_n967), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(KEYINPUT127), .ZN(new_n982));
  AOI21_X1  g781(.A(KEYINPUT63), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  AND4_X1   g782(.A1(KEYINPUT63), .A2(new_n982), .A3(G211gat), .A4(new_n979), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n977), .B1(new_n983), .B2(new_n984), .ZN(G1354gat));
  AOI21_X1  g784(.A(G218gat), .B1(new_n965), .B2(new_n294), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n293), .A2(new_n362), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n986), .B1(new_n968), .B2(new_n987), .ZN(G1355gat));
endmodule


