//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(KEYINPUT64), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT64), .A2(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(G143), .A3(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT64), .A2(G146), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT64), .A2(G146), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n188), .A2(G143), .ZN(new_n197));
  AOI22_X1  g011(.A1(new_n192), .A2(G128), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT65), .B1(new_n188), .B2(G143), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n191), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n189), .A2(new_n205), .A3(G143), .A4(new_n190), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n201), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT11), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G137), .ZN(new_n210));
  INV_X1    g024(.A(G137), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT11), .A3(G134), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(G137), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n210), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n209), .A2(G137), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n211), .A2(G134), .ZN(new_n217));
  OAI21_X1  g031(.A(G131), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n215), .A2(new_n218), .A3(KEYINPUT68), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT68), .B1(new_n215), .B2(new_n218), .ZN(new_n220));
  OAI22_X1  g034(.A1(new_n198), .A2(new_n207), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n196), .A2(new_n197), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n194), .A2(new_n195), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G143), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n224), .B1(new_n227), .B2(new_n199), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n202), .B1(new_n226), .B2(G143), .ZN(new_n229));
  INV_X1    g043(.A(new_n206), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n200), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n215), .A2(new_n218), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n215), .A2(new_n218), .A3(KEYINPUT68), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n232), .A2(new_n237), .A3(KEYINPUT69), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n204), .A2(new_n206), .ZN(new_n239));
  AND2_X1   g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  NOR2_X1   g054(.A1(KEYINPUT0), .A2(G128), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n239), .A2(new_n240), .B1(new_n224), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n210), .A2(new_n212), .A3(new_n214), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G131), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n215), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n223), .A2(KEYINPUT30), .A3(new_n238), .A4(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT30), .ZN(new_n249));
  INV_X1    g063(.A(new_n233), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n250), .B1(new_n198), .B2(new_n207), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n240), .B1(new_n229), .B2(new_n230), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n224), .A2(new_n242), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n252), .A2(KEYINPUT66), .A3(new_n246), .A4(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT66), .B1(new_n243), .B2(new_n246), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n249), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G119), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n258), .A2(G116), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT67), .B(G116), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(G119), .ZN(new_n261));
  XOR2_X1   g075(.A(KEYINPUT2), .B(G113), .Z(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n248), .A2(new_n257), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n263), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n223), .A2(new_n265), .A3(new_n238), .A4(new_n247), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  OR2_X1    g081(.A1(KEYINPUT70), .A2(G237), .ZN(new_n268));
  NAND2_X1  g082(.A1(KEYINPUT70), .A2(G237), .ZN(new_n269));
  AOI21_X1  g083(.A(G953), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G210), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT26), .B(G101), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n273), .B(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT29), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n263), .B1(new_n255), .B2(new_n256), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n266), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT72), .B(KEYINPUT28), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n247), .A2(new_n221), .A3(new_n265), .ZN(new_n281));
  OAI22_X1  g095(.A1(new_n279), .A2(new_n280), .B1(KEYINPUT28), .B2(new_n281), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n276), .B(new_n277), .C1(new_n282), .C2(new_n275), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n281), .A2(KEYINPUT28), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n266), .A2(KEYINPUT74), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n223), .A2(new_n247), .A3(new_n238), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n263), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n221), .A2(new_n222), .B1(new_n246), .B2(new_n243), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n265), .A4(new_n238), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n285), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n284), .B1(new_n291), .B2(KEYINPUT28), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n275), .A2(new_n277), .ZN(new_n293));
  AOI21_X1  g107(.A(G902), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n283), .B1(new_n294), .B2(KEYINPUT75), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n296));
  AOI211_X1 g110(.A(new_n296), .B(G902), .C1(new_n292), .C2(new_n293), .ZN(new_n297));
  OAI21_X1  g111(.A(G472), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n275), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n264), .A2(new_n299), .A3(new_n266), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT31), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n264), .A2(KEYINPUT31), .A3(new_n299), .A4(new_n266), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n282), .A2(new_n275), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(G472), .A2(G902), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(KEYINPUT73), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n302), .A2(new_n303), .B1(new_n282), .B2(new_n275), .ZN(new_n310));
  INV_X1    g124(.A(new_n307), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT32), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n308), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n306), .A2(KEYINPUT32), .A3(new_n307), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n298), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT83), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT80), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  OR3_X1    g135(.A1(new_n321), .A2(KEYINPUT16), .A3(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n318), .B1(new_n323), .B2(new_n188), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n320), .A2(KEYINPUT80), .A3(new_n322), .A4(G146), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n226), .A2(new_n319), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT81), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n226), .A2(new_n319), .A3(KEYINPUT81), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n324), .A2(new_n325), .A3(new_n330), .ZN(new_n331));
  XOR2_X1   g145(.A(KEYINPUT24), .B(G110), .Z(new_n332));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n199), .A2(G119), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n258), .A2(G128), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n258), .A2(G128), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n199), .A2(G119), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT77), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n332), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n340), .A2(KEYINPUT79), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n199), .A2(KEYINPUT23), .A3(G119), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n342), .B(new_n337), .C1(new_n335), .C2(KEYINPUT23), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(G110), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n344), .B1(new_n340), .B2(KEYINPUT79), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n331), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n336), .A2(new_n339), .A3(new_n332), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n323), .A2(new_n188), .ZN(new_n348));
  AOI21_X1  g162(.A(G146), .B1(new_n320), .B2(new_n322), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OR2_X1    g164(.A1(new_n343), .A2(KEYINPUT78), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n343), .A2(KEYINPUT78), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n352), .A2(G110), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n350), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n317), .B1(new_n346), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n351), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n356), .B(new_n347), .C1(new_n349), .C2(new_n348), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n341), .A2(new_n345), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n357), .B(KEYINPUT83), .C1(new_n358), .C2(new_n331), .ZN(new_n359));
  INV_X1    g173(.A(G953), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(G221), .A3(G234), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(KEYINPUT82), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT22), .B(G137), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n362), .B(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n355), .A2(new_n359), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n346), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n367), .A2(KEYINPUT83), .A3(new_n357), .A4(new_n364), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G234), .ZN(new_n370));
  OAI21_X1  g184(.A(G217), .B1(new_n370), .B2(G902), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n371), .B(KEYINPUT76), .ZN(new_n372));
  INV_X1    g186(.A(G902), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(KEYINPUT84), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n376), .A2(KEYINPUT85), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(KEYINPUT85), .ZN(new_n378));
  AOI21_X1  g192(.A(G902), .B1(new_n366), .B2(new_n368), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT25), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n372), .B1(new_n379), .B2(new_n380), .ZN(new_n383));
  AOI211_X1 g197(.A(new_n377), .B(new_n378), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n316), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(G475), .A2(G902), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(G113), .B(G122), .ZN(new_n388));
  INV_X1    g202(.A(G104), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT70), .B(G237), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(G214), .A3(new_n360), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n193), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n270), .A2(G143), .A3(G214), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT18), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(new_n213), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n319), .A2(new_n188), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n399), .B1(new_n328), .B2(new_n329), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n395), .A2(new_n397), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n213), .B1(new_n393), .B2(new_n394), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT98), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT17), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n406), .B1(new_n405), .B2(KEYINPUT17), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n395), .A2(G131), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT17), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n393), .A2(new_n213), .A3(new_n394), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n348), .A2(new_n349), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n390), .B(new_n404), .C1(new_n409), .C2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n390), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n319), .B(KEYINPUT19), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n226), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n324), .A3(new_n325), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n420), .B1(new_n410), .B2(new_n412), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n402), .A2(new_n398), .A3(new_n400), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n417), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n387), .B1(new_n416), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT99), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n425), .B1(new_n424), .B2(new_n426), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n424), .A2(new_n426), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G475), .ZN(new_n431));
  INV_X1    g245(.A(new_n409), .ZN(new_n432));
  INV_X1    g246(.A(new_n415), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n422), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(new_n390), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n431), .B1(new_n435), .B2(new_n373), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n260), .A2(G122), .ZN(new_n438));
  INV_X1    g252(.A(G122), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G116), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(G107), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT13), .B1(new_n199), .B2(G143), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(new_n209), .ZN(new_n444));
  XNOR2_X1  g258(.A(G128), .B(G143), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n444), .B(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G107), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n439), .A2(G116), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n438), .B1(KEYINPUT14), .B2(new_n449), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n450), .A2(KEYINPUT100), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n438), .A2(KEYINPUT14), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n452), .B1(new_n450), .B2(KEYINPUT100), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n448), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n445), .B(new_n209), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n455), .B1(G107), .B2(new_n441), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n447), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT9), .B(G234), .ZN(new_n458));
  INV_X1    g272(.A(G217), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n458), .A2(new_n459), .A3(G953), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n447), .B(new_n460), .C1(new_n454), .C2(new_n456), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(KEYINPUT101), .A3(new_n373), .ZN(new_n465));
  INV_X1    g279(.A(G478), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(KEYINPUT15), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n467), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n437), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(G214), .B1(G237), .B2(G902), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT94), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT3), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n448), .A3(G104), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT87), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n478), .A2(new_n475), .A3(new_n448), .A4(G104), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G101), .ZN(new_n481));
  OAI211_X1 g295(.A(KEYINPUT86), .B(KEYINPUT3), .C1(new_n389), .C2(G107), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n448), .A2(G104), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT3), .B1(new_n389), .B2(G107), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT86), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n480), .A2(new_n481), .A3(new_n482), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n484), .A2(new_n485), .ZN(new_n489));
  INV_X1    g303(.A(new_n483), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n489), .A2(new_n482), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n481), .B1(new_n491), .B2(new_n480), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n486), .A2(new_n482), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n477), .A2(new_n479), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n494), .B(G101), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n263), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n261), .A2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g314(.A(G113), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT5), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n501), .B1(new_n259), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n261), .A2(new_n262), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n389), .A2(G107), .ZN(new_n507));
  OAI21_X1  g321(.A(G101), .B1(new_n507), .B2(new_n483), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n487), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n499), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(G110), .B(G122), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT95), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n487), .A2(KEYINPUT96), .A3(new_n508), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n515), .A2(new_n506), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT8), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n514), .B(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n506), .B2(new_n515), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n511), .A2(new_n514), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n243), .A2(new_n321), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n228), .A2(new_n231), .A3(new_n321), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n360), .A2(G224), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT7), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n522), .A2(KEYINPUT97), .A3(new_n523), .A4(new_n527), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n523), .B(new_n527), .C1(new_n321), .C2(new_n243), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT97), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n523), .ZN(new_n532));
  OAI22_X1  g346(.A1(new_n532), .A2(new_n521), .B1(new_n526), .B2(new_n525), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n528), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(G902), .B1(new_n520), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n509), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(new_n505), .A3(new_n504), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n493), .B2(new_n498), .ZN(new_n538));
  INV_X1    g352(.A(new_n514), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n537), .B(new_n514), .C1(new_n493), .C2(new_n498), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(KEYINPUT6), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n532), .A2(new_n521), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(new_n524), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT6), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n538), .A2(new_n545), .A3(new_n539), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n542), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n535), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(G210), .B1(G237), .B2(G902), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n535), .A2(new_n547), .A3(new_n549), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n474), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n360), .A2(G952), .ZN(new_n554));
  NAND2_X1  g368(.A1(G234), .A2(G237), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G898), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n360), .B1(KEYINPUT21), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(KEYINPUT21), .B2(new_n557), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n555), .A2(G902), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n556), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n553), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n472), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT89), .ZN(new_n564));
  XNOR2_X1  g378(.A(G110), .B(G140), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n360), .A2(G227), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n246), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n509), .A2(new_n228), .A3(new_n231), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G128), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n204), .A2(new_n206), .A3(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n487), .B(new_n508), .C1(new_n573), .C2(new_n207), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n569), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT12), .B1(new_n246), .B2(KEYINPUT88), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n575), .B(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT10), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n536), .A2(KEYINPUT10), .A3(new_n232), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n243), .B(new_n497), .C1(new_n488), .C2(new_n492), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n580), .A2(new_n581), .A3(new_n582), .A4(new_n569), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n568), .B1(new_n578), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n246), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(new_n583), .A3(new_n568), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n564), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n570), .A2(new_n574), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n577), .B1(new_n590), .B2(new_n246), .ZN(new_n591));
  AOI211_X1 g405(.A(new_n569), .B(new_n576), .C1(new_n570), .C2(new_n574), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n583), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n567), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(KEYINPUT89), .A3(new_n587), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n589), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G469), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT90), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n594), .A2(KEYINPUT89), .A3(new_n587), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT89), .B1(new_n594), .B2(new_n587), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n373), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT90), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n602), .A3(G469), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n583), .A2(new_n568), .ZN(new_n604));
  OR2_X1    g418(.A1(new_n604), .A2(KEYINPUT91), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(KEYINPUT91), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n578), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n568), .B1(new_n586), .B2(new_n583), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT92), .ZN(new_n609));
  OR2_X1    g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n597), .A3(new_n373), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n598), .A2(new_n603), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT93), .ZN(new_n615));
  OAI21_X1  g429(.A(G221), .B1(new_n458), .B2(G902), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n615), .B1(new_n614), .B2(new_n616), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n385), .B(new_n563), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  AND2_X1   g434(.A1(new_n308), .A2(new_n312), .ZN(new_n621));
  OAI21_X1  g435(.A(G472), .B1(new_n310), .B2(G902), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n624), .B(new_n384), .C1(new_n617), .C2(new_n618), .ZN(new_n625));
  INV_X1    g439(.A(new_n428), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n627));
  INV_X1    g441(.A(new_n429), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n434), .A2(new_n390), .ZN(new_n630));
  INV_X1    g444(.A(new_n416), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n373), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(G475), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT33), .B1(new_n460), .B2(KEYINPUT102), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n464), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n635), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n462), .A2(new_n463), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n466), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  AOI211_X1 g453(.A(G478), .B(G902), .C1(new_n462), .C2(new_n463), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n466), .A2(new_n373), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n634), .A2(new_n642), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n643), .A2(new_n562), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n625), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT34), .B(G104), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  INV_X1    g461(.A(new_n553), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n424), .B(new_n426), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n633), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n561), .B(KEYINPUT103), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n470), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n653));
  OR3_X1    g467(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n653), .B1(new_n652), .B2(new_n650), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n625), .A2(new_n648), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT105), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G107), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  NAND2_X1  g474(.A1(new_n367), .A2(new_n357), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n364), .A2(KEYINPUT36), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n375), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n369), .A2(new_n380), .A3(new_n373), .ZN(new_n665));
  INV_X1    g479(.A(new_n372), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n664), .B1(new_n667), .B2(new_n381), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n472), .A2(new_n562), .A3(new_n669), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n670), .B(new_n624), .C1(new_n617), .C2(new_n618), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT37), .B(G110), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G12));
  NAND2_X1  g487(.A1(new_n553), .A2(new_n668), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n556), .B(KEYINPUT107), .Z(new_n675));
  NOR3_X1   g489(.A1(new_n560), .A2(G900), .A3(new_n360), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT106), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n470), .A2(new_n633), .A3(new_n649), .A4(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n316), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n681), .B1(new_n617), .B2(new_n618), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  XNOR2_X1  g497(.A(KEYINPUT109), .B(KEYINPUT39), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n678), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n603), .A2(new_n613), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n602), .B1(new_n601), .B2(G469), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n616), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT93), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n685), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT40), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n471), .A2(new_n474), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n693), .A2(new_n634), .A3(new_n669), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n291), .A2(new_n275), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n695), .A2(new_n300), .ZN(new_n696));
  OAI21_X1  g510(.A(G472), .B1(new_n696), .B2(G902), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n314), .A2(new_n315), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n551), .A2(new_n552), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT38), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n694), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT108), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n692), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G143), .ZN(G45));
  OAI211_X1 g518(.A(new_n642), .B(new_n678), .C1(new_n430), .C2(new_n436), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n674), .A2(new_n705), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n316), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n617), .B2(new_n618), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  INV_X1    g523(.A(new_n644), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n612), .A2(new_n373), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G469), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n616), .A3(new_n613), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n385), .A2(new_n710), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT41), .B(G113), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  NAND4_X1  g531(.A1(new_n712), .A2(new_n553), .A3(new_n616), .A4(new_n613), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n385), .A2(new_n655), .A3(new_n654), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  NAND2_X1  g535(.A1(new_n668), .A2(new_n561), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n718), .A2(new_n472), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n316), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  OAI21_X1  g539(.A(new_n304), .B1(new_n299), .B2(new_n292), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n307), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n622), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n384), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n377), .A2(new_n378), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(new_n381), .B2(new_n667), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(KEYINPUT110), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n728), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n693), .A2(new_n699), .A3(new_n634), .ZN(new_n735));
  INV_X1    g549(.A(new_n651), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n735), .A2(new_n713), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  NOR4_X1   g553(.A1(new_n718), .A2(new_n669), .A3(new_n705), .A4(new_n728), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n321), .ZN(G27));
  INV_X1    g555(.A(KEYINPUT42), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n597), .A2(new_n373), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n584), .A2(new_n588), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n743), .B1(new_n744), .B2(G469), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n613), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n474), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n616), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n699), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n316), .A3(new_n384), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n742), .B1(new_n752), .B2(new_n705), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n313), .B1(new_n310), .B2(new_n311), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n315), .A2(new_n754), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n730), .A2(new_n733), .B1(new_n755), .B2(new_n298), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n750), .A2(new_n742), .A3(new_n705), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(KEYINPUT111), .B(G131), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(G33));
  INV_X1    g575(.A(new_n679), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n751), .A2(new_n316), .A3(new_n384), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  NOR2_X1   g578(.A1(new_n634), .A2(KEYINPUT112), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(KEYINPUT43), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n437), .A2(new_n642), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n437), .B(new_n642), .C1(new_n765), .C2(KEYINPUT43), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT113), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n768), .A2(new_n772), .A3(new_n769), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n624), .A2(new_n669), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT44), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n771), .A2(new_n774), .A3(KEYINPUT44), .A4(new_n773), .ZN(new_n778));
  INV_X1    g592(.A(new_n685), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT46), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT45), .B1(new_n589), .B2(new_n595), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n584), .A2(new_n588), .A3(new_n782), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n781), .A2(new_n597), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n780), .B1(new_n784), .B2(new_n743), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n613), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n784), .A2(new_n780), .A3(new_n743), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n616), .B(new_n779), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n788), .A2(new_n474), .A3(new_n699), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n777), .A2(new_n778), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(KEYINPUT114), .B(G137), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(G39));
  OAI21_X1  g606(.A(new_n616), .B1(new_n786), .B2(new_n787), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(KEYINPUT47), .B(new_n616), .C1(new_n786), .C2(new_n787), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n798));
  INV_X1    g612(.A(new_n705), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n699), .A2(new_n474), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n732), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n316), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n797), .A2(new_n798), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n798), .B1(new_n797), .B2(new_n802), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(G140), .Z(G42));
  NAND2_X1  g620(.A1(new_n712), .A2(new_n613), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n749), .ZN(new_n809));
  AOI211_X1 g623(.A(new_n675), .B(new_n809), .C1(new_n769), .C2(new_n768), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n728), .A2(new_n669), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OR4_X1    g626(.A1(new_n732), .A2(new_n809), .A3(new_n556), .A4(new_n698), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n813), .A2(new_n634), .A3(new_n642), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n714), .A2(new_n474), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n700), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n816), .B2(new_n815), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n675), .B1(new_n768), .B2(new_n769), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n734), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n812), .B(new_n814), .C1(KEYINPUT50), .C2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n818), .A2(KEYINPUT50), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n795), .B(new_n796), .C1(new_n616), .C2(new_n807), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n823), .B1(new_n824), .B2(new_n800), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n822), .B1(new_n820), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n822), .B(KEYINPUT51), .C1(new_n820), .C2(new_n825), .ZN(new_n829));
  OAI221_X1 g643(.A(new_n554), .B1(new_n820), .B2(new_n718), .C1(new_n813), .C2(new_n643), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n831), .A2(KEYINPUT120), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n810), .A2(new_n756), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n833), .B(KEYINPUT48), .Z(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(KEYINPUT120), .B2(new_n831), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n828), .A2(new_n829), .A3(new_n832), .A4(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n437), .A2(new_n642), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n471), .B2(new_n437), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n651), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n625), .A2(new_n648), .A3(new_n839), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n734), .A2(new_n737), .B1(new_n723), .B2(new_n316), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n715), .A3(new_n720), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n619), .A2(new_n671), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n759), .ZN(new_n845));
  INV_X1    g659(.A(new_n678), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n650), .A2(new_n846), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n471), .A2(new_n800), .A3(new_n847), .A4(new_n668), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n316), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(new_n690), .B2(new_n689), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n751), .A2(new_n799), .A3(new_n811), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n763), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT116), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n316), .B(new_n848), .C1(new_n617), .C2(new_n618), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT116), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n854), .A2(new_n855), .A3(new_n763), .A4(new_n851), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n845), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n844), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  INV_X1    g673(.A(new_n740), .ZN(new_n860));
  INV_X1    g674(.A(new_n735), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n669), .A2(new_n616), .A3(new_n678), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(new_n698), .A3(new_n862), .A4(new_n746), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n682), .A2(new_n708), .A3(new_n860), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT117), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n689), .A2(new_n690), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n740), .B1(new_n866), .B2(new_n681), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n868), .A3(new_n708), .A4(new_n863), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n864), .A2(KEYINPUT52), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n858), .A2(new_n859), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n865), .A2(new_n869), .A3(KEYINPUT52), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n844), .A3(new_n857), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT52), .B1(new_n865), .B2(new_n869), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT53), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n874), .A2(new_n878), .A3(KEYINPUT54), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n859), .B1(new_n876), .B2(new_n877), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n842), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n841), .A2(KEYINPUT118), .A3(new_n720), .A4(new_n715), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n623), .B1(new_n689), .B2(new_n690), .ZN(new_n885));
  INV_X1    g699(.A(new_n839), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n885), .A2(new_n886), .A3(new_n384), .A4(new_n553), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(KEYINPUT53), .A3(new_n619), .A4(new_n671), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n889), .A2(new_n872), .A3(new_n857), .A4(new_n873), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n880), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n879), .B1(new_n891), .B2(KEYINPUT54), .ZN(new_n892));
  OAI22_X1  g706(.A1(new_n836), .A2(new_n892), .B1(G952), .B2(G953), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n767), .B1(new_n730), .B2(new_n733), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n807), .B(KEYINPUT49), .Z(new_n895));
  NOR2_X1   g709(.A1(new_n700), .A2(new_n748), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n893), .B1(new_n698), .B2(new_n897), .ZN(G75));
  NOR2_X1   g712(.A1(new_n360), .A2(G952), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n373), .B1(new_n880), .B2(new_n890), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT56), .B1(new_n901), .B2(G210), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n542), .A2(new_n546), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n544), .ZN(new_n904));
  XNOR2_X1  g718(.A(KEYINPUT121), .B(KEYINPUT55), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n904), .B(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n900), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n901), .B2(G210), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n910), .A2(KEYINPUT122), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(KEYINPUT122), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n907), .B1(new_n911), .B2(new_n912), .ZN(G51));
  XNOR2_X1  g727(.A(new_n743), .B(KEYINPUT57), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n891), .A2(KEYINPUT54), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n880), .B2(new_n890), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n914), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n612), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n901), .A2(new_n784), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n899), .B1(new_n919), .B2(new_n920), .ZN(G54));
  NAND2_X1  g735(.A1(new_n416), .A2(new_n423), .ZN(new_n922));
  AND2_X1   g736(.A1(KEYINPUT58), .A2(G475), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n901), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n922), .B1(new_n901), .B2(new_n923), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n899), .ZN(G60));
  AND2_X1   g740(.A1(new_n636), .A2(new_n638), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n641), .B(KEYINPUT59), .Z(new_n928));
  OAI211_X1 g742(.A(new_n927), .B(new_n928), .C1(new_n915), .C2(new_n917), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n900), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n927), .B1(new_n892), .B2(new_n928), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(G63));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n933));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT60), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n880), .B2(new_n890), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n663), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n900), .B1(new_n936), .B2(new_n369), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n933), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n936), .A2(new_n369), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n941), .A2(KEYINPUT61), .A3(new_n900), .A4(new_n937), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(G66));
  OAI21_X1  g757(.A(new_n559), .B1(G224), .B2(new_n360), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT123), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n844), .B2(G953), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n903), .B1(G898), .B2(new_n360), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(G69));
  NAND2_X1  g762(.A1(new_n248), .A2(new_n257), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(new_n418), .Z(new_n950));
  NAND2_X1  g764(.A1(new_n756), .A2(new_n861), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n763), .B1(new_n951), .B2(new_n788), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n845), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n790), .B(new_n953), .C1(new_n803), .C2(new_n804), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n682), .A2(new_n708), .A3(new_n860), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT124), .ZN(new_n957));
  AOI21_X1  g771(.A(G953), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n360), .A2(G900), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n950), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n957), .A2(new_n703), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT62), .ZN(new_n962));
  INV_X1    g776(.A(new_n790), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n805), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n957), .A2(new_n965), .A3(new_n703), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n691), .A2(new_n385), .A3(new_n800), .A4(new_n838), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n962), .A2(new_n964), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n968), .A2(new_n360), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n960), .B1(new_n969), .B2(new_n950), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n360), .B1(G227), .B2(G900), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n971), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n960), .B(new_n973), .C1(new_n969), .C2(new_n950), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(G72));
  XNOR2_X1  g789(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n976));
  NAND2_X1  g790(.A1(G472), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n276), .B2(new_n300), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n874), .A2(new_n878), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n955), .A2(new_n844), .A3(new_n957), .ZN(new_n981));
  INV_X1    g795(.A(new_n978), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n267), .B(KEYINPUT126), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n984), .A2(new_n299), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n900), .B(new_n980), .C1(new_n983), .C2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n844), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n982), .B1(new_n968), .B2(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n984), .A2(new_n299), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n988), .A2(KEYINPUT127), .A3(new_n989), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n986), .B1(new_n992), .B2(new_n993), .ZN(G57));
endmodule


