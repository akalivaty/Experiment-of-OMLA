//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n802, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  AND2_X1   g001(.A1(G211gat), .A2(G218gat), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(KEYINPUT22), .B2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G211gat), .B(G218gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n205), .B(new_n202), .C1(KEYINPUT22), .C2(new_n203), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT66), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT24), .ZN(new_n213));
  INV_X1    g012(.A(G183gat), .ZN(new_n214));
  INV_X1    g013(.A(G190gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT24), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n211), .A2(KEYINPUT66), .A3(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n213), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT67), .ZN(new_n220));
  NOR2_X1   g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT64), .B1(new_n221), .B2(KEYINPUT23), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n223), .B(new_n224), .C1(G169gat), .C2(G176gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  AND3_X1   g025(.A1(new_n222), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n212), .A2(KEYINPUT24), .B1(new_n214), .B2(new_n215), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(new_n229), .A3(new_n218), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n231));
  INV_X1    g030(.A(G169gat), .ZN(new_n232));
  INV_X1    g031(.A(G176gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n224), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n220), .A2(new_n227), .A3(new_n230), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n211), .A2(new_n217), .ZN(new_n240));
  NAND3_X1  g039(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n216), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n221), .A2(KEYINPUT23), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n222), .A2(new_n225), .A3(new_n226), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n237), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n239), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G226gat), .A2(G233gat), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT26), .B1(new_n234), .B2(new_n235), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT26), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n221), .B1(new_n250), .B2(new_n226), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n211), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT69), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n254), .B(new_n211), .C1(new_n249), .C2(new_n251), .ZN(new_n255));
  AND2_X1   g054(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n215), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n258), .A2(KEYINPUT68), .A3(KEYINPUT28), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT27), .B(G183gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n261));
  OR2_X1    g060(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n260), .A2(new_n215), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n253), .A2(new_n255), .A3(new_n264), .ZN(new_n265));
  AND3_X1   g064(.A1(new_n247), .A2(new_n248), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n267), .B1(new_n247), .B2(new_n265), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n210), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n267), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n242), .A2(new_n243), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT25), .B1(new_n271), .B2(new_n227), .ZN(new_n272));
  AND4_X1   g071(.A1(new_n229), .A2(new_n213), .A3(new_n216), .A4(new_n218), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n229), .B1(new_n228), .B2(new_n218), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NOR3_X1   g074(.A1(new_n245), .A2(new_n236), .A3(new_n237), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n272), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n253), .A2(new_n255), .A3(new_n264), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n270), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n247), .A2(new_n248), .A3(new_n265), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(new_n209), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT76), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n269), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT76), .A4(new_n209), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(KEYINPUT37), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G8gat), .B(G36gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(G64gat), .B(G92gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT89), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT89), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n285), .A2(new_n291), .A3(new_n288), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n283), .A2(new_n284), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT37), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT87), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT87), .ZN(new_n296));
  AOI211_X1 g095(.A(new_n296), .B(KEYINPUT37), .C1(new_n283), .C2(new_n284), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n290), .B(new_n292), .C1(new_n295), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT38), .ZN(new_n299));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G155gat), .B(G162gat), .Z(new_n302));
  XNOR2_X1  g101(.A(G141gat), .B(G148gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(KEYINPUT2), .B2(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(G141gat), .B(G148gat), .Z(new_n305));
  XNOR2_X1  g104(.A(G155gat), .B(G162gat), .ZN(new_n306));
  INV_X1    g105(.A(G162gat), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT2), .B1(new_n307), .B2(KEYINPUT77), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(G127gat), .B(G134gat), .Z(new_n311));
  INV_X1    g110(.A(G120gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G113gat), .ZN(new_n313));
  INV_X1    g112(.A(G113gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G120gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n311), .B1(KEYINPUT71), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G113gat), .B(G120gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT71), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT1), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT1), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n322), .B1(new_n316), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n318), .A2(KEYINPUT70), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n311), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n321), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n310), .B1(new_n326), .B2(new_n321), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n301), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT78), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n304), .A2(new_n309), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(KEYINPUT3), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n321), .A2(new_n326), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(KEYINPUT3), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT4), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT1), .B1(new_n318), .B2(KEYINPUT70), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(KEYINPUT70), .B2(new_n318), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n340), .A2(new_n311), .B1(new_n317), .B2(new_n320), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n338), .B1(new_n341), .B2(new_n310), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n310), .A2(new_n321), .A3(new_n338), .A4(new_n326), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n337), .B(new_n300), .C1(new_n342), .C2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n346), .B(new_n301), .C1(new_n328), .C2(new_n329), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n331), .A2(new_n345), .A3(KEYINPUT5), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n327), .A2(KEYINPUT4), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT80), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n350), .A3(new_n343), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n301), .A2(KEYINPUT5), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n327), .A2(KEYINPUT80), .A3(KEYINPUT4), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n351), .A2(new_n337), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n337), .A2(new_n353), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n358), .A2(KEYINPUT81), .A3(new_n352), .A4(new_n351), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n348), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  XOR2_X1   g159(.A(G57gat), .B(G85gat), .Z(new_n361));
  XNOR2_X1  g160(.A(G1gat), .B(G29gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT6), .ZN(new_n367));
  INV_X1    g166(.A(new_n365), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n348), .A2(new_n356), .A3(new_n359), .A4(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n366), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n360), .A2(KEYINPUT6), .A3(new_n365), .ZN(new_n371));
  INV_X1    g170(.A(new_n288), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n293), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT88), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n295), .A2(new_n297), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n269), .A2(new_n281), .A3(KEYINPUT86), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n378), .B(KEYINPUT37), .C1(KEYINPUT86), .C2(new_n269), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT38), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(new_n380), .A3(new_n288), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n376), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n379), .A2(new_n380), .A3(new_n288), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n383), .B(KEYINPUT88), .C1(new_n295), .C2(new_n297), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n299), .A2(new_n375), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  AND2_X1   g184(.A1(G228gat), .A2(G233gat), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT29), .B1(new_n207), .B2(new_n208), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n332), .B1(new_n387), .B2(KEYINPUT3), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n386), .B1(new_n388), .B2(KEYINPUT82), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n210), .B1(new_n333), .B2(KEYINPUT29), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n388), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n390), .B(new_n388), .C1(KEYINPUT82), .C2(new_n386), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT83), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n392), .A2(KEYINPUT83), .A3(new_n393), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n397), .A2(G22gat), .ZN(new_n398));
  XOR2_X1   g197(.A(G78gat), .B(G106gat), .Z(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT31), .B(G50gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n397), .A2(G22gat), .ZN(new_n402));
  AND4_X1   g201(.A1(new_n396), .A2(new_n398), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n398), .A2(new_n402), .B1(new_n396), .B2(new_n401), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n349), .A2(new_n350), .A3(new_n343), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n301), .B1(new_n407), .B2(new_n357), .ZN(new_n408));
  OR3_X1    g207(.A1(new_n328), .A2(new_n329), .A3(new_n301), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(KEYINPUT39), .A3(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT84), .B(KEYINPUT39), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n301), .B(new_n411), .C1(new_n407), .C2(new_n357), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n368), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT85), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT40), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT40), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n413), .A2(KEYINPUT85), .A3(new_n416), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n415), .A2(new_n366), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n283), .A2(new_n284), .A3(new_n288), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n373), .A2(KEYINPUT30), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT30), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n293), .A2(new_n421), .A3(new_n372), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n406), .B1(new_n418), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n385), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n370), .A2(new_n371), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n405), .B1(new_n427), .B2(new_n423), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT36), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n247), .A2(new_n341), .A3(new_n265), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT72), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n335), .B1(new_n277), .B2(new_n278), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n247), .A2(KEYINPUT72), .A3(new_n341), .A4(new_n265), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g234(.A1(G227gat), .A2(G233gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G71gat), .B(G99gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(G43gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT74), .B(G15gat), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n439), .B(new_n440), .Z(new_n441));
  NAND4_X1  g240(.A1(new_n437), .A2(KEYINPUT32), .A3(KEYINPUT33), .A4(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT73), .ZN(new_n443));
  INV_X1    g242(.A(new_n441), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT33), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n437), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n442), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT75), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(new_n435), .B2(new_n436), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(KEYINPUT34), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT32), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n435), .B2(new_n436), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n452), .B1(new_n446), .B2(KEYINPUT73), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n447), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT34), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n449), .B(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n446), .A2(KEYINPUT73), .ZN(new_n457));
  INV_X1    g256(.A(new_n452), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n437), .A2(new_n445), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n460), .A2(new_n443), .A3(new_n441), .ZN(new_n461));
  INV_X1    g260(.A(new_n442), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n456), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n429), .B1(new_n454), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n459), .A2(new_n463), .A3(new_n456), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n450), .B1(new_n447), .B2(new_n453), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n467), .A3(KEYINPUT36), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n428), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n466), .A2(new_n467), .A3(new_n405), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n427), .A2(new_n423), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT35), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n466), .A2(new_n467), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n427), .A2(new_n423), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT35), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n473), .A2(new_n474), .A3(new_n475), .A4(new_n405), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n426), .A2(new_n469), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(G50gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(G43gat), .ZN(new_n479));
  INV_X1    g278(.A(G43gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(G50gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT92), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT92), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(KEYINPUT15), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT14), .ZN(new_n487));
  INV_X1    g286(.A(G29gat), .ZN(new_n488));
  INV_X1    g287(.A(G36gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n490), .A2(new_n491), .B1(G29gat), .B2(G36gat), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(KEYINPUT95), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT95), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n495), .A2(new_n487), .A3(new_n488), .A4(new_n489), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n496), .A3(new_n491), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT96), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(G29gat), .A2(G36gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT97), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT93), .B(KEYINPUT15), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n481), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n480), .A2(KEYINPUT94), .A3(G50gat), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n504), .A2(new_n479), .A3(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n486), .B(new_n501), .C1(new_n502), .C2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n493), .B1(new_n499), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT17), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G15gat), .B(G22gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT16), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(G1gat), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(G1gat), .B2(new_n511), .ZN(new_n514));
  XOR2_X1   g313(.A(new_n514), .B(G8gat), .Z(new_n515));
  OAI211_X1 g314(.A(new_n493), .B(KEYINPUT17), .C1(new_n499), .C2(new_n507), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n510), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n515), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n508), .ZN(new_n519));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT18), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n515), .B(new_n508), .Z(new_n524));
  XOR2_X1   g323(.A(new_n520), .B(KEYINPUT13), .Z(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n517), .A2(KEYINPUT18), .A3(new_n519), .A4(new_n520), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n523), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(G169gat), .B(G197gat), .Z(new_n529));
  XNOR2_X1  g328(.A(G113gat), .B(G141gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(KEYINPUT90), .B(KEYINPUT11), .Z(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT91), .B(KEYINPUT12), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n535), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n523), .A2(new_n526), .A3(new_n537), .A4(new_n527), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(KEYINPUT98), .A2(G57gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(G64gat), .ZN(new_n542));
  INV_X1    g341(.A(G71gat), .ZN(new_n543));
  INV_X1    g342(.A(G78gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT9), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OR2_X1    g346(.A1(G57gat), .A2(G64gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(G57gat), .A2(G64gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(KEYINPUT9), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n545), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n543), .A2(new_n544), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT21), .ZN(new_n555));
  XOR2_X1   g354(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n515), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n515), .B2(new_n555), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n561), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n563), .B1(new_n558), .B2(new_n559), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n554), .A2(KEYINPUT21), .ZN(new_n566));
  XOR2_X1   g365(.A(G183gat), .B(G211gat), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n568), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n562), .A2(new_n564), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G127gat), .B(G155gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n573), .B(new_n574), .Z(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n569), .A2(new_n575), .A3(new_n571), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(G85gat), .ZN(new_n580));
  INV_X1    g379(.A(G92gat), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT101), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT101), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n583), .A2(G85gat), .A3(G92gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(new_n584), .A3(KEYINPUT7), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(KEYINPUT8), .A2(new_n586), .B1(new_n580), .B2(new_n581), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT7), .ZN(new_n588));
  OAI211_X1 g387(.A(KEYINPUT101), .B(new_n588), .C1(new_n580), .C2(new_n581), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n585), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(G99gat), .ZN(new_n591));
  INV_X1    g390(.A(G106gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n590), .A2(new_n586), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n586), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n585), .A2(new_n595), .A3(new_n587), .A4(new_n589), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n510), .A2(new_n516), .A3(new_n597), .ZN(new_n598));
  AND3_X1   g397(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n597), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(new_n508), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G190gat), .B(G218gat), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT102), .ZN(new_n604));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n605), .B(new_n606), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n602), .A2(new_n604), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n608), .B1(new_n602), .B2(new_n604), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n603), .A2(KEYINPUT102), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  OR3_X1    g411(.A1(new_n609), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n612), .B1(new_n609), .B2(new_n610), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT103), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n590), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n554), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n597), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT10), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n554), .A2(new_n596), .A3(new_n594), .A4(new_n618), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n600), .A2(KEYINPUT10), .A3(new_n554), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT104), .ZN(new_n626));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(KEYINPUT105), .Z(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT104), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n623), .A2(new_n630), .A3(new_n624), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n620), .A2(new_n622), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n628), .ZN(new_n634));
  XNOR2_X1  g433(.A(G120gat), .B(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(G176gat), .B(G204gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n632), .A2(new_n634), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n634), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n628), .B1(new_n623), .B2(new_n624), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n637), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n579), .A2(new_n616), .A3(new_n644), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n477), .A2(new_n540), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n427), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g448(.A(KEYINPUT16), .B(G8gat), .Z(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(new_n424), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT42), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n646), .A2(new_n424), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(G8gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(G1325gat));
  AOI21_X1  g454(.A(G15gat), .B1(new_n646), .B2(new_n473), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n465), .A2(new_n468), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n646), .A2(G15gat), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(G1326gat));
  NAND2_X1  g459(.A1(new_n646), .A2(new_n406), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT106), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT43), .B(G22gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  NOR2_X1   g463(.A1(new_n477), .A2(new_n616), .ZN(new_n665));
  INV_X1    g464(.A(new_n579), .ZN(new_n666));
  AND4_X1   g465(.A1(new_n539), .A2(new_n665), .A3(new_n666), .A4(new_n644), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n667), .A2(new_n488), .A3(new_n647), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT45), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n536), .A2(KEYINPUT107), .A3(new_n538), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT107), .B1(new_n536), .B2(new_n538), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n672), .A2(new_n644), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n579), .B(KEYINPUT108), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n665), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n477), .A2(KEYINPUT44), .A3(new_n616), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n673), .B(new_n674), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G29gat), .B1(new_n678), .B2(new_n427), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n669), .A2(new_n679), .ZN(G1328gat));
  NAND3_X1  g479(.A1(new_n667), .A2(new_n489), .A3(new_n424), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(KEYINPUT46), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT109), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(KEYINPUT46), .ZN(new_n685));
  OAI21_X1  g484(.A(G36gat), .B1(new_n678), .B2(new_n423), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(G1329gat));
  NAND3_X1  g486(.A1(new_n667), .A2(new_n480), .A3(new_n473), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT110), .Z(new_n689));
  OAI21_X1  g488(.A(G43gat), .B1(new_n678), .B2(new_n657), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(KEYINPUT47), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n688), .B(KEYINPUT110), .ZN(new_n693));
  INV_X1    g492(.A(new_n690), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n691), .A2(new_n695), .ZN(G1330gat));
  OAI21_X1  g495(.A(G50gat), .B1(new_n678), .B2(new_n405), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n667), .A2(new_n478), .A3(new_n406), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT111), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT48), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1331gat));
  NAND3_X1  g500(.A1(new_n415), .A2(new_n366), .A3(new_n417), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n405), .B1(new_n702), .B2(new_n423), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n382), .A2(new_n384), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n374), .B1(new_n298), .B2(KEYINPUT38), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n471), .A2(new_n406), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n466), .A2(new_n467), .A3(KEYINPUT36), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT36), .B1(new_n466), .B2(new_n467), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n466), .A2(new_n467), .A3(new_n405), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n475), .B1(new_n711), .B2(new_n474), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n470), .A2(KEYINPUT35), .A3(new_n471), .ZN(new_n713));
  OAI22_X1  g512(.A1(new_n706), .A2(new_n710), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n672), .A2(new_n644), .ZN(new_n715));
  AND4_X1   g514(.A1(new_n714), .A2(new_n579), .A3(new_n616), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n647), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n424), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT49), .B(G64gat), .Z(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n719), .B2(new_n721), .ZN(G1333gat));
  NAND3_X1  g521(.A1(new_n716), .A2(G71gat), .A3(new_n658), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n716), .A2(new_n473), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n724), .B2(G71gat), .ZN(new_n725));
  XOR2_X1   g524(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1334gat));
  NAND2_X1  g526(.A1(new_n716), .A2(new_n406), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g528(.A1(new_n676), .A2(new_n677), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n666), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  OR3_X1    g532(.A1(new_n733), .A2(KEYINPUT113), .A3(new_n427), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT113), .B1(new_n733), .B2(new_n427), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(G85gat), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT114), .B1(new_n477), .B2(new_n616), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n672), .A2(new_n579), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT114), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n714), .A2(new_n739), .A3(new_n615), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n737), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n743), .A2(new_n580), .A3(new_n647), .A4(new_n643), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n736), .A2(new_n744), .ZN(G1336gat));
  AOI21_X1  g544(.A(new_n581), .B1(new_n732), .B2(new_n424), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n743), .A2(new_n581), .A3(new_n424), .A4(new_n643), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n741), .A2(KEYINPUT115), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT115), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n737), .A2(new_n740), .A3(new_n752), .A4(new_n738), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n751), .A2(new_n742), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT116), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n741), .A2(new_n742), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n751), .A2(new_n757), .A3(new_n742), .A4(new_n753), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n423), .A2(G92gat), .A3(new_n644), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n746), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n750), .B1(new_n761), .B2(new_n749), .ZN(G1337gat));
  OAI21_X1  g561(.A(G99gat), .B1(new_n733), .B2(new_n657), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n743), .A2(new_n591), .A3(new_n473), .A4(new_n643), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(G1338gat));
  AOI21_X1  g564(.A(new_n592), .B1(new_n732), .B2(new_n406), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n405), .A2(G106gat), .A3(new_n644), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT53), .B1(new_n743), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n766), .B1(new_n759), .B2(new_n768), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(G1339gat));
  NAND3_X1  g572(.A1(new_n623), .A2(new_n628), .A3(new_n624), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n632), .A2(KEYINPUT54), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT54), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n638), .B1(new_n641), .B2(new_n776), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n775), .A2(KEYINPUT55), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT55), .B1(new_n775), .B2(new_n777), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n780), .B(new_n639), .C1(new_n670), .C2(new_n671), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n524), .A2(new_n525), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n520), .B1(new_n517), .B2(new_n519), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n533), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n784), .A2(new_n538), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n643), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n615), .B1(new_n781), .B2(new_n786), .ZN(new_n787));
  AND4_X1   g586(.A1(new_n615), .A2(new_n780), .A3(new_n639), .A4(new_n785), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n674), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n645), .A2(new_n672), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n470), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n424), .A2(new_n427), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(new_n314), .A3(new_n672), .ZN(new_n796));
  OAI21_X1  g595(.A(G113gat), .B1(new_n794), .B2(new_n540), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g597(.A(new_n798), .B(KEYINPUT117), .Z(G1340gat));
  NOR2_X1   g598(.A1(new_n794), .A2(new_n644), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(new_n312), .ZN(G1341gat));
  INV_X1    g600(.A(G127gat), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n794), .A2(new_n802), .A3(new_n674), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT118), .ZN(new_n804));
  AOI21_X1  g603(.A(G127gat), .B1(new_n795), .B2(new_n579), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(G1342gat));
  NAND2_X1  g605(.A1(new_n795), .A2(new_n615), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(G134gat), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT56), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(G134gat), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(G1343gat));
  INV_X1    g610(.A(G141gat), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n789), .A2(new_n791), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n814), .A3(new_n406), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n775), .A2(new_n777), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n775), .A2(KEYINPUT55), .A3(new_n777), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(new_n639), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n786), .B1(new_n820), .B2(new_n540), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n616), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n820), .A2(new_n616), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n785), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n790), .B1(new_n825), .B2(new_n666), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT57), .B1(new_n826), .B2(new_n405), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n657), .A2(new_n793), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n815), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n812), .B1(new_n830), .B2(new_n672), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n813), .A2(new_n829), .A3(new_n812), .A4(new_n406), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(new_n540), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT58), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n815), .A2(new_n827), .A3(new_n539), .A4(new_n829), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT58), .B1(new_n835), .B2(G141gat), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT119), .B1(new_n832), .B2(new_n540), .ZN(new_n837));
  AOI211_X1 g636(.A(new_n405), .B(new_n828), .C1(new_n789), .C2(new_n791), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n838), .A2(new_n839), .A3(new_n812), .A4(new_n539), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n836), .A2(KEYINPUT120), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT120), .B1(new_n836), .B2(new_n841), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n834), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(KEYINPUT121), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n846), .B(new_n834), .C1(new_n842), .C2(new_n843), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(G1344gat));
  INV_X1    g647(.A(G148gat), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n838), .A2(new_n849), .A3(new_n643), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n405), .B1(new_n789), .B2(new_n791), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n852), .A2(new_n814), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n823), .A2(KEYINPUT122), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n823), .A2(KEYINPUT122), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n785), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n579), .B1(new_n856), .B2(new_n822), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n645), .A2(new_n539), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n814), .B(new_n406), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n643), .A3(new_n829), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n851), .B1(new_n861), .B2(G148gat), .ZN(new_n862));
  AOI211_X1 g661(.A(KEYINPUT59), .B(new_n849), .C1(new_n830), .C2(new_n643), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n850), .B1(new_n862), .B2(new_n863), .ZN(G1345gat));
  AOI21_X1  g663(.A(G155gat), .B1(new_n838), .B2(new_n579), .ZN(new_n865));
  INV_X1    g664(.A(new_n830), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n674), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n865), .B1(new_n867), .B2(G155gat), .ZN(G1346gat));
  XOR2_X1   g667(.A(KEYINPUT77), .B(G162gat), .Z(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(new_n838), .B2(new_n615), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n866), .A2(new_n616), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n869), .ZN(G1347gat));
  NOR2_X1   g671(.A1(new_n647), .A2(new_n423), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n792), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(G169gat), .B1(new_n874), .B2(new_n540), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT123), .ZN(new_n876));
  INV_X1    g675(.A(new_n874), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n232), .A3(new_n672), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(G1348gat));
  AOI22_X1  g678(.A1(new_n877), .A2(new_n643), .B1(KEYINPUT124), .B2(G176gat), .ZN(new_n880));
  NOR2_X1   g679(.A1(KEYINPUT124), .A2(G176gat), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n880), .B(new_n881), .Z(G1349gat));
  NAND3_X1  g681(.A1(new_n877), .A2(new_n260), .A3(new_n579), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n884));
  OAI21_X1  g683(.A(G183gat), .B1(new_n874), .B2(new_n674), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT60), .ZN(G1350gat));
  XNOR2_X1  g686(.A(KEYINPUT61), .B(G190gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n616), .ZN(new_n890));
  MUX2_X1   g689(.A(new_n888), .B(new_n889), .S(new_n890), .Z(G1351gat));
  NAND2_X1  g690(.A1(new_n657), .A2(new_n873), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n853), .A2(new_n859), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G197gat), .B1(new_n894), .B2(new_n540), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n852), .A2(new_n893), .ZN(new_n896));
  INV_X1    g695(.A(G197gat), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n672), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n895), .B1(new_n896), .B2(new_n898), .ZN(G1352gat));
  NAND3_X1  g698(.A1(new_n860), .A2(new_n643), .A3(new_n893), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(G204gat), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n896), .A2(G204gat), .A3(new_n644), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT62), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(G1353gat));
  NAND3_X1  g703(.A1(new_n860), .A2(new_n579), .A3(new_n893), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G211gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(KEYINPUT126), .A3(KEYINPUT63), .ZN(new_n907));
  OR3_X1    g706(.A1(new_n896), .A2(G211gat), .A3(new_n666), .ZN(new_n908));
  NAND2_X1  g707(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n909));
  OR2_X1    g708(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n905), .A2(G211gat), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n907), .A2(new_n908), .A3(new_n911), .ZN(G1354gat));
  OAI21_X1  g711(.A(G218gat), .B1(new_n894), .B2(new_n616), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n616), .A2(G218gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n896), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


