

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726;

  NOR2_X1 U369 ( .A1(n721), .A2(n723), .ZN(n365) );
  AND2_X1 U370 ( .A1(n641), .A2(n640), .ZN(n644) );
  XNOR2_X1 U371 ( .A(n377), .B(n348), .ZN(n533) );
  XNOR2_X2 U372 ( .A(n587), .B(KEYINPUT33), .ZN(n673) );
  XNOR2_X2 U373 ( .A(n550), .B(KEYINPUT38), .ZN(n659) );
  INV_X2 U374 ( .A(n527), .ZN(n550) );
  XNOR2_X2 U375 ( .A(n522), .B(n523), .ZN(n561) );
  NOR2_X1 U376 ( .A1(n683), .A2(n695), .ZN(n364) );
  NOR2_X1 U377 ( .A1(n688), .A2(n695), .ZN(n363) );
  NOR2_X1 U378 ( .A1(n367), .A2(n695), .ZN(n615) );
  OR2_X1 U379 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U380 ( .A1(n645), .A2(n644), .ZN(n585) );
  XNOR2_X2 U381 ( .A(KEYINPUT1), .B(n533), .ZN(n645) );
  INV_X1 U382 ( .A(KEYINPUT48), .ZN(n388) );
  AND2_X2 U383 ( .A1(n611), .A2(n610), .ZN(n690) );
  NOR2_X1 U384 ( .A1(n608), .A2(n411), .ZN(n410) );
  NAND2_X1 U385 ( .A1(n387), .A2(n725), .ZN(n608) );
  XNOR2_X1 U386 ( .A(n389), .B(n388), .ZN(n387) );
  AND2_X1 U387 ( .A1(n547), .A2(n349), .ZN(n390) );
  NAND2_X1 U388 ( .A1(n639), .A2(n605), .ZN(n411) );
  XNOR2_X1 U389 ( .A(n546), .B(n356), .ZN(n723) );
  NOR2_X1 U390 ( .A1(n518), .A2(n511), .ZN(n535) );
  NOR2_X1 U391 ( .A1(n657), .A2(n661), .ZN(n543) );
  AND2_X1 U392 ( .A1(n533), .A2(n644), .ZN(n576) );
  XNOR2_X1 U393 ( .A(n415), .B(n494), .ZN(n692) );
  XNOR2_X2 U394 ( .A(n376), .B(n375), .ZN(n726) );
  INV_X1 U395 ( .A(G146), .ZN(n500) );
  NAND2_X1 U396 ( .A1(n713), .A2(G224), .ZN(n407) );
  BUF_X1 U397 ( .A(n517), .Z(n651) );
  NOR2_X1 U398 ( .A1(n679), .A2(G902), .ZN(n377) );
  XNOR2_X1 U399 ( .A(n414), .B(n496), .ZN(n641) );
  OR2_X1 U400 ( .A1(n692), .A2(G902), .ZN(n414) );
  XNOR2_X1 U401 ( .A(n476), .B(G134), .ZN(n395) );
  XNOR2_X1 U402 ( .A(G131), .B(G137), .ZN(n476) );
  XNOR2_X1 U403 ( .A(n447), .B(n357), .ZN(n492) );
  INV_X1 U404 ( .A(KEYINPUT8), .ZN(n357) );
  XOR2_X1 U405 ( .A(KEYINPUT6), .B(n651), .Z(n586) );
  XNOR2_X1 U406 ( .A(n413), .B(G146), .ZN(n451) );
  INV_X1 U407 ( .A(G125), .ZN(n413) );
  XNOR2_X1 U408 ( .A(G107), .B(G104), .ZN(n479) );
  XNOR2_X1 U409 ( .A(n409), .B(n430), .ZN(n408) );
  XOR2_X1 U410 ( .A(KEYINPUT17), .B(KEYINPUT80), .Z(n430) );
  INV_X1 U411 ( .A(n451), .ZN(n409) );
  INV_X1 U412 ( .A(KEYINPUT0), .ZN(n406) );
  NAND2_X1 U413 ( .A1(n560), .A2(n406), .ZN(n404) );
  XOR2_X1 U414 ( .A(n506), .B(KEYINPUT72), .Z(n429) );
  XOR2_X1 U415 ( .A(KEYINPUT83), .B(KEYINPUT23), .Z(n490) );
  XNOR2_X1 U416 ( .A(KEYINPUT84), .B(KEYINPUT24), .ZN(n489) );
  XNOR2_X1 U417 ( .A(G128), .B(G119), .ZN(n487) );
  XOR2_X1 U418 ( .A(G137), .B(G110), .Z(n488) );
  XNOR2_X1 U419 ( .A(n451), .B(n412), .ZN(n710) );
  XNOR2_X1 U420 ( .A(G140), .B(KEYINPUT10), .ZN(n412) );
  XNOR2_X1 U421 ( .A(n382), .B(n381), .ZN(n380) );
  INV_X1 U422 ( .A(KEYINPUT104), .ZN(n381) );
  INV_X1 U423 ( .A(KEYINPUT36), .ZN(n530) );
  NOR2_X1 U424 ( .A1(n573), .A2(n567), .ZN(n568) );
  XNOR2_X1 U425 ( .A(n355), .B(KEYINPUT22), .ZN(n570) );
  NAND2_X1 U426 ( .A1(n575), .A2(n562), .ZN(n355) );
  NOR2_X1 U427 ( .A1(n651), .A2(n528), .ZN(n520) );
  XNOR2_X1 U428 ( .A(G478), .B(n450), .ZN(n540) );
  NOR2_X1 U429 ( .A1(n570), .A2(n645), .ZN(n572) );
  XNOR2_X1 U430 ( .A(n394), .B(n391), .ZN(n616) );
  XNOR2_X1 U431 ( .A(n504), .B(n392), .ZN(n391) );
  XNOR2_X1 U432 ( .A(n393), .B(n505), .ZN(n392) );
  NAND2_X1 U433 ( .A1(n690), .A2(G472), .ZN(n373) );
  INV_X1 U434 ( .A(KEYINPUT64), .ZN(n369) );
  NAND2_X1 U435 ( .A1(n690), .A2(G478), .ZN(n399) );
  INV_X1 U436 ( .A(KEYINPUT47), .ZN(n359) );
  INV_X1 U437 ( .A(KEYINPUT4), .ZN(n432) );
  XNOR2_X1 U438 ( .A(KEYINPUT69), .B(G101), .ZN(n421) );
  NOR2_X1 U439 ( .A1(G953), .A2(G237), .ZN(n501) );
  OR2_X1 U440 ( .A1(G902), .A2(G237), .ZN(n499) );
  NOR2_X1 U441 ( .A1(n641), .A2(n518), .ZN(n519) );
  XNOR2_X1 U442 ( .A(n508), .B(n507), .ZN(n517) );
  NOR2_X1 U443 ( .A1(G902), .A2(n616), .ZN(n508) );
  XNOR2_X1 U444 ( .A(n500), .B(KEYINPUT88), .ZN(n393) );
  XNOR2_X1 U445 ( .A(G116), .B(G113), .ZN(n505) );
  XNOR2_X1 U446 ( .A(n423), .B(n422), .ZN(n506) );
  XOR2_X1 U447 ( .A(KEYINPUT3), .B(G119), .Z(n422) );
  XNOR2_X1 U448 ( .A(n421), .B(n420), .ZN(n423) );
  INV_X1 U449 ( .A(KEYINPUT79), .ZN(n420) );
  INV_X1 U450 ( .A(G953), .ZN(n704) );
  XNOR2_X1 U451 ( .A(n368), .B(n603), .ZN(n705) );
  NOR2_X1 U452 ( .A1(n602), .A2(n601), .ZN(n368) );
  XNOR2_X1 U453 ( .A(n362), .B(n361), .ZN(n445) );
  XNOR2_X1 U454 ( .A(n442), .B(n444), .ZN(n362) );
  XNOR2_X1 U455 ( .A(G122), .B(G143), .ZN(n453) );
  XNOR2_X1 U456 ( .A(n482), .B(n378), .ZN(n679) );
  XNOR2_X1 U457 ( .A(n711), .B(n481), .ZN(n378) );
  XOR2_X1 U458 ( .A(G110), .B(G101), .Z(n478) );
  XNOR2_X1 U459 ( .A(n408), .B(n407), .ZN(n436) );
  XNOR2_X1 U460 ( .A(n572), .B(KEYINPUT101), .ZN(n595) );
  NAND2_X2 U461 ( .A1(n403), .A2(n400), .ZN(n575) );
  AND2_X1 U462 ( .A1(n405), .A2(n404), .ZN(n403) );
  NOR2_X1 U463 ( .A1(n560), .A2(n406), .ZN(n401) );
  XOR2_X1 U464 ( .A(n710), .B(n491), .Z(n494) );
  XNOR2_X1 U465 ( .A(n493), .B(n495), .ZN(n415) );
  XNOR2_X1 U466 ( .A(n385), .B(KEYINPUT106), .ZN(n725) );
  XNOR2_X1 U467 ( .A(n549), .B(n353), .ZN(n386) );
  INV_X1 U468 ( .A(KEYINPUT42), .ZN(n356) );
  XNOR2_X1 U469 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n538) );
  XNOR2_X1 U470 ( .A(n530), .B(KEYINPUT109), .ZN(n531) );
  XNOR2_X1 U471 ( .A(n592), .B(n591), .ZN(n722) );
  NOR2_X1 U472 ( .A1(n590), .A2(n589), .ZN(n592) );
  INV_X1 U473 ( .A(KEYINPUT32), .ZN(n375) );
  OR2_X1 U474 ( .A1(n570), .A2(n569), .ZN(n376) );
  NOR2_X1 U475 ( .A1(n596), .A2(n595), .ZN(n623) );
  XNOR2_X1 U476 ( .A(n574), .B(KEYINPUT100), .ZN(n724) );
  NOR2_X1 U477 ( .A1(n573), .A2(n566), .ZN(n360) );
  NAND2_X1 U478 ( .A1(n372), .A2(n371), .ZN(n370) );
  XNOR2_X1 U479 ( .A(n373), .B(n352), .ZN(n372) );
  XNOR2_X1 U480 ( .A(n399), .B(n398), .ZN(n397) );
  INV_X1 U481 ( .A(n689), .ZN(n398) );
  XNOR2_X1 U482 ( .A(n687), .B(n686), .ZN(n688) );
  NOR2_X1 U483 ( .A1(n608), .A2(n552), .ZN(n712) );
  XOR2_X1 U484 ( .A(KEYINPUT68), .B(G469), .Z(n348) );
  AND2_X1 U485 ( .A1(n526), .A2(n525), .ZN(n349) );
  AND2_X1 U486 ( .A1(n712), .A2(n705), .ZN(n350) );
  OR2_X1 U487 ( .A1(n595), .A2(n564), .ZN(n351) );
  XOR2_X1 U488 ( .A(n616), .B(n416), .Z(n352) );
  XNOR2_X1 U489 ( .A(KEYINPUT105), .B(KEYINPUT43), .ZN(n353) );
  XOR2_X1 U490 ( .A(n606), .B(KEYINPUT67), .Z(n354) );
  NOR2_X1 U491 ( .A1(n713), .A2(G952), .ZN(n695) );
  XNOR2_X1 U492 ( .A(n682), .B(n418), .ZN(n683) );
  XNOR2_X1 U493 ( .A(n612), .B(n613), .ZN(n367) );
  INV_X1 U494 ( .A(n695), .ZN(n371) );
  AND2_X1 U495 ( .A1(n572), .A2(n360), .ZN(n574) );
  NAND2_X1 U496 ( .A1(n492), .A2(G221), .ZN(n493) );
  NAND2_X1 U497 ( .A1(n524), .A2(n358), .ZN(n525) );
  XNOR2_X1 U498 ( .A(n628), .B(n359), .ZN(n358) );
  INV_X1 U499 ( .A(n443), .ZN(n361) );
  NAND2_X1 U500 ( .A1(n390), .A2(n638), .ZN(n389) );
  XNOR2_X1 U501 ( .A(n363), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U502 ( .A(n364), .B(KEYINPUT120), .ZN(G54) );
  XNOR2_X1 U503 ( .A(n365), .B(KEYINPUT46), .ZN(n547) );
  NAND2_X1 U504 ( .A1(n366), .A2(n354), .ZN(n611) );
  NAND2_X1 U505 ( .A1(n410), .A2(n705), .ZN(n366) );
  NAND2_X1 U506 ( .A1(n402), .A2(n401), .ZN(n400) );
  XNOR2_X1 U507 ( .A(n452), .B(n424), .ZN(n426) );
  NAND2_X1 U508 ( .A1(n713), .A2(G227), .ZN(n477) );
  XNOR2_X2 U509 ( .A(n369), .B(G953), .ZN(n713) );
  XNOR2_X1 U510 ( .A(n370), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U511 ( .A1(n351), .A2(n374), .ZN(n571) );
  NAND2_X1 U512 ( .A1(n726), .A2(KEYINPUT44), .ZN(n374) );
  NOR2_X1 U513 ( .A1(n670), .A2(n379), .ZN(n671) );
  INV_X1 U514 ( .A(n610), .ZN(n379) );
  NAND2_X1 U515 ( .A1(n609), .A2(n705), .ZN(n610) );
  NAND2_X1 U516 ( .A1(n380), .A2(n658), .ZN(n548) );
  NAND2_X1 U517 ( .A1(n383), .A2(n631), .ZN(n382) );
  XNOR2_X1 U518 ( .A(n529), .B(n384), .ZN(n383) );
  INV_X1 U519 ( .A(KEYINPUT103), .ZN(n384) );
  NAND2_X1 U520 ( .A1(n386), .A2(n550), .ZN(n385) );
  XNOR2_X1 U521 ( .A(n506), .B(n711), .ZN(n394) );
  XNOR2_X2 U522 ( .A(n475), .B(n395), .ZN(n711) );
  XNOR2_X1 U523 ( .A(n426), .B(n443), .ZN(n427) );
  NAND2_X1 U524 ( .A1(n397), .A2(n371), .ZN(n396) );
  XNOR2_X1 U525 ( .A(n396), .B(KEYINPUT121), .ZN(G63) );
  INV_X1 U526 ( .A(n561), .ZN(n402) );
  NAND2_X1 U527 ( .A1(n561), .A2(n406), .ZN(n405) );
  XNOR2_X1 U528 ( .A(KEYINPUT62), .B(KEYINPUT110), .ZN(n416) );
  XOR2_X1 U529 ( .A(n469), .B(KEYINPUT75), .Z(n417) );
  XOR2_X1 U530 ( .A(n681), .B(n680), .Z(n418) );
  XNOR2_X1 U531 ( .A(KEYINPUT76), .B(n607), .ZN(n419) );
  XNOR2_X1 U532 ( .A(n480), .B(n500), .ZN(n481) );
  NOR2_X1 U533 ( .A1(n608), .A2(n419), .ZN(n609) );
  INV_X1 U534 ( .A(KEYINPUT59), .ZN(n684) );
  XNOR2_X1 U535 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U536 ( .A(n532), .B(n531), .ZN(n534) );
  XNOR2_X1 U537 ( .A(KEYINPUT54), .B(KEYINPUT117), .ZN(n439) );
  XOR2_X2 U538 ( .A(G113), .B(G104), .Z(n452) );
  XOR2_X1 U539 ( .A(KEYINPUT16), .B(KEYINPUT71), .Z(n424) );
  XNOR2_X1 U540 ( .A(G107), .B(G122), .ZN(n425) );
  XNOR2_X1 U541 ( .A(n425), .B(G116), .ZN(n443) );
  XNOR2_X1 U542 ( .A(n427), .B(G110), .ZN(n428) );
  XNOR2_X1 U543 ( .A(n429), .B(n428), .ZN(n696) );
  XNOR2_X2 U544 ( .A(G143), .B(G128), .ZN(n442) );
  INV_X1 U545 ( .A(n442), .ZN(n431) );
  NAND2_X1 U546 ( .A1(n431), .A2(KEYINPUT4), .ZN(n434) );
  NAND2_X1 U547 ( .A1(n432), .A2(n442), .ZN(n433) );
  NAND2_X1 U548 ( .A1(n434), .A2(n433), .ZN(n475) );
  XOR2_X1 U549 ( .A(n475), .B(KEYINPUT18), .Z(n435) );
  XNOR2_X1 U550 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U551 ( .A(n696), .B(n437), .ZN(n468) );
  XNOR2_X1 U552 ( .A(n468), .B(KEYINPUT55), .ZN(n438) );
  XOR2_X1 U553 ( .A(n439), .B(n438), .Z(n613) );
  XOR2_X1 U554 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n441) );
  XNOR2_X1 U555 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n440) );
  XNOR2_X1 U556 ( .A(n441), .B(n440), .ZN(n446) );
  XOR2_X1 U557 ( .A(G134), .B(KEYINPUT95), .Z(n444) );
  XOR2_X1 U558 ( .A(n446), .B(n445), .Z(n449) );
  NAND2_X1 U559 ( .A1(n713), .A2(G234), .ZN(n447) );
  NAND2_X1 U560 ( .A1(G217), .A2(n492), .ZN(n448) );
  XNOR2_X1 U561 ( .A(n449), .B(n448), .ZN(n689) );
  NOR2_X1 U562 ( .A1(n689), .A2(G902), .ZN(n450) );
  XNOR2_X1 U563 ( .A(n453), .B(n452), .ZN(n457) );
  XOR2_X1 U564 ( .A(KEYINPUT90), .B(KEYINPUT11), .Z(n455) );
  XNOR2_X1 U565 ( .A(KEYINPUT92), .B(KEYINPUT91), .ZN(n454) );
  XNOR2_X1 U566 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U567 ( .A(n457), .B(n456), .ZN(n461) );
  XOR2_X1 U568 ( .A(G131), .B(KEYINPUT12), .Z(n459) );
  NAND2_X1 U569 ( .A1(n501), .A2(G214), .ZN(n458) );
  XNOR2_X1 U570 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U571 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U572 ( .A(n710), .B(n462), .ZN(n685) );
  NOR2_X1 U573 ( .A1(n685), .A2(G902), .ZN(n466) );
  XOR2_X1 U574 ( .A(KEYINPUT94), .B(KEYINPUT13), .Z(n464) );
  XNOR2_X1 U575 ( .A(KEYINPUT93), .B(G475), .ZN(n463) );
  XNOR2_X1 U576 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U577 ( .A(n466), .B(n465), .ZN(n513) );
  NOR2_X1 U578 ( .A1(n540), .A2(n513), .ZN(n634) );
  AND2_X1 U579 ( .A1(n540), .A2(n513), .ZN(n537) );
  NOR2_X1 U580 ( .A1(n634), .A2(n537), .ZN(n467) );
  XNOR2_X1 U581 ( .A(n467), .B(KEYINPUT98), .ZN(n656) );
  NAND2_X1 U582 ( .A1(n656), .A2(KEYINPUT47), .ZN(n515) );
  XOR2_X1 U583 ( .A(G902), .B(KEYINPUT15), .Z(n605) );
  INV_X1 U584 ( .A(n605), .ZN(n604) );
  NAND2_X1 U585 ( .A1(n468), .A2(n604), .ZN(n470) );
  AND2_X1 U586 ( .A1(G210), .A2(n499), .ZN(n469) );
  XNOR2_X2 U587 ( .A(n470), .B(n417), .ZN(n527) );
  NAND2_X1 U588 ( .A1(G237), .A2(G234), .ZN(n471) );
  XNOR2_X1 U589 ( .A(n471), .B(KEYINPUT14), .ZN(n472) );
  NAND2_X1 U590 ( .A1(G952), .A2(n472), .ZN(n669) );
  NOR2_X1 U591 ( .A1(G953), .A2(n669), .ZN(n558) );
  NAND2_X1 U592 ( .A1(G902), .A2(n472), .ZN(n556) );
  OR2_X1 U593 ( .A1(n713), .A2(n556), .ZN(n473) );
  NOR2_X1 U594 ( .A1(G900), .A2(n473), .ZN(n474) );
  NOR2_X1 U595 ( .A1(n558), .A2(n474), .ZN(n518) );
  XNOR2_X1 U596 ( .A(n478), .B(n477), .ZN(n482) );
  XNOR2_X1 U597 ( .A(n479), .B(G140), .ZN(n480) );
  XOR2_X1 U598 ( .A(KEYINPUT25), .B(KEYINPUT86), .Z(n486) );
  XOR2_X1 U599 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n484) );
  NAND2_X1 U600 ( .A1(G234), .A2(n604), .ZN(n483) );
  XNOR2_X1 U601 ( .A(n484), .B(n483), .ZN(n497) );
  NAND2_X1 U602 ( .A1(n497), .A2(G217), .ZN(n485) );
  XNOR2_X1 U603 ( .A(n486), .B(n485), .ZN(n496) );
  XOR2_X1 U604 ( .A(n488), .B(n487), .Z(n495) );
  XNOR2_X1 U605 ( .A(n490), .B(n489), .ZN(n491) );
  NAND2_X1 U606 ( .A1(G221), .A2(n497), .ZN(n498) );
  XOR2_X1 U607 ( .A(KEYINPUT21), .B(n498), .Z(n640) );
  NAND2_X1 U608 ( .A1(G214), .A2(n499), .ZN(n658) );
  XOR2_X1 U609 ( .A(KEYINPUT5), .B(KEYINPUT87), .Z(n503) );
  NAND2_X1 U610 ( .A1(n501), .A2(G210), .ZN(n502) );
  XNOR2_X1 U611 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U612 ( .A(KEYINPUT70), .B(G472), .ZN(n507) );
  INV_X1 U613 ( .A(n517), .ZN(n578) );
  NAND2_X1 U614 ( .A1(n658), .A2(n578), .ZN(n509) );
  XOR2_X1 U615 ( .A(KEYINPUT30), .B(n509), .Z(n510) );
  NAND2_X1 U616 ( .A1(n576), .A2(n510), .ZN(n511) );
  NAND2_X1 U617 ( .A1(n527), .A2(n535), .ZN(n512) );
  XNOR2_X1 U618 ( .A(KEYINPUT107), .B(n512), .ZN(n514) );
  INV_X1 U619 ( .A(n513), .ZN(n541) );
  NOR2_X1 U620 ( .A1(n541), .A2(n540), .ZN(n584) );
  NAND2_X1 U621 ( .A1(n514), .A2(n584), .ZN(n627) );
  NAND2_X1 U622 ( .A1(n515), .A2(n627), .ZN(n516) );
  XNOR2_X1 U623 ( .A(n516), .B(KEYINPUT77), .ZN(n526) );
  NAND2_X1 U624 ( .A1(n519), .A2(n640), .ZN(n528) );
  XNOR2_X1 U625 ( .A(n520), .B(KEYINPUT28), .ZN(n521) );
  NAND2_X1 U626 ( .A1(n521), .A2(n533), .ZN(n544) );
  INV_X1 U627 ( .A(KEYINPUT19), .ZN(n523) );
  NAND2_X1 U628 ( .A1(n527), .A2(n658), .ZN(n522) );
  NOR2_X1 U629 ( .A1(n544), .A2(n561), .ZN(n628) );
  NAND2_X1 U630 ( .A1(n628), .A2(n656), .ZN(n524) );
  XNOR2_X1 U631 ( .A(KEYINPUT102), .B(n537), .ZN(n631) );
  NOR2_X1 U632 ( .A1(n586), .A2(n528), .ZN(n529) );
  NOR2_X1 U633 ( .A1(n550), .A2(n548), .ZN(n532) );
  XNOR2_X1 U634 ( .A(n645), .B(KEYINPUT78), .ZN(n565) );
  NAND2_X1 U635 ( .A1(n534), .A2(n565), .ZN(n638) );
  NAND2_X1 U636 ( .A1(n535), .A2(n659), .ZN(n536) );
  XNOR2_X1 U637 ( .A(n536), .B(KEYINPUT39), .ZN(n551) );
  AND2_X1 U638 ( .A1(n551), .A2(n537), .ZN(n539) );
  XNOR2_X1 U639 ( .A(n539), .B(n538), .ZN(n721) );
  NAND2_X1 U640 ( .A1(n541), .A2(n540), .ZN(n661) );
  NAND2_X1 U641 ( .A1(n659), .A2(n658), .ZN(n657) );
  INV_X1 U642 ( .A(KEYINPUT41), .ZN(n542) );
  XNOR2_X1 U643 ( .A(n543), .B(n542), .ZN(n674) );
  INV_X1 U644 ( .A(n544), .ZN(n545) );
  NAND2_X1 U645 ( .A1(n674), .A2(n545), .ZN(n546) );
  NOR2_X1 U646 ( .A1(n548), .A2(n645), .ZN(n549) );
  NAND2_X1 U647 ( .A1(n551), .A2(n634), .ZN(n639) );
  INV_X1 U648 ( .A(n639), .ZN(n552) );
  INV_X1 U649 ( .A(n661), .ZN(n553) );
  NAND2_X1 U650 ( .A1(n553), .A2(n640), .ZN(n554) );
  XNOR2_X1 U651 ( .A(n554), .B(KEYINPUT99), .ZN(n562) );
  NOR2_X1 U652 ( .A1(n704), .A2(G898), .ZN(n555) );
  XNOR2_X1 U653 ( .A(n555), .B(KEYINPUT81), .ZN(n697) );
  NOR2_X1 U654 ( .A1(n556), .A2(n697), .ZN(n557) );
  NOR2_X1 U655 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U656 ( .A(n559), .B(KEYINPUT82), .ZN(n560) );
  INV_X1 U657 ( .A(n641), .ZN(n566) );
  NAND2_X1 U658 ( .A1(n651), .A2(n566), .ZN(n596) );
  INV_X1 U659 ( .A(KEYINPUT44), .ZN(n563) );
  OR2_X1 U660 ( .A1(n596), .A2(n563), .ZN(n564) );
  INV_X1 U661 ( .A(n586), .ZN(n573) );
  NAND2_X1 U662 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U663 ( .A(KEYINPUT74), .B(n568), .Z(n569) );
  XNOR2_X1 U664 ( .A(n571), .B(KEYINPUT66), .ZN(n602) );
  NAND2_X1 U665 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U666 ( .A1(n578), .A2(n577), .ZN(n618) );
  INV_X1 U667 ( .A(n575), .ZN(n580) );
  NOR2_X1 U668 ( .A1(n585), .A2(n651), .ZN(n579) );
  XNOR2_X1 U669 ( .A(n579), .B(KEYINPUT89), .ZN(n653) );
  NOR2_X1 U670 ( .A1(n580), .A2(n653), .ZN(n581) );
  XOR2_X1 U671 ( .A(KEYINPUT31), .B(n581), .Z(n635) );
  NOR2_X1 U672 ( .A1(n618), .A2(n635), .ZN(n582) );
  NOR2_X1 U673 ( .A1(n656), .A2(n582), .ZN(n583) );
  NOR2_X1 U674 ( .A1(n724), .A2(n583), .ZN(n594) );
  INV_X1 U675 ( .A(n584), .ZN(n590) );
  NAND2_X1 U676 ( .A1(n673), .A2(n575), .ZN(n588) );
  XNOR2_X1 U677 ( .A(KEYINPUT34), .B(n588), .ZN(n589) );
  XNOR2_X1 U678 ( .A(KEYINPUT35), .B(KEYINPUT73), .ZN(n591) );
  NAND2_X1 U679 ( .A1(n722), .A2(KEYINPUT44), .ZN(n593) );
  AND2_X1 U680 ( .A1(n594), .A2(n593), .ZN(n600) );
  NOR2_X1 U681 ( .A1(n623), .A2(n726), .ZN(n598) );
  NOR2_X1 U682 ( .A1(n722), .A2(KEYINPUT44), .ZN(n597) );
  NAND2_X1 U683 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U684 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U685 ( .A(KEYINPUT45), .B(KEYINPUT65), .ZN(n603) );
  NAND2_X1 U686 ( .A1(n605), .A2(KEYINPUT2), .ZN(n606) );
  NAND2_X1 U687 ( .A1(KEYINPUT2), .A2(n639), .ZN(n607) );
  NAND2_X1 U688 ( .A1(n690), .A2(G210), .ZN(n612) );
  XNOR2_X1 U689 ( .A(KEYINPUT56), .B(KEYINPUT118), .ZN(n614) );
  XNOR2_X1 U690 ( .A(n615), .B(n614), .ZN(G51) );
  NAND2_X1 U691 ( .A1(n631), .A2(n618), .ZN(n617) );
  XNOR2_X1 U692 ( .A(n617), .B(G104), .ZN(G6) );
  XOR2_X1 U693 ( .A(KEYINPUT111), .B(KEYINPUT27), .Z(n620) );
  NAND2_X1 U694 ( .A1(n618), .A2(n634), .ZN(n619) );
  XNOR2_X1 U695 ( .A(n620), .B(n619), .ZN(n622) );
  XOR2_X1 U696 ( .A(G107), .B(KEYINPUT26), .Z(n621) );
  XNOR2_X1 U697 ( .A(n622), .B(n621), .ZN(G9) );
  XOR2_X1 U698 ( .A(G110), .B(n623), .Z(G12) );
  XOR2_X1 U699 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n625) );
  NAND2_X1 U700 ( .A1(n628), .A2(n634), .ZN(n624) );
  XNOR2_X1 U701 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U702 ( .A(G128), .B(n626), .ZN(G30) );
  XNOR2_X1 U703 ( .A(G143), .B(n627), .ZN(G45) );
  XOR2_X1 U704 ( .A(G146), .B(KEYINPUT113), .Z(n630) );
  NAND2_X1 U705 ( .A1(n628), .A2(n631), .ZN(n629) );
  XNOR2_X1 U706 ( .A(n630), .B(n629), .ZN(G48) );
  NAND2_X1 U707 ( .A1(n631), .A2(n635), .ZN(n632) );
  XNOR2_X1 U708 ( .A(n632), .B(KEYINPUT114), .ZN(n633) );
  XNOR2_X1 U709 ( .A(G113), .B(n633), .ZN(G15) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n636), .B(G116), .ZN(G18) );
  XOR2_X1 U712 ( .A(G125), .B(KEYINPUT37), .Z(n637) );
  XNOR2_X1 U713 ( .A(n638), .B(n637), .ZN(G27) );
  XNOR2_X1 U714 ( .A(G134), .B(n639), .ZN(G36) );
  NOR2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n643) );
  XNOR2_X1 U716 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n642) );
  XNOR2_X1 U717 ( .A(n643), .B(n642), .ZN(n649) );
  XNOR2_X1 U718 ( .A(KEYINPUT116), .B(KEYINPUT50), .ZN(n647) );
  NOR2_X1 U719 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n647), .B(n646), .ZN(n648) );
  NOR2_X1 U721 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U722 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U723 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U724 ( .A(KEYINPUT51), .B(n654), .Z(n655) );
  NAND2_X1 U725 ( .A1(n674), .A2(n655), .ZN(n666) );
  NOR2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n663) );
  NOR2_X1 U727 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U728 ( .A1(n661), .A2(n660), .ZN(n662) );
  OR2_X1 U729 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U730 ( .A1(n673), .A2(n664), .ZN(n665) );
  NAND2_X1 U731 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U732 ( .A(KEYINPUT52), .B(n667), .Z(n668) );
  NOR2_X1 U733 ( .A1(n669), .A2(n668), .ZN(n672) );
  NOR2_X1 U734 ( .A1(KEYINPUT2), .A2(n350), .ZN(n670) );
  NOR2_X1 U735 ( .A1(n672), .A2(n671), .ZN(n676) );
  NAND2_X1 U736 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U737 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U738 ( .A1(n677), .A2(G953), .ZN(n678) );
  XNOR2_X1 U739 ( .A(n678), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U740 ( .A1(n690), .A2(G469), .ZN(n682) );
  XOR2_X1 U741 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n681) );
  XNOR2_X1 U742 ( .A(n679), .B(KEYINPUT119), .ZN(n680) );
  NAND2_X1 U743 ( .A1(n690), .A2(G475), .ZN(n687) );
  NAND2_X1 U744 ( .A1(n690), .A2(G217), .ZN(n691) );
  XNOR2_X1 U745 ( .A(n691), .B(KEYINPUT122), .ZN(n693) );
  XNOR2_X1 U746 ( .A(n692), .B(n693), .ZN(n694) );
  NOR2_X1 U747 ( .A1(n695), .A2(n694), .ZN(G66) );
  XNOR2_X1 U748 ( .A(n696), .B(KEYINPUT125), .ZN(n698) );
  NAND2_X1 U749 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U750 ( .A(n699), .B(KEYINPUT126), .ZN(n709) );
  XOR2_X1 U751 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n701) );
  NAND2_X1 U752 ( .A1(G224), .A2(G953), .ZN(n700) );
  XNOR2_X1 U753 ( .A(n701), .B(n700), .ZN(n702) );
  NAND2_X1 U754 ( .A1(G898), .A2(n702), .ZN(n703) );
  XNOR2_X1 U755 ( .A(n703), .B(KEYINPUT124), .ZN(n707) );
  NAND2_X1 U756 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U757 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U758 ( .A(n709), .B(n708), .Z(G69) );
  XOR2_X1 U759 ( .A(n711), .B(n710), .Z(n715) );
  XOR2_X1 U760 ( .A(n715), .B(n712), .Z(n714) );
  NAND2_X1 U761 ( .A1(n714), .A2(n713), .ZN(n719) );
  XNOR2_X1 U762 ( .A(G227), .B(n715), .ZN(n716) );
  NAND2_X1 U763 ( .A1(n716), .A2(G900), .ZN(n717) );
  NAND2_X1 U764 ( .A1(n717), .A2(G953), .ZN(n718) );
  NAND2_X1 U765 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U766 ( .A(KEYINPUT127), .B(n720), .Z(G72) );
  XOR2_X1 U767 ( .A(n721), .B(G131), .Z(G33) );
  XOR2_X1 U768 ( .A(G122), .B(n722), .Z(G24) );
  XOR2_X1 U769 ( .A(G137), .B(n723), .Z(G39) );
  XOR2_X1 U770 ( .A(n724), .B(G101), .Z(G3) );
  XNOR2_X1 U771 ( .A(G140), .B(n725), .ZN(G42) );
  XOR2_X1 U772 ( .A(n726), .B(G119), .Z(G21) );
endmodule

