//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n550, new_n551, new_n552, new_n553, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n562, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n581,
    new_n582, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n460), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(new_n460), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n469), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n462), .A2(new_n464), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n474), .A2(G137), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n461), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT67), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  OR2_X1    g057(.A1(new_n474), .A2(KEYINPUT68), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n474), .A2(KEYINPUT68), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OAI21_X1  g062(.A(KEYINPUT69), .B1(G100), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NOR3_X1   g064(.A1(KEYINPUT69), .A2(G100), .A3(G2105), .ZN(new_n490));
  NOR3_X1   g065(.A1(new_n489), .A2(new_n490), .A3(new_n461), .ZN(new_n491));
  OR2_X1    g066(.A1(new_n471), .A2(G112), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n473), .A2(new_n471), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n491), .A2(new_n492), .B1(new_n493), .B2(G124), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n497), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n462), .A2(new_n464), .A3(new_n460), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(new_n465), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT71), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n467), .A2(new_n471), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT4), .B1(new_n502), .B2(new_n497), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(new_n498), .C1(new_n499), .C2(new_n465), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n501), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n462), .A2(new_n464), .A3(G126), .ZN(new_n509));
  NAND2_X1  g084(.A1(G114), .A2(G2104), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n471), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n477), .A2(G102), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n508), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n510), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(new_n467), .B2(G126), .ZN(new_n516));
  OAI211_X1 g091(.A(KEYINPUT70), .B(new_n512), .C1(new_n516), .C2(new_n471), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n507), .A2(new_n518), .ZN(G164));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G651), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n521), .A2(KEYINPUT72), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(KEYINPUT72), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n522), .A2(new_n523), .B1(KEYINPUT6), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G543), .ZN(new_n528));
  OR3_X1    g103(.A1(new_n528), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n529));
  OAI21_X1  g104(.A(KEYINPUT5), .B1(new_n528), .B2(KEYINPUT73), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(G50), .A2(new_n527), .B1(new_n534), .B2(G88), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT74), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n532), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n524), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(G166));
  NAND2_X1  g115(.A1(new_n525), .A2(G89), .ZN(new_n541));
  NAND2_X1  g116(.A1(G63), .A2(G651), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n531), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n526), .B(KEYINPUT75), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n543), .B1(new_n544), .B2(G51), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT7), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n545), .A2(new_n547), .ZN(G286));
  INV_X1    g123(.A(G286), .ZN(G168));
  AOI22_X1  g124(.A1(new_n532), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n524), .ZN(new_n551));
  INV_X1    g126(.A(G90), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n533), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n544), .B2(G52), .ZN(G171));
  AOI22_X1  g129(.A1(new_n532), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n524), .ZN(new_n556));
  INV_X1    g131(.A(G81), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n533), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n544), .B2(G43), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT76), .Z(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G188));
  AOI22_X1  g141(.A1(new_n532), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n524), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT80), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n568), .A2(new_n569), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n534), .A2(G91), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n572), .A2(KEYINPUT79), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(KEYINPUT79), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n570), .A2(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n527), .A2(G53), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT77), .B1(new_n576), .B2(KEYINPUT78), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(KEYINPUT9), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n577), .B(KEYINPUT9), .C1(KEYINPUT77), .C2(new_n576), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(G299));
  NAND2_X1  g155(.A1(new_n544), .A2(G52), .ZN(new_n581));
  INV_X1    g156(.A(new_n553), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G301));
  XNOR2_X1  g158(.A(new_n539), .B(KEYINPUT81), .ZN(G303));
  NAND2_X1  g159(.A1(new_n527), .A2(G49), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n534), .A2(G87), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n532), .B2(G74), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G288));
  AOI22_X1  g163(.A1(G48), .A2(new_n527), .B1(new_n534), .B2(G86), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n532), .A2(KEYINPUT82), .A3(G61), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n531), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G73), .ZN(new_n594));
  OAI21_X1  g169(.A(KEYINPUT83), .B1(new_n594), .B2(new_n528), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n590), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  NOR3_X1   g171(.A1(new_n594), .A2(new_n528), .A3(KEYINPUT83), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n589), .A2(new_n598), .ZN(G305));
  AND2_X1   g174(.A1(new_n544), .A2(G47), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n532), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n601), .A2(new_n524), .B1(new_n533), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n534), .A2(G92), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT10), .Z(new_n608));
  AOI22_X1  g183(.A1(new_n532), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT84), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G651), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n544), .A2(G54), .ZN(new_n612));
  AND3_X1   g187(.A1(new_n608), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n606), .B1(new_n613), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  INV_X1    g191(.A(G299), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G297));
  OAI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G280));
  XNOR2_X1  g194(.A(KEYINPUT85), .B(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(G860), .B2(new_n620), .ZN(G148));
  NAND2_X1  g196(.A1(new_n613), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n486), .A2(G135), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n471), .A2(G111), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n461), .B1(new_n627), .B2(KEYINPUT87), .ZN(new_n628));
  OAI221_X1 g203(.A(new_n628), .B1(KEYINPUT87), .B2(new_n627), .C1(G99), .C2(G2105), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n493), .A2(G123), .ZN(new_n630));
  AND2_X1   g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT88), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2096), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n469), .A2(new_n477), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT13), .B(G2100), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n634), .A2(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(G2427), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT90), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT89), .B(G2438), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT91), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n649), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G1341), .B(G1348), .Z(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT92), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n654), .B2(new_n655), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n649), .A2(new_n653), .ZN(new_n659));
  INV_X1    g234(.A(new_n648), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n647), .B(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n661), .A2(new_n652), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n657), .B(new_n655), .C1(new_n659), .C2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n656), .B(G14), .C1(new_n658), .C2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT93), .B(KEYINPUT17), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XOR2_X1   g245(.A(G2067), .B(G2678), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT94), .ZN(new_n673));
  INV_X1    g248(.A(new_n670), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n667), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n674), .B(new_n675), .C1(new_n669), .C2(new_n671), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n674), .A2(new_n671), .A3(new_n667), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT18), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n673), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2096), .B(G2100), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n684), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n685), .A2(new_n686), .ZN(new_n690));
  AOI22_X1  g265(.A1(new_n688), .A2(KEYINPUT20), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n690), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n692), .A2(new_n684), .A3(new_n687), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n691), .B(new_n693), .C1(KEYINPUT20), .C2(new_n688), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT95), .ZN(new_n695));
  INV_X1    g270(.A(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1986), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1991), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT96), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n697), .B(new_n702), .Z(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  NAND2_X1  g279(.A1(new_n493), .A2(G119), .ZN(new_n705));
  NOR2_X1   g280(.A1(G95), .A2(G2105), .ZN(new_n706));
  OAI21_X1  g281(.A(G2104), .B1(new_n471), .B2(G107), .ZN(new_n707));
  INV_X1    g282(.A(G131), .ZN(new_n708));
  OAI221_X1 g283(.A(new_n705), .B1(new_n706), .B2(new_n707), .C1(new_n485), .C2(new_n708), .ZN(new_n709));
  MUX2_X1   g284(.A(G25), .B(new_n709), .S(G29), .Z(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT35), .B(G1991), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT97), .Z(new_n712));
  XOR2_X1   g287(.A(new_n710), .B(new_n712), .Z(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n604), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n714), .B2(G24), .ZN(new_n716));
  INV_X1    g291(.A(G1986), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n713), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(G22), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G166), .B2(new_n714), .ZN(new_n720));
  INV_X1    g295(.A(G1971), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT98), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G16), .B2(G23), .ZN(new_n724));
  OR3_X1    g299(.A1(new_n723), .A2(G16), .A3(G23), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n724), .B(new_n725), .C1(G288), .C2(new_n714), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT33), .B(G1976), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n714), .A2(G6), .ZN(new_n729));
  INV_X1    g304(.A(G305), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(new_n714), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT32), .B(G1981), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n722), .A2(new_n728), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n718), .B1(new_n734), .B2(KEYINPUT34), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n716), .A2(new_n717), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n735), .B(new_n736), .C1(KEYINPUT34), .C2(new_n734), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT36), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n559), .A2(new_n714), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n714), .B2(G19), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(G1341), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT31), .B(G11), .Z(new_n743));
  AND2_X1   g318(.A1(KEYINPUT24), .A2(G34), .ZN(new_n744));
  NOR2_X1   g319(.A1(KEYINPUT24), .A2(G34), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n744), .A2(new_n745), .A3(G29), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n481), .B2(G29), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(G2084), .Z(new_n748));
  INV_X1    g323(.A(G29), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G27), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G164), .B2(new_n749), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G2078), .ZN(new_n752));
  OR2_X1    g327(.A1(G29), .A2(G32), .ZN(new_n753));
  NAND3_X1  g328(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT26), .Z(new_n755));
  AOI22_X1  g330(.A1(new_n493), .A2(G129), .B1(G105), .B2(new_n477), .ZN(new_n756));
  INV_X1    g331(.A(G141), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n755), .B(new_n756), .C1(new_n485), .C2(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n753), .B1(new_n758), .B2(new_n749), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT27), .B(G1996), .Z(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n759), .A2(new_n761), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n626), .A2(G29), .A3(new_n631), .ZN(new_n764));
  INV_X1    g339(.A(G28), .ZN(new_n765));
  AOI21_X1  g340(.A(G29), .B1(new_n765), .B2(KEYINPUT30), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(KEYINPUT30), .B2(new_n765), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n767), .ZN(new_n768));
  OR4_X1    g343(.A1(new_n743), .A2(new_n748), .A3(new_n752), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n714), .A2(G5), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G171), .B2(new_n714), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1961), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n714), .A2(G21), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G168), .B2(new_n714), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT101), .B(G1966), .Z(new_n775));
  XOR2_X1   g350(.A(new_n774), .B(new_n775), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n749), .A2(G33), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n477), .A2(G103), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT25), .Z(new_n779));
  AOI22_X1  g354(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n780));
  INV_X1    g355(.A(G139), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n779), .B1(new_n780), .B2(new_n471), .C1(new_n485), .C2(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT99), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n777), .B1(new_n783), .B2(new_n749), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT100), .B(G2072), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n784), .B(new_n785), .Z(new_n786));
  NOR4_X1   g361(.A1(new_n769), .A2(new_n772), .A3(new_n776), .A4(new_n786), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n787), .A2(KEYINPUT102), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(KEYINPUT102), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT103), .B(KEYINPUT23), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n714), .A2(G20), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G299), .B2(G16), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(G1956), .Z(new_n794));
  OR2_X1    g369(.A1(G104), .A2(G2105), .ZN(new_n795));
  INV_X1    g370(.A(G116), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n461), .B1(new_n796), .B2(G2105), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n493), .A2(G128), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G140), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n485), .B2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(new_n749), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n749), .A2(G26), .ZN(new_n803));
  OAI21_X1  g378(.A(KEYINPUT28), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(KEYINPUT28), .B2(new_n803), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G2067), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n749), .A2(G35), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G162), .B2(new_n749), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT29), .B(G2090), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n714), .A2(G4), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n613), .B2(new_n714), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n741), .A2(G1341), .B1(new_n813), .B2(G1348), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n811), .B(new_n814), .C1(G1348), .C2(new_n813), .ZN(new_n815));
  NOR4_X1   g390(.A1(new_n788), .A2(new_n789), .A3(new_n794), .A4(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n738), .A2(new_n742), .A3(new_n816), .ZN(G150));
  INV_X1    g392(.A(G150), .ZN(G311));
  NAND2_X1  g393(.A1(new_n544), .A2(G55), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n532), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(new_n524), .ZN(new_n821));
  INV_X1    g396(.A(G93), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n819), .B(new_n821), .C1(new_n822), .C2(new_n533), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT104), .B(G860), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT37), .Z(new_n826));
  NAND2_X1  g401(.A1(new_n613), .A2(G559), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT38), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n821), .B1(new_n533), .B2(new_n822), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n544), .B2(G55), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n544), .A2(G43), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(new_n558), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n823), .A2(new_n559), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT39), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n828), .B(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n826), .B1(new_n836), .B2(new_n824), .ZN(G145));
  XNOR2_X1  g412(.A(new_n758), .B(new_n800), .ZN(new_n838));
  OAI21_X1  g413(.A(KEYINPUT106), .B1(new_n511), .B2(new_n513), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT106), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n840), .B(new_n512), .C1(new_n516), .C2(new_n471), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n506), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT107), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n506), .A2(KEYINPUT107), .A3(new_n842), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n838), .B(new_n847), .ZN(new_n848));
  MUX2_X1   g423(.A(new_n783), .B(new_n782), .S(new_n848), .Z(new_n849));
  NAND2_X1  g424(.A1(new_n493), .A2(G130), .ZN(new_n850));
  NOR2_X1   g425(.A1(G106), .A2(G2105), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(new_n471), .B2(G118), .ZN(new_n852));
  INV_X1    g427(.A(G142), .ZN(new_n853));
  OAI221_X1 g428(.A(new_n850), .B1(new_n851), .B2(new_n852), .C1(new_n485), .C2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n709), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n637), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT108), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n849), .A2(new_n856), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n481), .B(KEYINPUT105), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n495), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n632), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n858), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n862), .B1(new_n859), .B2(new_n857), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n864), .A2(G37), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g442(.A1(new_n823), .A2(G868), .ZN(new_n868));
  INV_X1    g443(.A(G288), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n539), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n730), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n539), .B(G288), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(G305), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(G290), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n871), .A2(new_n873), .A3(new_n604), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT42), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n622), .B(new_n834), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n608), .A2(new_n611), .A3(new_n612), .ZN(new_n880));
  XNOR2_X1  g455(.A(G299), .B(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(G299), .A2(new_n613), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n880), .A2(new_n578), .A3(new_n575), .A4(new_n579), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT109), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT109), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n617), .A2(new_n887), .A3(new_n880), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n881), .A2(KEYINPUT41), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n882), .B1(new_n891), .B2(new_n879), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT110), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n878), .A2(new_n894), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n892), .A2(new_n893), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n868), .B1(new_n897), .B2(G868), .ZN(G295));
  AOI21_X1  g473(.A(new_n868), .B1(new_n897), .B2(G868), .ZN(G331));
  AND2_X1   g474(.A1(new_n889), .A2(new_n890), .ZN(new_n900));
  NAND2_X1  g475(.A1(G168), .A2(G301), .ZN(new_n901));
  NAND2_X1  g476(.A1(G286), .A2(G171), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n834), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT111), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n901), .A2(new_n833), .A3(new_n832), .A4(new_n902), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  OR3_X1    g482(.A1(new_n903), .A2(new_n834), .A3(new_n905), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT112), .B1(new_n900), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT112), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n891), .A2(new_n911), .A3(new_n908), .A4(new_n907), .ZN(new_n912));
  INV_X1    g487(.A(new_n881), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(new_n904), .A3(new_n906), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n910), .A2(new_n912), .A3(new_n877), .A4(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G37), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n910), .A2(new_n914), .A3(new_n912), .ZN(new_n918));
  INV_X1    g493(.A(new_n877), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT43), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n915), .A2(new_n916), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n881), .B1(new_n907), .B2(new_n908), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT113), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n885), .A2(KEYINPUT41), .A3(new_n888), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n904), .A2(new_n906), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n925), .B(new_n926), .C1(new_n913), .C2(KEYINPUT41), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n877), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n922), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT44), .B1(new_n921), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n929), .B1(new_n917), .B2(new_n920), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n922), .A2(new_n928), .A3(KEYINPUT43), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n931), .A2(new_n935), .ZN(G397));
  INV_X1    g511(.A(G1384), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT45), .B1(new_n847), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G40), .ZN(new_n939));
  NOR4_X1   g514(.A1(new_n472), .A2(new_n939), .A3(new_n475), .A4(new_n479), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(G1996), .A3(new_n758), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n943), .B(KEYINPUT114), .Z(new_n944));
  XNOR2_X1  g519(.A(new_n800), .B(G2067), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n941), .A2(G1996), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n944), .B(new_n946), .C1(new_n758), .C2(new_n948), .ZN(new_n949));
  OR3_X1    g524(.A1(new_n949), .A2(new_n712), .A3(new_n709), .ZN(new_n950));
  INV_X1    g525(.A(G2067), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n801), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n941), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n709), .B(new_n712), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n949), .B1(new_n942), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(G290), .A2(G1986), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n942), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT126), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT48), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n942), .A2(new_n758), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT125), .B1(new_n961), .B2(new_n946), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n962), .B1(new_n963), .B2(new_n948), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n961), .A2(new_n946), .A3(KEYINPUT125), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n964), .B(new_n965), .C1(new_n963), .C2(new_n948), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT47), .Z(new_n967));
  NOR3_X1   g542(.A1(new_n953), .A2(new_n960), .A3(new_n967), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n506), .A2(KEYINPUT107), .A3(new_n842), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT107), .B1(new_n506), .B2(new_n842), .ZN(new_n970));
  OAI211_X1 g545(.A(KEYINPUT45), .B(new_n937), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT115), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n847), .A2(KEYINPUT115), .A3(KEYINPUT45), .A4(new_n937), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n937), .B1(new_n507), .B2(new_n518), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n975), .A2(KEYINPUT116), .A3(new_n978), .A4(new_n940), .ZN(new_n979));
  INV_X1    g554(.A(G2078), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n973), .A2(new_n974), .A3(new_n978), .A4(new_n940), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT116), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n979), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n976), .A2(KEYINPUT50), .ZN(new_n987));
  AOI21_X1  g562(.A(G1384), .B1(new_n506), .B2(new_n842), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n989), .B1(new_n988), .B2(new_n990), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n940), .B(new_n987), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1961), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI211_X1 g570(.A(KEYINPUT45), .B(new_n937), .C1(new_n507), .C2(new_n518), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n940), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n988), .A2(KEYINPUT45), .ZN(new_n998));
  OR4_X1    g573(.A1(new_n985), .A2(new_n997), .A3(G2078), .A4(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n986), .A2(new_n995), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n775), .B1(new_n997), .B2(new_n998), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(new_n993), .B2(G2084), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1001), .B1(new_n1003), .B2(G286), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1002), .B(G168), .C1(new_n993), .C2(G2084), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(G8), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1001), .B1(new_n1005), .B2(G8), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT62), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(KEYINPUT51), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT62), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1010), .B(new_n1011), .C1(new_n1006), .C2(new_n1004), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1000), .A2(G171), .A3(new_n1009), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G8), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n979), .A2(new_n983), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n721), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n993), .A2(G2090), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AND2_X1   g593(.A1(KEYINPUT118), .A2(KEYINPUT55), .ZN(new_n1019));
  NOR2_X1   g594(.A1(KEYINPUT118), .A2(KEYINPUT55), .ZN(new_n1020));
  OAI211_X1 g595(.A(G303), .B(G8), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  AND2_X1   g596(.A1(G303), .A2(G8), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1021), .B1(new_n1022), .B2(new_n1019), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1018), .A2(new_n1023), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1003), .A2(G8), .A3(G168), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT63), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1013), .A2(new_n1024), .A3(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n940), .B1(new_n976), .B2(KEYINPUT50), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n988), .A2(new_n990), .ZN(new_n1030));
  OR3_X1    g605(.A1(new_n1029), .A2(G2090), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1014), .B1(new_n1016), .B2(new_n1031), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n1032), .A2(new_n1023), .ZN(new_n1033));
  XNOR2_X1  g608(.A(G305), .B(G1981), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1034), .B(KEYINPUT49), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n940), .A2(new_n988), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(G8), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(G8), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1038), .B1(G1976), .B2(new_n869), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1039), .B(new_n1040), .C1(G1976), .C2(new_n869), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1037), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1028), .A2(new_n1033), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1976), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1037), .A2(new_n1045), .A3(new_n869), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n730), .A2(new_n696), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1038), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1043), .B(new_n1025), .C1(new_n1018), .C2(new_n1023), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1048), .B1(new_n1049), .B2(KEYINPUT63), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1044), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT54), .B1(new_n1000), .B2(G171), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n984), .A2(new_n985), .B1(new_n994), .B2(new_n993), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n975), .A2(new_n940), .ZN(new_n1054));
  OR4_X1    g629(.A1(new_n985), .A2(new_n1054), .A3(G2078), .A4(new_n938), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1052), .B1(G171), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT124), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1053), .A2(KEYINPUT124), .A3(new_n1055), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1059), .A2(G171), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1000), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT54), .B1(new_n1062), .B2(G171), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1057), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1010), .B1(new_n1006), .B2(new_n1004), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1033), .A2(new_n1024), .A3(new_n1065), .A4(new_n1043), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1036), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT58), .B(G1341), .ZN(new_n1068));
  OAI22_X1  g643(.A1(new_n981), .A2(G1996), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n559), .ZN(new_n1070));
  AND2_X1   g645(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n571), .A2(new_n570), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n573), .A2(new_n574), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1074), .B1(new_n1077), .B2(KEYINPUT119), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1078), .B(G299), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT56), .B(G2072), .Z(new_n1080));
  NOR2_X1   g655(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n981), .A2(new_n1080), .B1(G1956), .B2(new_n1081), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1072), .A2(new_n1073), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT61), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1348), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n993), .A2(new_n1087), .B1(new_n1067), .B2(new_n951), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT60), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT123), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT60), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n1097), .B2(new_n1090), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n613), .B1(new_n1098), .B2(KEYINPUT123), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1093), .A2(new_n1094), .A3(new_n880), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1095), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1091), .A2(new_n1092), .A3(KEYINPUT60), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1083), .B(new_n1086), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1084), .A2(new_n1090), .A3(new_n1097), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1082), .B(KEYINPUT121), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1104), .A2(new_n613), .B1(new_n1079), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1066), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1051), .B1(new_n1064), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n604), .A2(new_n717), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n942), .B1(new_n956), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n955), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n968), .B1(new_n1108), .B2(new_n1111), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g687(.A1(new_n665), .A2(G319), .A3(new_n681), .ZN(new_n1114));
  NAND2_X1  g688(.A1(new_n1114), .A2(KEYINPUT127), .ZN(new_n1115));
  INV_X1    g689(.A(KEYINPUT127), .ZN(new_n1116));
  NAND4_X1  g690(.A1(new_n665), .A2(new_n1116), .A3(G319), .A4(new_n681), .ZN(new_n1117));
  NAND3_X1  g691(.A1(new_n1115), .A2(new_n703), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g692(.A(new_n1118), .ZN(new_n1119));
  OAI211_X1 g693(.A(new_n1119), .B(new_n866), .C1(new_n933), .C2(new_n934), .ZN(G225));
  INV_X1    g694(.A(G225), .ZN(G308));
endmodule


