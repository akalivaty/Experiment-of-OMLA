

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U556 ( .A(n551), .B(KEYINPUT65), .ZN(G160) );
  XOR2_X1 U557 ( .A(n776), .B(KEYINPUT89), .Z(n519) );
  AND2_X1 U558 ( .A1(G126), .A2(n888), .ZN(n520) );
  OR2_X1 U559 ( .A1(n757), .A2(n752), .ZN(n521) );
  AND2_X1 U560 ( .A1(n975), .A2(n823), .ZN(n522) );
  NOR2_X1 U561 ( .A1(n732), .A2(n731), .ZN(n523) );
  NOR2_X1 U562 ( .A1(n777), .A2(n519), .ZN(n524) );
  OR2_X1 U563 ( .A1(n714), .A2(n958), .ZN(n690) );
  XNOR2_X1 U564 ( .A(n714), .B(KEYINPUT91), .ZN(n709) );
  INV_X1 U565 ( .A(KEYINPUT32), .ZN(n748) );
  INV_X1 U566 ( .A(KEYINPUT87), .ZN(n715) );
  NOR2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n541) );
  NOR2_X1 U568 ( .A1(G2104), .A2(n544), .ZN(n888) );
  NOR2_X1 U569 ( .A1(n806), .A2(n522), .ZN(n807) );
  NOR2_X1 U570 ( .A1(n630), .A2(G651), .ZN(n642) );
  AND2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n887) );
  XOR2_X1 U572 ( .A(KEYINPUT1), .B(n525), .Z(n641) );
  XNOR2_X1 U573 ( .A(KEYINPUT6), .B(KEYINPUT76), .ZN(n529) );
  INV_X1 U574 ( .A(G651), .ZN(n532) );
  NOR2_X1 U575 ( .A1(G543), .A2(n532), .ZN(n525) );
  NAND2_X1 U576 ( .A1(G63), .A2(n641), .ZN(n527) );
  XOR2_X1 U577 ( .A(KEYINPUT0), .B(G543), .Z(n630) );
  NAND2_X1 U578 ( .A1(G51), .A2(n642), .ZN(n526) );
  NAND2_X1 U579 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U580 ( .A(n529), .B(n528), .ZN(n539) );
  NOR2_X1 U581 ( .A1(G543), .A2(G651), .ZN(n646) );
  NAND2_X1 U582 ( .A1(G89), .A2(n646), .ZN(n530) );
  XNOR2_X1 U583 ( .A(n530), .B(KEYINPUT4), .ZN(n531) );
  XNOR2_X1 U584 ( .A(n531), .B(KEYINPUT74), .ZN(n535) );
  OR2_X1 U585 ( .A1(n532), .A2(n630), .ZN(n533) );
  XNOR2_X1 U586 ( .A(KEYINPUT67), .B(n533), .ZN(n647) );
  NAND2_X1 U587 ( .A1(G76), .A2(n647), .ZN(n534) );
  NAND2_X1 U588 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U589 ( .A(KEYINPUT5), .B(n536), .ZN(n537) );
  XNOR2_X1 U590 ( .A(KEYINPUT75), .B(n537), .ZN(n538) );
  NOR2_X1 U591 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U592 ( .A(KEYINPUT7), .B(n540), .Z(G168) );
  XOR2_X2 U593 ( .A(KEYINPUT17), .B(n541), .Z(n892) );
  NAND2_X1 U594 ( .A1(G137), .A2(n892), .ZN(n543) );
  INV_X1 U595 ( .A(G2105), .ZN(n544) );
  NAND2_X1 U596 ( .A1(G125), .A2(n888), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n543), .A2(n542), .ZN(n547) );
  AND2_X1 U598 ( .A1(n544), .A2(G2104), .ZN(n891) );
  NAND2_X1 U599 ( .A1(G101), .A2(n891), .ZN(n545) );
  XNOR2_X1 U600 ( .A(KEYINPUT23), .B(n545), .ZN(n546) );
  NOR2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n550) );
  NAND2_X1 U602 ( .A1(n887), .A2(G113), .ZN(n548) );
  XNOR2_X1 U603 ( .A(n548), .B(KEYINPUT66), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U605 ( .A1(G64), .A2(n641), .ZN(n553) );
  NAND2_X1 U606 ( .A1(G52), .A2(n642), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n553), .A2(n552), .ZN(n559) );
  NAND2_X1 U608 ( .A1(G90), .A2(n646), .ZN(n555) );
  NAND2_X1 U609 ( .A1(G77), .A2(n647), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U611 ( .A(KEYINPUT69), .B(n556), .ZN(n557) );
  XNOR2_X1 U612 ( .A(KEYINPUT9), .B(n557), .ZN(n558) );
  NOR2_X1 U613 ( .A1(n559), .A2(n558), .ZN(G171) );
  NAND2_X1 U614 ( .A1(n892), .A2(G138), .ZN(n565) );
  NAND2_X1 U615 ( .A1(G114), .A2(n887), .ZN(n560) );
  XOR2_X1 U616 ( .A(KEYINPUT85), .B(n560), .Z(n562) );
  NAND2_X1 U617 ( .A1(G102), .A2(n891), .ZN(n561) );
  NAND2_X1 U618 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U619 ( .A1(n520), .A2(n563), .ZN(n564) );
  AND2_X1 U620 ( .A1(n565), .A2(n564), .ZN(G164) );
  AND2_X1 U621 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U622 ( .A(G57), .ZN(G237) );
  INV_X1 U623 ( .A(G132), .ZN(G219) );
  XOR2_X1 U624 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U625 ( .A1(G7), .A2(G661), .ZN(n566) );
  XNOR2_X1 U626 ( .A(n566), .B(KEYINPUT72), .ZN(n567) );
  XOR2_X1 U627 ( .A(KEYINPUT10), .B(n567), .Z(n922) );
  NAND2_X1 U628 ( .A1(n922), .A2(G567), .ZN(n568) );
  XOR2_X1 U629 ( .A(KEYINPUT11), .B(n568), .Z(G234) );
  NAND2_X1 U630 ( .A1(G56), .A2(n641), .ZN(n569) );
  XOR2_X1 U631 ( .A(KEYINPUT14), .B(n569), .Z(n575) );
  NAND2_X1 U632 ( .A1(n646), .A2(G81), .ZN(n570) );
  XNOR2_X1 U633 ( .A(n570), .B(KEYINPUT12), .ZN(n572) );
  NAND2_X1 U634 ( .A1(G68), .A2(n647), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U636 ( .A(KEYINPUT13), .B(n573), .Z(n574) );
  NOR2_X1 U637 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n642), .A2(G43), .ZN(n576) );
  NAND2_X1 U639 ( .A1(n577), .A2(n576), .ZN(n990) );
  INV_X1 U640 ( .A(G860), .ZN(n596) );
  OR2_X1 U641 ( .A1(n990), .A2(n596), .ZN(G153) );
  XNOR2_X1 U642 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U643 ( .A1(G868), .A2(G301), .ZN(n586) );
  NAND2_X1 U644 ( .A1(G66), .A2(n641), .ZN(n579) );
  NAND2_X1 U645 ( .A1(G92), .A2(n646), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U647 ( .A1(G79), .A2(n647), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G54), .A2(n642), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U651 ( .A(KEYINPUT15), .B(n584), .ZN(n971) );
  INV_X1 U652 ( .A(G868), .ZN(n661) );
  NAND2_X1 U653 ( .A1(n971), .A2(n661), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U655 ( .A1(G65), .A2(n641), .ZN(n588) );
  NAND2_X1 U656 ( .A1(G53), .A2(n642), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U658 ( .A1(G91), .A2(n646), .ZN(n590) );
  NAND2_X1 U659 ( .A1(G78), .A2(n647), .ZN(n589) );
  NAND2_X1 U660 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n970) );
  XOR2_X1 U662 ( .A(n970), .B(KEYINPUT70), .Z(G299) );
  XOR2_X1 U663 ( .A(KEYINPUT77), .B(n661), .Z(n593) );
  NOR2_X1 U664 ( .A1(G286), .A2(n593), .ZN(n595) );
  NOR2_X1 U665 ( .A1(G868), .A2(G299), .ZN(n594) );
  NOR2_X1 U666 ( .A1(n595), .A2(n594), .ZN(G297) );
  NAND2_X1 U667 ( .A1(n596), .A2(G559), .ZN(n597) );
  INV_X1 U668 ( .A(n971), .ZN(n697) );
  NAND2_X1 U669 ( .A1(n597), .A2(n697), .ZN(n598) );
  XNOR2_X1 U670 ( .A(n598), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U671 ( .A1(n971), .A2(n661), .ZN(n599) );
  XOR2_X1 U672 ( .A(KEYINPUT78), .B(n599), .Z(n600) );
  NOR2_X1 U673 ( .A1(G559), .A2(n600), .ZN(n602) );
  NOR2_X1 U674 ( .A1(G868), .A2(n990), .ZN(n601) );
  NOR2_X1 U675 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U676 ( .A1(G123), .A2(n888), .ZN(n603) );
  XNOR2_X1 U677 ( .A(n603), .B(KEYINPUT18), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n887), .A2(G111), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U680 ( .A1(G99), .A2(n891), .ZN(n607) );
  NAND2_X1 U681 ( .A1(G135), .A2(n892), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U683 ( .A1(n609), .A2(n608), .ZN(n939) );
  XNOR2_X1 U684 ( .A(n939), .B(G2096), .ZN(n610) );
  INV_X1 U685 ( .A(G2100), .ZN(n855) );
  NAND2_X1 U686 ( .A1(n610), .A2(n855), .ZN(G156) );
  NAND2_X1 U687 ( .A1(G93), .A2(n646), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G55), .A2(n642), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U690 ( .A1(G80), .A2(n647), .ZN(n613) );
  XNOR2_X1 U691 ( .A(KEYINPUT79), .B(n613), .ZN(n614) );
  NOR2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n641), .A2(G67), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n660) );
  NAND2_X1 U695 ( .A1(n697), .A2(G559), .ZN(n658) );
  XNOR2_X1 U696 ( .A(n990), .B(n658), .ZN(n618) );
  NOR2_X1 U697 ( .A1(G860), .A2(n618), .ZN(n619) );
  XOR2_X1 U698 ( .A(n660), .B(n619), .Z(G145) );
  NAND2_X1 U699 ( .A1(G85), .A2(n646), .ZN(n621) );
  NAND2_X1 U700 ( .A1(G47), .A2(n642), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U702 ( .A1(n641), .A2(G60), .ZN(n622) );
  XOR2_X1 U703 ( .A(KEYINPUT68), .B(n622), .Z(n623) );
  NOR2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n647), .A2(G72), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(G290) );
  NAND2_X1 U707 ( .A1(G49), .A2(n642), .ZN(n628) );
  NAND2_X1 U708 ( .A1(G74), .A2(G651), .ZN(n627) );
  NAND2_X1 U709 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U710 ( .A1(n641), .A2(n629), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n630), .A2(G87), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n632), .A2(n631), .ZN(G288) );
  XOR2_X1 U713 ( .A(KEYINPUT80), .B(KEYINPUT2), .Z(n634) );
  NAND2_X1 U714 ( .A1(G73), .A2(n647), .ZN(n633) );
  XNOR2_X1 U715 ( .A(n634), .B(n633), .ZN(n638) );
  NAND2_X1 U716 ( .A1(G86), .A2(n646), .ZN(n636) );
  NAND2_X1 U717 ( .A1(G48), .A2(n642), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n641), .A2(G61), .ZN(n639) );
  NAND2_X1 U721 ( .A1(n640), .A2(n639), .ZN(G305) );
  NAND2_X1 U722 ( .A1(G62), .A2(n641), .ZN(n644) );
  NAND2_X1 U723 ( .A1(G50), .A2(n642), .ZN(n643) );
  NAND2_X1 U724 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U725 ( .A(KEYINPUT81), .B(n645), .ZN(n651) );
  NAND2_X1 U726 ( .A1(G88), .A2(n646), .ZN(n649) );
  NAND2_X1 U727 ( .A1(G75), .A2(n647), .ZN(n648) );
  AND2_X1 U728 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U729 ( .A1(n651), .A2(n650), .ZN(G303) );
  XNOR2_X1 U730 ( .A(KEYINPUT19), .B(G290), .ZN(n652) );
  XNOR2_X1 U731 ( .A(n652), .B(G288), .ZN(n655) );
  XNOR2_X1 U732 ( .A(G299), .B(n990), .ZN(n653) );
  XNOR2_X1 U733 ( .A(n653), .B(n660), .ZN(n654) );
  XNOR2_X1 U734 ( .A(n655), .B(n654), .ZN(n657) );
  XOR2_X1 U735 ( .A(G305), .B(G303), .Z(n656) );
  XNOR2_X1 U736 ( .A(n657), .B(n656), .ZN(n910) );
  XNOR2_X1 U737 ( .A(n658), .B(n910), .ZN(n659) );
  NAND2_X1 U738 ( .A1(n659), .A2(G868), .ZN(n663) );
  NAND2_X1 U739 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U740 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U741 ( .A(KEYINPUT82), .B(n664), .ZN(G295) );
  NAND2_X1 U742 ( .A1(G2084), .A2(G2078), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n665), .B(KEYINPUT83), .ZN(n666) );
  XNOR2_X1 U744 ( .A(n666), .B(KEYINPUT20), .ZN(n667) );
  NAND2_X1 U745 ( .A1(n667), .A2(G2090), .ZN(n668) );
  XNOR2_X1 U746 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U747 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U748 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U749 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NOR2_X1 U750 ( .A1(G219), .A2(G220), .ZN(n670) );
  XOR2_X1 U751 ( .A(KEYINPUT22), .B(n670), .Z(n671) );
  NOR2_X1 U752 ( .A1(G218), .A2(n671), .ZN(n672) );
  NAND2_X1 U753 ( .A1(G96), .A2(n672), .ZN(n842) );
  NAND2_X1 U754 ( .A1(n842), .A2(G2106), .ZN(n676) );
  NAND2_X1 U755 ( .A1(G108), .A2(G120), .ZN(n673) );
  NOR2_X1 U756 ( .A1(G237), .A2(n673), .ZN(n674) );
  NAND2_X1 U757 ( .A1(G69), .A2(n674), .ZN(n843) );
  NAND2_X1 U758 ( .A1(n843), .A2(G567), .ZN(n675) );
  NAND2_X1 U759 ( .A1(n676), .A2(n675), .ZN(n866) );
  NAND2_X1 U760 ( .A1(G661), .A2(G483), .ZN(n677) );
  NOR2_X1 U761 ( .A1(n866), .A2(n677), .ZN(n841) );
  NAND2_X1 U762 ( .A1(n841), .A2(G36), .ZN(n678) );
  XNOR2_X1 U763 ( .A(KEYINPUT84), .B(n678), .ZN(G176) );
  INV_X1 U764 ( .A(G303), .ZN(G166) );
  XOR2_X1 U765 ( .A(KEYINPUT93), .B(KEYINPUT27), .Z(n683) );
  NAND2_X1 U766 ( .A1(G160), .A2(G40), .ZN(n779) );
  INV_X1 U767 ( .A(n779), .ZN(n681) );
  NOR2_X1 U768 ( .A1(G1384), .A2(G164), .ZN(n680) );
  XNOR2_X1 U769 ( .A(n680), .B(KEYINPUT64), .ZN(n778) );
  NAND2_X1 U770 ( .A1(n681), .A2(n778), .ZN(n714) );
  NAND2_X1 U771 ( .A1(G2072), .A2(n709), .ZN(n682) );
  XNOR2_X1 U772 ( .A(n683), .B(n682), .ZN(n685) );
  INV_X1 U773 ( .A(G1956), .ZN(n969) );
  NOR2_X1 U774 ( .A1(n709), .A2(n969), .ZN(n684) );
  NOR2_X1 U775 ( .A1(n685), .A2(n684), .ZN(n701) );
  NOR2_X1 U776 ( .A1(n970), .A2(n701), .ZN(n686) );
  XOR2_X1 U777 ( .A(n686), .B(KEYINPUT28), .Z(n705) );
  NAND2_X1 U778 ( .A1(n714), .A2(G1348), .ZN(n689) );
  NAND2_X1 U779 ( .A1(G2067), .A2(n709), .ZN(n687) );
  XOR2_X1 U780 ( .A(n687), .B(KEYINPUT95), .Z(n688) );
  NAND2_X1 U781 ( .A1(n689), .A2(n688), .ZN(n695) );
  XOR2_X1 U782 ( .A(G1996), .B(KEYINPUT94), .Z(n958) );
  XNOR2_X1 U783 ( .A(n690), .B(KEYINPUT26), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n714), .A2(G1341), .ZN(n691) );
  NAND2_X1 U785 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U786 ( .A1(n990), .A2(n693), .ZN(n698) );
  NAND2_X1 U787 ( .A1(n698), .A2(n697), .ZN(n694) );
  NAND2_X1 U788 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U789 ( .A(n696), .B(KEYINPUT96), .ZN(n700) );
  OR2_X1 U790 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U791 ( .A1(n700), .A2(n699), .ZN(n703) );
  NAND2_X1 U792 ( .A1(n970), .A2(n701), .ZN(n702) );
  NAND2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U794 ( .A1(n705), .A2(n704), .ZN(n707) );
  XNOR2_X1 U795 ( .A(KEYINPUT97), .B(KEYINPUT29), .ZN(n706) );
  XNOR2_X1 U796 ( .A(n707), .B(n706), .ZN(n713) );
  XNOR2_X1 U797 ( .A(G2078), .B(KEYINPUT25), .ZN(n708) );
  XNOR2_X1 U798 ( .A(n708), .B(KEYINPUT92), .ZN(n952) );
  NAND2_X1 U799 ( .A1(n709), .A2(n952), .ZN(n711) );
  INV_X1 U800 ( .A(G1961), .ZN(n997) );
  NAND2_X1 U801 ( .A1(n714), .A2(n997), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n723) );
  NAND2_X1 U803 ( .A1(n723), .A2(G171), .ZN(n712) );
  NAND2_X1 U804 ( .A1(n713), .A2(n712), .ZN(n740) );
  NAND2_X1 U805 ( .A1(n714), .A2(G8), .ZN(n716) );
  XNOR2_X1 U806 ( .A(n716), .B(n715), .ZN(n734) );
  NOR2_X1 U807 ( .A1(G1966), .A2(n734), .ZN(n717) );
  XNOR2_X1 U808 ( .A(KEYINPUT90), .B(n717), .ZN(n732) );
  INV_X1 U809 ( .A(G8), .ZN(n739) );
  NOR2_X1 U810 ( .A1(G2084), .A2(n714), .ZN(n730) );
  OR2_X1 U811 ( .A1(n739), .A2(n730), .ZN(n718) );
  NOR2_X1 U812 ( .A1(n732), .A2(n718), .ZN(n720) );
  INV_X1 U813 ( .A(KEYINPUT30), .ZN(n719) );
  XNOR2_X1 U814 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U815 ( .A1(n721), .A2(G168), .ZN(n722) );
  XNOR2_X1 U816 ( .A(n722), .B(KEYINPUT98), .ZN(n725) );
  NOR2_X1 U817 ( .A1(n723), .A2(G171), .ZN(n724) );
  NOR2_X1 U818 ( .A1(n725), .A2(n724), .ZN(n727) );
  INV_X1 U819 ( .A(KEYINPUT31), .ZN(n726) );
  XNOR2_X1 U820 ( .A(n727), .B(n726), .ZN(n741) );
  NAND2_X1 U821 ( .A1(n740), .A2(n741), .ZN(n729) );
  INV_X1 U822 ( .A(KEYINPUT99), .ZN(n728) );
  XNOR2_X1 U823 ( .A(n729), .B(n728), .ZN(n733) );
  AND2_X1 U824 ( .A1(n730), .A2(G8), .ZN(n731) );
  AND2_X1 U825 ( .A1(n733), .A2(n523), .ZN(n751) );
  NOR2_X1 U826 ( .A1(G2090), .A2(n714), .ZN(n736) );
  INV_X1 U827 ( .A(n734), .ZN(n771) );
  INV_X1 U828 ( .A(n771), .ZN(n775) );
  NOR2_X1 U829 ( .A1(G1971), .A2(n775), .ZN(n735) );
  NOR2_X1 U830 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U831 ( .A1(n737), .A2(G303), .ZN(n738) );
  OR2_X1 U832 ( .A1(n739), .A2(n738), .ZN(n743) );
  AND2_X1 U833 ( .A1(n740), .A2(n743), .ZN(n742) );
  NAND2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n747) );
  INV_X1 U835 ( .A(n743), .ZN(n745) );
  AND2_X1 U836 ( .A1(G286), .A2(G8), .ZN(n744) );
  OR2_X1 U837 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U838 ( .A1(n747), .A2(n746), .ZN(n749) );
  XNOR2_X1 U839 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X1 U840 ( .A1(n751), .A2(n750), .ZN(n768) );
  NOR2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n757) );
  NOR2_X1 U842 ( .A1(G1971), .A2(G303), .ZN(n752) );
  OR2_X1 U843 ( .A1(n768), .A2(n521), .ZN(n753) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n980) );
  NAND2_X1 U845 ( .A1(n753), .A2(n980), .ZN(n755) );
  NAND2_X1 U846 ( .A1(n771), .A2(KEYINPUT100), .ZN(n754) );
  NOR2_X1 U847 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U848 ( .A1(KEYINPUT33), .A2(n756), .ZN(n763) );
  INV_X1 U849 ( .A(n757), .ZN(n981) );
  OR2_X1 U850 ( .A1(KEYINPUT100), .A2(n981), .ZN(n760) );
  NAND2_X1 U851 ( .A1(n757), .A2(KEYINPUT33), .ZN(n758) );
  NAND2_X1 U852 ( .A1(n758), .A2(KEYINPUT100), .ZN(n759) );
  NAND2_X1 U853 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U854 ( .A1(n775), .A2(n761), .ZN(n762) );
  NOR2_X1 U855 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U856 ( .A(G1981), .B(G305), .Z(n977) );
  NAND2_X1 U857 ( .A1(n764), .A2(n977), .ZN(n765) );
  NAND2_X1 U858 ( .A1(G166), .A2(G8), .ZN(n766) );
  NOR2_X1 U859 ( .A1(G2090), .A2(n766), .ZN(n767) );
  NOR2_X1 U860 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U861 ( .A(KEYINPUT101), .B(n769), .Z(n770) );
  NOR2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n777) );
  NOR2_X1 U863 ( .A1(G1981), .A2(G305), .ZN(n772) );
  XOR2_X1 U864 ( .A(KEYINPUT88), .B(n772), .Z(n773) );
  XNOR2_X1 U865 ( .A(KEYINPUT24), .B(n773), .ZN(n774) );
  NOR2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U867 ( .A1(n765), .A2(n524), .ZN(n808) );
  NOR2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n823) );
  NAND2_X1 U869 ( .A1(G104), .A2(n891), .ZN(n781) );
  NAND2_X1 U870 ( .A1(G140), .A2(n892), .ZN(n780) );
  NAND2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U872 ( .A(KEYINPUT34), .B(n782), .ZN(n787) );
  NAND2_X1 U873 ( .A1(G116), .A2(n887), .ZN(n784) );
  NAND2_X1 U874 ( .A1(G128), .A2(n888), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U876 ( .A(KEYINPUT35), .B(n785), .Z(n786) );
  NOR2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U878 ( .A(KEYINPUT36), .B(n788), .ZN(n884) );
  XNOR2_X1 U879 ( .A(G2067), .B(KEYINPUT37), .ZN(n821) );
  NOR2_X1 U880 ( .A1(n884), .A2(n821), .ZN(n932) );
  NAND2_X1 U881 ( .A1(n823), .A2(n932), .ZN(n819) );
  NAND2_X1 U882 ( .A1(G129), .A2(n888), .ZN(n790) );
  NAND2_X1 U883 ( .A1(G141), .A2(n892), .ZN(n789) );
  NAND2_X1 U884 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U885 ( .A1(n891), .A2(G105), .ZN(n791) );
  XOR2_X1 U886 ( .A(KEYINPUT38), .B(n791), .Z(n792) );
  NOR2_X1 U887 ( .A1(n793), .A2(n792), .ZN(n795) );
  NAND2_X1 U888 ( .A1(n887), .A2(G117), .ZN(n794) );
  NAND2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n898) );
  AND2_X1 U890 ( .A1(n898), .A2(G1996), .ZN(n804) );
  NAND2_X1 U891 ( .A1(G107), .A2(n887), .ZN(n797) );
  NAND2_X1 U892 ( .A1(G119), .A2(n888), .ZN(n796) );
  NAND2_X1 U893 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U894 ( .A(KEYINPUT86), .B(n798), .ZN(n802) );
  NAND2_X1 U895 ( .A1(G95), .A2(n891), .ZN(n800) );
  NAND2_X1 U896 ( .A1(G131), .A2(n892), .ZN(n799) );
  NAND2_X1 U897 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n883) );
  INV_X1 U899 ( .A(G1991), .ZN(n846) );
  NOR2_X1 U900 ( .A1(n883), .A2(n846), .ZN(n803) );
  NOR2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n936) );
  INV_X1 U902 ( .A(n936), .ZN(n805) );
  NAND2_X1 U903 ( .A1(n805), .A2(n823), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n819), .A2(n810), .ZN(n806) );
  XNOR2_X1 U905 ( .A(G1986), .B(G290), .ZN(n975) );
  NAND2_X1 U906 ( .A1(n808), .A2(n807), .ZN(n826) );
  XOR2_X1 U907 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n809) );
  XNOR2_X1 U908 ( .A(KEYINPUT104), .B(n809), .ZN(n818) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n898), .ZN(n929) );
  INV_X1 U910 ( .A(n810), .ZN(n815) );
  AND2_X1 U911 ( .A1(n846), .A2(n883), .ZN(n811) );
  XOR2_X1 U912 ( .A(KEYINPUT103), .B(n811), .Z(n940) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n812) );
  XNOR2_X1 U914 ( .A(KEYINPUT102), .B(n812), .ZN(n813) );
  NOR2_X1 U915 ( .A1(n940), .A2(n813), .ZN(n814) );
  NOR2_X1 U916 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U917 ( .A1(n929), .A2(n816), .ZN(n817) );
  XNOR2_X1 U918 ( .A(n818), .B(n817), .ZN(n820) );
  NAND2_X1 U919 ( .A1(n820), .A2(n819), .ZN(n822) );
  NAND2_X1 U920 ( .A1(n884), .A2(n821), .ZN(n935) );
  NAND2_X1 U921 ( .A1(n822), .A2(n935), .ZN(n824) );
  NAND2_X1 U922 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U923 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U924 ( .A(n827), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U925 ( .A(G2443), .B(G2451), .ZN(n837) );
  XOR2_X1 U926 ( .A(G2446), .B(G2430), .Z(n829) );
  XNOR2_X1 U927 ( .A(KEYINPUT107), .B(G2438), .ZN(n828) );
  XNOR2_X1 U928 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U929 ( .A(G2435), .B(G2454), .Z(n831) );
  XNOR2_X1 U930 ( .A(G1341), .B(G1348), .ZN(n830) );
  XNOR2_X1 U931 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U932 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U933 ( .A(G2427), .B(KEYINPUT106), .ZN(n834) );
  XNOR2_X1 U934 ( .A(n835), .B(n834), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(n838) );
  NAND2_X1 U936 ( .A1(n838), .A2(G14), .ZN(n917) );
  XOR2_X1 U937 ( .A(KEYINPUT108), .B(n917), .Z(G401) );
  NAND2_X1 U938 ( .A1(G2106), .A2(n922), .ZN(G217) );
  AND2_X1 U939 ( .A1(G15), .A2(G2), .ZN(n839) );
  NAND2_X1 U940 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U941 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U942 ( .A1(n841), .A2(n840), .ZN(G188) );
  XNOR2_X1 U943 ( .A(G120), .B(KEYINPUT109), .ZN(G236) );
  INV_X1 U945 ( .A(G108), .ZN(G238) );
  INV_X1 U946 ( .A(G96), .ZN(G221) );
  NOR2_X1 U947 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U948 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U949 ( .A(G1976), .B(KEYINPUT41), .ZN(n854) );
  XNOR2_X1 U950 ( .A(G1971), .B(n997), .ZN(n845) );
  XOR2_X1 U951 ( .A(G1986), .B(n969), .Z(n844) );
  XNOR2_X1 U952 ( .A(n845), .B(n844), .ZN(n850) );
  XOR2_X1 U953 ( .A(G1966), .B(G1981), .Z(n848) );
  XOR2_X1 U954 ( .A(G1996), .B(n846), .Z(n847) );
  XNOR2_X1 U955 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U956 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U957 ( .A(KEYINPUT112), .B(G2474), .ZN(n851) );
  XNOR2_X1 U958 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U959 ( .A(n854), .B(n853), .ZN(G229) );
  XNOR2_X1 U960 ( .A(n855), .B(KEYINPUT110), .ZN(n857) );
  XNOR2_X1 U961 ( .A(KEYINPUT111), .B(KEYINPUT43), .ZN(n856) );
  XNOR2_X1 U962 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U963 ( .A(KEYINPUT42), .B(G2090), .Z(n859) );
  XNOR2_X1 U964 ( .A(G2067), .B(G2072), .ZN(n858) );
  XNOR2_X1 U965 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U966 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U967 ( .A(G2678), .B(G2096), .ZN(n862) );
  XNOR2_X1 U968 ( .A(n863), .B(n862), .ZN(n865) );
  XOR2_X1 U969 ( .A(G2084), .B(G2078), .Z(n864) );
  XNOR2_X1 U970 ( .A(n865), .B(n864), .ZN(G227) );
  INV_X1 U971 ( .A(n866), .ZN(G319) );
  NAND2_X1 U972 ( .A1(G124), .A2(n888), .ZN(n867) );
  XNOR2_X1 U973 ( .A(n867), .B(KEYINPUT44), .ZN(n869) );
  NAND2_X1 U974 ( .A1(n887), .A2(G112), .ZN(n868) );
  NAND2_X1 U975 ( .A1(n869), .A2(n868), .ZN(n873) );
  NAND2_X1 U976 ( .A1(G100), .A2(n891), .ZN(n871) );
  NAND2_X1 U977 ( .A1(G136), .A2(n892), .ZN(n870) );
  NAND2_X1 U978 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U979 ( .A1(n873), .A2(n872), .ZN(G162) );
  NAND2_X1 U980 ( .A1(G103), .A2(n891), .ZN(n875) );
  NAND2_X1 U981 ( .A1(G139), .A2(n892), .ZN(n874) );
  NAND2_X1 U982 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U983 ( .A(KEYINPUT113), .B(n876), .Z(n882) );
  NAND2_X1 U984 ( .A1(n888), .A2(G127), .ZN(n877) );
  XNOR2_X1 U985 ( .A(n877), .B(KEYINPUT114), .ZN(n879) );
  NAND2_X1 U986 ( .A1(G115), .A2(n887), .ZN(n878) );
  NAND2_X1 U987 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  NOR2_X1 U989 ( .A1(n882), .A2(n881), .ZN(n923) );
  XNOR2_X1 U990 ( .A(n923), .B(G162), .ZN(n886) );
  XNOR2_X1 U991 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U992 ( .A(n886), .B(n885), .ZN(n901) );
  NAND2_X1 U993 ( .A1(G118), .A2(n887), .ZN(n890) );
  NAND2_X1 U994 ( .A1(G130), .A2(n888), .ZN(n889) );
  NAND2_X1 U995 ( .A1(n890), .A2(n889), .ZN(n897) );
  NAND2_X1 U996 ( .A1(G106), .A2(n891), .ZN(n894) );
  NAND2_X1 U997 ( .A1(G142), .A2(n892), .ZN(n893) );
  NAND2_X1 U998 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U999 ( .A(n895), .B(KEYINPUT45), .Z(n896) );
  NOR2_X1 U1000 ( .A1(n897), .A2(n896), .ZN(n899) );
  XNOR2_X1 U1001 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U1002 ( .A(n901), .B(n900), .Z(n908) );
  XNOR2_X1 U1003 ( .A(n939), .B(KEYINPUT115), .ZN(n902) );
  XNOR2_X1 U1004 ( .A(n902), .B(KEYINPUT116), .ZN(n903) );
  XOR2_X1 U1005 ( .A(n903), .B(KEYINPUT46), .Z(n905) );
  XNOR2_X1 U1006 ( .A(G160), .B(KEYINPUT48), .ZN(n904) );
  XNOR2_X1 U1007 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1008 ( .A(G164), .B(n906), .ZN(n907) );
  XNOR2_X1 U1009 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n909), .ZN(G395) );
  XOR2_X1 U1011 ( .A(KEYINPUT117), .B(n910), .Z(n912) );
  XOR2_X1 U1012 ( .A(n971), .B(G286), .Z(n911) );
  XNOR2_X1 U1013 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1014 ( .A(G171), .B(n913), .Z(n914) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n914), .ZN(G397) );
  NOR2_X1 U1016 ( .A1(G229), .A2(G227), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(KEYINPUT118), .ZN(n915) );
  XNOR2_X1 U1018 ( .A(n916), .B(n915), .ZN(n919) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n917), .ZN(n918) );
  NOR2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(G69), .ZN(G235) );
  INV_X1 U1025 ( .A(n922), .ZN(G223) );
  XOR2_X1 U1026 ( .A(G2072), .B(n923), .Z(n925) );
  XOR2_X1 U1027 ( .A(G164), .B(G2078), .Z(n924) );
  NOR2_X1 U1028 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1029 ( .A(KEYINPUT120), .B(n926), .ZN(n927) );
  XNOR2_X1 U1030 ( .A(n927), .B(KEYINPUT50), .ZN(n934) );
  XOR2_X1 U1031 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1032 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1033 ( .A(n930), .B(KEYINPUT51), .ZN(n931) );
  NOR2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n945) );
  NAND2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n938) );
  XOR2_X1 U1037 ( .A(G160), .B(G2084), .Z(n937) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n943) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1040 ( .A(KEYINPUT119), .B(n941), .Z(n942) );
  NAND2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(KEYINPUT52), .B(n946), .ZN(n947) );
  INV_X1 U1044 ( .A(KEYINPUT55), .ZN(n1025) );
  NAND2_X1 U1045 ( .A1(n947), .A2(n1025), .ZN(n948) );
  NAND2_X1 U1046 ( .A1(n948), .A2(G29), .ZN(n1032) );
  XNOR2_X1 U1047 ( .A(G2090), .B(G35), .ZN(n963) );
  XNOR2_X1 U1048 ( .A(G2067), .B(G26), .ZN(n950) );
  XNOR2_X1 U1049 ( .A(G33), .B(G2072), .ZN(n949) );
  NOR2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n957) );
  XOR2_X1 U1051 ( .A(G25), .B(G1991), .Z(n951) );
  NAND2_X1 U1052 ( .A1(n951), .A2(G28), .ZN(n955) );
  XNOR2_X1 U1053 ( .A(G27), .B(n952), .ZN(n953) );
  XNOR2_X1 U1054 ( .A(KEYINPUT121), .B(n953), .ZN(n954) );
  NOR2_X1 U1055 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n960) );
  XOR2_X1 U1057 ( .A(n958), .B(G32), .Z(n959) );
  NOR2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1059 ( .A(KEYINPUT53), .B(n961), .ZN(n962) );
  NOR2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1061 ( .A(G2084), .B(KEYINPUT54), .Z(n964) );
  XNOR2_X1 U1062 ( .A(G34), .B(n964), .ZN(n965) );
  NAND2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n1026) );
  NOR2_X1 U1064 ( .A1(G29), .A2(KEYINPUT55), .ZN(n967) );
  NAND2_X1 U1065 ( .A1(n1026), .A2(n967), .ZN(n968) );
  NAND2_X1 U1066 ( .A1(G11), .A2(n968), .ZN(n1030) );
  INV_X1 U1067 ( .A(G16), .ZN(n1021) );
  XOR2_X1 U1068 ( .A(n1021), .B(KEYINPUT56), .Z(n996) );
  XOR2_X1 U1069 ( .A(n970), .B(n969), .Z(n973) );
  XOR2_X1 U1070 ( .A(n971), .B(G1348), .Z(n972) );
  NAND2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n994) );
  XNOR2_X1 U1073 ( .A(G1966), .B(G168), .ZN(n976) );
  XNOR2_X1 U1074 ( .A(n976), .B(KEYINPUT122), .ZN(n978) );
  NAND2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1076 ( .A(n979), .B(KEYINPUT57), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1078 ( .A(n982), .B(KEYINPUT123), .ZN(n985) );
  XOR2_X1 U1079 ( .A(G303), .B(G1971), .Z(n983) );
  XNOR2_X1 U1080 ( .A(n983), .B(KEYINPUT124), .ZN(n984) );
  NAND2_X1 U1081 ( .A1(n985), .A2(n984), .ZN(n987) );
  XNOR2_X1 U1082 ( .A(G171), .B(n997), .ZN(n986) );
  NOR2_X1 U1083 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(G1341), .B(n990), .ZN(n991) );
  NOR2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n1023) );
  XNOR2_X1 U1089 ( .A(G1966), .B(G21), .ZN(n999) );
  XOR2_X1 U1090 ( .A(n997), .B(G5), .Z(n998) );
  NOR2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1010) );
  XOR2_X1 U1092 ( .A(G1341), .B(G19), .Z(n1001) );
  XOR2_X1 U1093 ( .A(G1956), .B(G20), .Z(n1000) );
  NAND2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1007) );
  XOR2_X1 U1095 ( .A(G1981), .B(G6), .Z(n1005) );
  XOR2_X1 U1096 ( .A(KEYINPUT59), .B(G4), .Z(n1002) );
  XNOR2_X1 U1097 ( .A(KEYINPUT125), .B(n1002), .ZN(n1003) );
  XNOR2_X1 U1098 ( .A(n1003), .B(G1348), .ZN(n1004) );
  NAND2_X1 U1099 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1101 ( .A(n1008), .B(KEYINPUT60), .ZN(n1009) );
  NAND2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(G1976), .B(G23), .ZN(n1012) );
  XNOR2_X1 U1104 ( .A(G1971), .B(G22), .ZN(n1011) );
  NOR2_X1 U1105 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XOR2_X1 U1106 ( .A(G1986), .B(G24), .Z(n1013) );
  NAND2_X1 U1107 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1108 ( .A(KEYINPUT58), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1109 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1110 ( .A(n1018), .B(KEYINPUT61), .ZN(n1019) );
  XNOR2_X1 U1111 ( .A(n1019), .B(KEYINPUT126), .ZN(n1020) );
  NAND2_X1 U1112 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1113 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1114 ( .A(n1024), .B(KEYINPUT127), .ZN(n1028) );
  OR2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1033), .ZN(G150) );
  INV_X1 U1120 ( .A(G150), .ZN(G311) );
endmodule

