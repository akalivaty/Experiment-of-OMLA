//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012, new_n1013;
  INV_X1    g000(.A(KEYINPUT99), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G228gat), .A2(G233gat), .ZN(new_n205));
  AND2_X1   g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G155gat), .B(G162gat), .ZN(new_n209));
  INV_X1    g008(.A(G155gat), .ZN(new_n210));
  INV_X1    g009(.A(G162gat), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT2), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n208), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G141gat), .ZN(new_n214));
  INV_X1    g013(.A(G148gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n213), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT29), .ZN(new_n225));
  NAND2_X1  g024(.A1(G211gat), .A2(G218gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT22), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G204gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G197gat), .ZN(new_n230));
  INV_X1    g029(.A(G197gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G204gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n228), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(G211gat), .B(G218gat), .Z(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G211gat), .B(G218gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(G197gat), .B(G204gat), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n236), .B1(new_n228), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n225), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n224), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n233), .A2(new_n234), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n236), .A2(new_n237), .A3(new_n228), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n213), .A2(new_n223), .A3(new_n240), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n244), .B1(new_n245), .B2(new_n225), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n205), .B1(new_n241), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G22gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n225), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n244), .A2(KEYINPUT71), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n242), .A2(new_n251), .A3(new_n243), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n205), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n213), .A2(new_n223), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT29), .B1(new_n242), .B2(new_n243), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n255), .B1(new_n256), .B2(KEYINPUT3), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n253), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n247), .A2(new_n248), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n248), .B1(new_n247), .B2(new_n258), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n204), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n253), .A2(new_n254), .A3(new_n257), .ZN(new_n262));
  INV_X1    g061(.A(new_n246), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n254), .B1(new_n263), .B2(new_n257), .ZN(new_n264));
  OAI21_X1  g063(.A(G22gat), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n247), .A2(new_n258), .A3(new_n248), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n266), .A3(new_n203), .ZN(new_n267));
  XOR2_X1   g066(.A(KEYINPUT31), .B(G50gat), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n261), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n269), .B1(new_n261), .B2(new_n267), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(G8gat), .B(G36gat), .Z(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT73), .ZN(new_n274));
  XNOR2_X1  g073(.A(G64gat), .B(G92gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n250), .A2(new_n252), .ZN(new_n277));
  INV_X1    g076(.A(G226gat), .ZN(new_n278));
  INV_X1    g077(.A(G233gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n282), .B1(KEYINPUT23), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G169gat), .ZN(new_n285));
  INV_X1    g084(.A(G176gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT23), .ZN(new_n287));
  INV_X1    g086(.A(G190gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  OR2_X1    g090(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(G190gat), .A3(new_n293), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n291), .A2(KEYINPUT64), .A3(KEYINPUT25), .A4(new_n294), .ZN(new_n295));
  AND2_X1   g094(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n288), .A2(new_n296), .B1(new_n282), .B2(KEYINPUT23), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n283), .A2(KEYINPUT23), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n285), .A2(new_n286), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n297), .A2(new_n294), .A3(new_n300), .A4(KEYINPUT25), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT64), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n297), .A2(new_n294), .A3(new_n300), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n295), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n299), .A2(KEYINPUT26), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT26), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n282), .B1(new_n310), .B2(new_n283), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT27), .B(G183gat), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n312), .A2(KEYINPUT28), .A3(new_n288), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT28), .B1(new_n312), .B2(new_n288), .ZN(new_n314));
  OAI221_X1 g113(.A(new_n308), .B1(new_n309), .B2(new_n311), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n281), .B1(new_n307), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n307), .A2(new_n315), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n280), .B1(new_n317), .B2(new_n225), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT72), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT29), .B1(new_n307), .B2(new_n315), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT72), .B1(new_n321), .B2(new_n280), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n277), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n244), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n318), .A2(new_n316), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n276), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n317), .A2(new_n225), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(new_n319), .A3(new_n281), .ZN(new_n328));
  INV_X1    g127(.A(new_n316), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(new_n322), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n277), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n325), .ZN(new_n333));
  INV_X1    g132(.A(new_n276), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n326), .A2(new_n335), .A3(KEYINPUT30), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n337));
  INV_X1    g136(.A(G134gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G127gat), .ZN(new_n339));
  INV_X1    g138(.A(G127gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G134gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G113gat), .B(G120gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n342), .B1(new_n343), .B2(KEYINPUT1), .ZN(new_n344));
  INV_X1    g143(.A(G120gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G113gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT65), .B(G113gat), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n347), .B1(new_n348), .B2(G120gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT1), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n339), .A2(new_n341), .A3(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n344), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n337), .A2(new_n352), .A3(new_n245), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT4), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n352), .B2(new_n255), .ZN(new_n355));
  INV_X1    g154(.A(G113gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT65), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT65), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G113gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n359), .A3(G120gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n346), .ZN(new_n361));
  INV_X1    g160(.A(new_n351), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n356), .A2(G120gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n350), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n361), .A2(new_n362), .B1(new_n365), .B2(new_n342), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n224), .ZN(new_n367));
  XOR2_X1   g166(.A(KEYINPUT74), .B(KEYINPUT4), .Z(new_n368));
  OAI211_X1 g167(.A(new_n353), .B(new_n355), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G225gat), .A2(G233gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT39), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n352), .A2(new_n255), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n361), .A2(new_n362), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n375), .A2(new_n344), .B1(new_n223), .B2(new_n213), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n373), .B1(new_n377), .B2(new_n370), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n369), .A2(new_n373), .A3(new_n371), .ZN(new_n380));
  XNOR2_X1  g179(.A(G1gat), .B(G29gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT0), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT77), .ZN(new_n383));
  XNOR2_X1  g182(.A(G57gat), .B(G85gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT77), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n382), .B(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n384), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n380), .A2(KEYINPUT78), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT78), .B1(new_n380), .B2(new_n390), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n379), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT40), .ZN(new_n394));
  OR2_X1    g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n368), .B1(new_n352), .B2(new_n255), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n366), .A2(new_n224), .A3(KEYINPUT4), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n398), .A2(KEYINPUT75), .A3(new_n353), .A4(new_n370), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n353), .A2(new_n396), .A3(new_n397), .A4(new_n370), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT75), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g202(.A(KEYINPUT76), .B(new_n371), .C1(new_n374), .C2(new_n376), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT5), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n352), .A2(new_n255), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n370), .B1(new_n367), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(KEYINPUT76), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n369), .A2(KEYINPUT5), .A3(new_n371), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n390), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n393), .A2(new_n394), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n325), .B1(new_n330), .B2(new_n331), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT30), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(new_n417), .A3(new_n334), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n336), .A2(new_n395), .A3(new_n415), .A4(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT79), .B(KEYINPUT37), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n332), .A2(new_n333), .A3(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n328), .A2(new_n322), .A3(new_n329), .A4(new_n277), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n324), .B1(new_n318), .B2(new_n316), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT37), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT38), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n421), .A2(new_n425), .A3(new_n426), .A4(new_n276), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n413), .A2(KEYINPUT6), .A3(new_n414), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n411), .B1(new_n403), .B2(new_n409), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT6), .B1(new_n429), .B2(new_n390), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT5), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n431), .B1(new_n407), .B2(KEYINPUT76), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT76), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n433), .B1(new_n377), .B2(new_n370), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n402), .B2(new_n399), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n414), .B1(new_n436), .B2(new_n411), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n430), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n427), .A2(new_n428), .A3(new_n438), .A4(new_n335), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n334), .B1(new_n416), .B2(new_n420), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT37), .B1(new_n323), .B2(new_n325), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n426), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n272), .B(new_n419), .C1(new_n439), .C2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT80), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n438), .A2(new_n428), .A3(new_n335), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n440), .A2(new_n441), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT38), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n448), .A3(new_n427), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n449), .A2(KEYINPUT80), .A3(new_n272), .A4(new_n419), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n336), .A2(new_n418), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n438), .A2(new_n428), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n272), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n317), .A2(new_n366), .ZN(new_n457));
  INV_X1    g256(.A(G227gat), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n458), .A2(new_n279), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n307), .A2(new_n352), .A3(new_n315), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  XOR2_X1   g260(.A(G15gat), .B(G43gat), .Z(new_n462));
  XNOR2_X1  g261(.A(G71gat), .B(G99gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT33), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n461), .A2(KEYINPUT32), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT66), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n461), .A2(KEYINPUT66), .A3(KEYINPUT32), .A4(new_n465), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n461), .A2(KEYINPUT32), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT33), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n461), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n473), .A3(new_n464), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n460), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n352), .B1(new_n307), .B2(new_n315), .ZN(new_n477));
  OAI22_X1  g276(.A1(new_n476), .A2(new_n477), .B1(new_n458), .B2(new_n279), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT68), .B1(new_n478), .B2(KEYINPUT34), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n459), .B1(new_n457), .B2(new_n460), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT68), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT34), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n478), .A2(KEYINPUT34), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n479), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n475), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n483), .A2(new_n484), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n470), .A2(new_n487), .A3(new_n479), .A4(new_n474), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT70), .B(KEYINPUT36), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n470), .A2(KEYINPUT67), .A3(new_n474), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT67), .B1(new_n470), .B2(new_n474), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n485), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT69), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n488), .A2(KEYINPUT36), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n495), .B1(new_n494), .B2(new_n496), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n491), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n451), .A2(new_n456), .A3(new_n499), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n336), .A2(new_n418), .B1(new_n438), .B2(new_n428), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n272), .A2(new_n488), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(new_n494), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT35), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT82), .ZN(new_n505));
  XOR2_X1   g304(.A(KEYINPUT81), .B(KEYINPUT35), .Z(new_n506));
  NAND4_X1  g305(.A1(new_n486), .A2(new_n272), .A3(new_n488), .A4(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n505), .B1(new_n508), .B2(new_n501), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n454), .A2(new_n507), .A3(KEYINPUT82), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n500), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT88), .ZN(new_n513));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514));
  OR3_X1    g313(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n515), .A2(new_n516), .B1(G29gat), .B2(G36gat), .ZN(new_n517));
  INV_X1    g316(.A(G43gat), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT15), .B1(new_n518), .B2(G50gat), .ZN(new_n519));
  INV_X1    g318(.A(G50gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(G43gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT83), .B(G43gat), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n521), .B1(new_n524), .B2(new_n520), .ZN(new_n525));
  OAI22_X1  g324(.A1(new_n525), .A2(KEYINPUT15), .B1(new_n521), .B2(new_n519), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n523), .B1(new_n526), .B2(new_n517), .ZN(new_n527));
  XNOR2_X1  g326(.A(G15gat), .B(G22gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT16), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n528), .B1(new_n529), .B2(G1gat), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(G1gat), .B2(new_n528), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT85), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT84), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n533), .B(G8gat), .C1(KEYINPUT84), .C2(new_n531), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT86), .ZN(new_n535));
  INV_X1    g334(.A(G8gat), .ZN(new_n536));
  OAI211_X1 g335(.A(KEYINPUT84), .B(new_n536), .C1(new_n531), .C2(new_n532), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n527), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT86), .B1(new_n527), .B2(new_n539), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n541), .B1(new_n537), .B2(new_n534), .ZN(new_n542));
  OAI211_X1 g341(.A(KEYINPUT18), .B(new_n514), .C1(new_n540), .C2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT87), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n514), .B1(new_n540), .B2(new_n542), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT18), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n514), .B(KEYINPUT13), .Z(new_n547));
  NAND2_X1  g346(.A1(new_n534), .A2(new_n537), .ZN(new_n548));
  INV_X1    g347(.A(new_n527), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n545), .A2(new_n546), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT11), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(new_n285), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(G197gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT12), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n551), .A3(new_n557), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  OR3_X1    g361(.A1(new_n512), .A2(new_n513), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n513), .B1(new_n512), .B2(new_n562), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n453), .ZN(new_n566));
  XNOR2_X1  g365(.A(G190gat), .B(G218gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT8), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(G85gat), .B2(G92gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(G85gat), .A2(G92gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT94), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT7), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G99gat), .B(G106gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT94), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n571), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT7), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n575), .B1(new_n574), .B2(new_n578), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n539), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n582), .A2(new_n527), .B1(KEYINPUT41), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n582), .A2(new_n527), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n567), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n567), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n584), .B(new_n588), .C1(new_n527), .C2(new_n582), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n583), .A2(KEYINPUT41), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n587), .B(new_n589), .C1(KEYINPUT41), .C2(new_n583), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G134gat), .B(G162gat), .Z(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n595), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n592), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G183gat), .B(G211gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G127gat), .B(G155gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT89), .ZN(new_n606));
  XOR2_X1   g405(.A(G71gat), .B(G78gat), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G57gat), .B(G64gat), .Z(new_n609));
  NAND3_X1  g408(.A1(new_n606), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(KEYINPUT9), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n607), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT90), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT21), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n610), .A2(KEYINPUT90), .A3(new_n612), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT91), .ZN(new_n619));
  NAND2_X1  g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT91), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n615), .A2(new_n622), .A3(new_n616), .A4(new_n617), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n619), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n621), .B1(new_n619), .B2(new_n623), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n604), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n610), .A2(KEYINPUT90), .A3(new_n612), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT90), .B1(new_n610), .B2(new_n612), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n622), .B1(new_n629), .B2(new_n616), .ZN(new_n630));
  INV_X1    g429(.A(new_n623), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n620), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n619), .A2(new_n621), .A3(new_n623), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n632), .A2(new_n633), .A3(new_n603), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n626), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n636), .B1(new_n626), .B2(new_n634), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n602), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n615), .A2(new_n617), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT92), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n640), .A2(new_n641), .ZN(new_n644));
  OAI21_X1  g443(.A(KEYINPUT21), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n548), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n646), .B(KEYINPUT93), .Z(new_n647));
  NOR3_X1   g446(.A1(new_n624), .A2(new_n625), .A3(new_n604), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n603), .B1(new_n632), .B2(new_n633), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n635), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n626), .A2(new_n634), .A3(new_n636), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(new_n651), .A3(new_n601), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n639), .A2(new_n647), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n647), .B1(new_n639), .B2(new_n652), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n600), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT95), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n639), .A2(new_n652), .ZN(new_n658));
  INV_X1    g457(.A(new_n647), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n639), .A2(new_n652), .A3(new_n647), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(KEYINPUT95), .A3(new_n600), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n615), .B(new_n617), .C1(new_n580), .C2(new_n581), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT10), .ZN(new_n666));
  INV_X1    g465(.A(new_n581), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n667), .A2(new_n612), .A3(new_n610), .A4(new_n579), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT96), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT96), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n665), .A2(new_n671), .A3(new_n668), .A4(new_n666), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n580), .A2(new_n581), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT10), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n629), .A2(KEYINPUT92), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n675), .B1(new_n676), .B2(new_n642), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(G230gat), .A2(G233gat), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n680), .B1(new_n665), .B2(new_n668), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT97), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G120gat), .B(G148gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(G176gat), .B(G204gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n687), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n681), .A2(new_n689), .A3(new_n683), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n664), .A2(new_n691), .ZN(new_n692));
  AND4_X1   g491(.A1(new_n202), .A2(new_n565), .A3(new_n566), .A4(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n692), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n563), .B2(new_n564), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n202), .B1(new_n695), .B2(new_n566), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT98), .B(G1gat), .Z(new_n697));
  OR3_X1    g496(.A1(new_n693), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n697), .B1(new_n693), .B2(new_n696), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(G1324gat));
  INV_X1    g499(.A(new_n695), .ZN(new_n701));
  OAI21_X1  g500(.A(G8gat), .B1(new_n701), .B2(new_n452), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n703));
  INV_X1    g502(.A(new_n452), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT16), .B(G8gat), .Z(new_n705));
  NAND3_X1  g504(.A1(new_n695), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n706), .A2(new_n707), .A3(new_n703), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n706), .B2(new_n703), .ZN(new_n709));
  OAI221_X1 g508(.A(new_n702), .B1(new_n703), .B2(new_n706), .C1(new_n708), .C2(new_n709), .ZN(G1325gat));
  OR3_X1    g509(.A1(new_n701), .A2(G15gat), .A3(new_n489), .ZN(new_n711));
  OAI21_X1  g510(.A(G15gat), .B1(new_n701), .B2(new_n499), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(G1326gat));
  OAI21_X1  g512(.A(KEYINPUT101), .B1(new_n701), .B2(new_n272), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT101), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n695), .A2(new_n715), .A3(new_n455), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT43), .B(G22gat), .Z(new_n717));
  AND3_X1   g516(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n714), .B2(new_n716), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(G1327gat));
  NOR2_X1   g519(.A1(new_n662), .A2(new_n691), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n600), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n724), .B1(new_n563), .B2(new_n564), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n453), .A2(G29gat), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT102), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT102), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n725), .A2(new_n729), .A3(new_n726), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n728), .A2(KEYINPUT45), .A3(new_n730), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n511), .A2(KEYINPUT103), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT103), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n736), .B(new_n504), .C1(new_n509), .C2(new_n510), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n500), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT104), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT104), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n500), .A2(new_n735), .A3(new_n740), .A4(new_n737), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n600), .A2(KEYINPUT44), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n739), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT44), .B1(new_n512), .B2(new_n600), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n722), .A2(new_n562), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(G29gat), .B1(new_n747), .B2(new_n453), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n734), .A3(new_n748), .ZN(G1328gat));
  OAI21_X1  g548(.A(G36gat), .B1(new_n747), .B2(new_n452), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n452), .A2(G36gat), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n725), .A2(KEYINPUT46), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT46), .B1(new_n725), .B2(new_n751), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n750), .B1(new_n752), .B2(new_n753), .ZN(G1329gat));
  INV_X1    g553(.A(new_n489), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n565), .A2(new_n755), .A3(new_n723), .ZN(new_n756));
  INV_X1    g555(.A(new_n524), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n756), .A2(new_n757), .B1(KEYINPUT105), .B2(KEYINPUT47), .ZN(new_n758));
  INV_X1    g557(.A(new_n499), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n745), .A2(new_n759), .A3(new_n524), .A4(new_n746), .ZN(new_n760));
  OR2_X1    g559(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n758), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n758), .B2(new_n760), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(G1330gat));
  NOR3_X1   g563(.A1(new_n747), .A2(new_n520), .A3(new_n272), .ZN(new_n765));
  AOI21_X1  g564(.A(G50gat), .B1(new_n725), .B2(new_n455), .ZN(new_n766));
  OR3_X1    g565(.A1(new_n765), .A2(new_n766), .A3(KEYINPUT48), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT48), .B1(new_n765), .B2(new_n766), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(G1331gat));
  INV_X1    g568(.A(new_n691), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n664), .A2(new_n561), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n739), .A2(new_n741), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n453), .ZN(new_n773));
  XOR2_X1   g572(.A(KEYINPUT106), .B(G57gat), .Z(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1332gat));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n772), .A2(new_n776), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n452), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT108), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n782), .B(new_n784), .ZN(G1333gat));
  OAI21_X1  g584(.A(G71gat), .B1(new_n779), .B2(new_n499), .ZN(new_n786));
  OR3_X1    g585(.A1(new_n772), .A2(G71gat), .A3(new_n489), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n786), .A2(KEYINPUT50), .A3(new_n787), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(G1334gat));
  NAND2_X1  g591(.A1(new_n780), .A2(new_n455), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(G78gat), .ZN(G1335gat));
  INV_X1    g593(.A(G85gat), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n662), .A2(new_n561), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n691), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n797), .B1(new_n743), .B2(new_n744), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n795), .B1(new_n798), .B2(new_n566), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n662), .A2(new_n561), .A3(new_n600), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n738), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT51), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n738), .A2(new_n803), .A3(new_n800), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NOR4_X1   g604(.A1(new_n805), .A2(G85gat), .A3(new_n453), .A4(new_n770), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n799), .A2(new_n806), .ZN(G1336gat));
  INV_X1    g606(.A(G92gat), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n798), .B2(new_n704), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n803), .A2(KEYINPUT110), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n801), .B(new_n810), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n770), .A2(G92gat), .A3(new_n452), .ZN(new_n812));
  XOR2_X1   g611(.A(new_n812), .B(KEYINPUT109), .Z(new_n813));
  NOR2_X1   g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT52), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n798), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT111), .B1(new_n816), .B2(new_n452), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n798), .A2(new_n818), .A3(new_n704), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n808), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n821));
  INV_X1    g620(.A(new_n812), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n821), .B1(new_n805), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n815), .B1(new_n820), .B2(new_n823), .ZN(G1337gat));
  OR4_X1    g623(.A1(G99gat), .A2(new_n805), .A3(new_n489), .A4(new_n770), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n816), .A2(new_n499), .ZN(new_n826));
  INV_X1    g625(.A(G99gat), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT112), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n825), .B(new_n830), .C1(new_n827), .C2(new_n826), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(G1338gat));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n834));
  INV_X1    g633(.A(new_n797), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n745), .A2(new_n455), .A3(new_n835), .ZN(new_n836));
  XNOR2_X1  g635(.A(KEYINPUT113), .B(G106gat), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n272), .A2(G106gat), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n691), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n811), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n834), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n837), .B1(new_n798), .B2(new_n455), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n802), .A2(new_n691), .A3(new_n804), .A4(new_n840), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n834), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n833), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n839), .A2(new_n834), .A3(new_n845), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n811), .A2(new_n841), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT53), .B1(new_n844), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n851), .A3(KEYINPUT114), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n848), .A2(new_n852), .ZN(G1339gat));
  NOR2_X1   g652(.A1(new_n704), .A2(new_n453), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n662), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n679), .A2(new_n858), .A3(new_n680), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n677), .B1(new_n670), .B2(new_n672), .ZN(new_n860));
  INV_X1    g659(.A(new_n680), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT54), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI211_X1 g661(.A(new_n680), .B(new_n677), .C1(new_n670), .C2(new_n672), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n859), .B(new_n687), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT55), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n857), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n860), .A2(new_n861), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n681), .A2(KEYINPUT54), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n860), .A2(new_n861), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n689), .B1(new_n869), .B2(new_n858), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n868), .A2(new_n870), .A3(KEYINPUT115), .A4(KEYINPUT55), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n690), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n873), .B1(new_n865), .B2(new_n864), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n561), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n550), .A2(new_n547), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n540), .A2(new_n514), .A3(new_n542), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n556), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n560), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n691), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n599), .B1(new_n875), .B2(new_n880), .ZN(new_n881));
  AND4_X1   g680(.A1(new_n599), .A2(new_n872), .A3(new_n874), .A4(new_n879), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n856), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n657), .A2(new_n663), .A3(new_n562), .A4(new_n770), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n855), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n489), .A2(new_n455), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT116), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(G113gat), .B1(new_n889), .B2(new_n562), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n502), .A2(new_n494), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n885), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n348), .A3(new_n561), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n890), .A2(new_n894), .ZN(G1340gat));
  AOI21_X1  g694(.A(G120gat), .B1(new_n893), .B2(new_n691), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n770), .A2(new_n345), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n888), .B2(new_n897), .ZN(G1341gat));
  OAI21_X1  g697(.A(G127gat), .B1(new_n889), .B2(new_n856), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n893), .A2(new_n340), .A3(new_n662), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(G1342gat));
  OAI21_X1  g700(.A(G134gat), .B1(new_n889), .B2(new_n600), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n453), .B1(new_n883), .B2(new_n884), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n599), .A2(new_n452), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT117), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  AND4_X1   g705(.A1(new_n338), .A2(new_n903), .A3(new_n892), .A4(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT56), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT118), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n902), .B(new_n910), .C1(new_n908), .C2(new_n907), .ZN(G1343gat));
  NOR2_X1   g710(.A1(new_n759), .A2(new_n272), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n885), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n562), .A2(G141gat), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n759), .A2(new_n855), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n455), .A2(KEYINPUT57), .ZN(new_n917));
  AND4_X1   g716(.A1(new_n562), .A2(new_n657), .A3(new_n663), .A4(new_n770), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n883), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g719(.A(KEYINPUT119), .B(new_n856), .C1(new_n881), .C2(new_n882), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n883), .A2(new_n884), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT57), .B1(new_n923), .B2(new_n455), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n561), .B(new_n916), .C1(new_n922), .C2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n915), .B1(new_n925), .B2(G141gat), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT58), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n925), .A2(G141gat), .ZN(new_n930));
  INV_X1    g729(.A(new_n915), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n929), .B1(new_n932), .B2(KEYINPUT58), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n926), .A2(KEYINPUT120), .A3(new_n927), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n928), .B1(new_n933), .B2(new_n934), .ZN(G1344gat));
  NAND2_X1  g734(.A1(new_n903), .A2(new_n912), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n937), .A2(new_n215), .A3(new_n452), .A4(new_n691), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n922), .A2(new_n924), .ZN(new_n939));
  INV_X1    g738(.A(new_n916), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI211_X1 g740(.A(KEYINPUT59), .B(new_n215), .C1(new_n941), .C2(new_n691), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT59), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT57), .ZN(new_n944));
  AOI211_X1 g743(.A(new_n944), .B(new_n272), .C1(new_n883), .C2(new_n884), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n924), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n946), .A2(new_n691), .A3(new_n916), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n943), .B1(new_n947), .B2(G148gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n938), .B1(new_n942), .B2(new_n948), .ZN(G1345gat));
  NAND3_X1  g748(.A1(new_n913), .A2(new_n210), .A3(new_n662), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n941), .A2(new_n662), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n950), .B1(new_n952), .B2(new_n210), .ZN(G1346gat));
  NAND3_X1  g752(.A1(new_n937), .A2(new_n211), .A3(new_n906), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n941), .A2(new_n599), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n954), .B1(new_n956), .B2(new_n211), .ZN(G1347gat));
  NOR2_X1   g756(.A1(new_n566), .A2(new_n452), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n923), .A2(new_n886), .A3(new_n958), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n959), .A2(new_n285), .A3(new_n562), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n566), .B1(new_n883), .B2(new_n884), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n961), .A2(new_n704), .A3(new_n892), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(new_n561), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n960), .B1(new_n963), .B2(new_n285), .ZN(G1348gat));
  NAND3_X1  g763(.A1(new_n962), .A2(new_n286), .A3(new_n691), .ZN(new_n965));
  OAI21_X1  g764(.A(G176gat), .B1(new_n959), .B2(new_n770), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(G1349gat));
  NAND3_X1  g766(.A1(new_n962), .A2(new_n312), .A3(new_n662), .ZN(new_n968));
  OAI21_X1  g767(.A(G183gat), .B1(new_n959), .B2(new_n856), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT60), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n971), .A2(KEYINPUT121), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n970), .B(new_n972), .ZN(G1350gat));
  NAND3_X1  g772(.A1(new_n962), .A2(new_n288), .A3(new_n599), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT122), .ZN(new_n975));
  OAI21_X1  g774(.A(G190gat), .B1(new_n959), .B2(new_n600), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT61), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(G1351gat));
  AND2_X1   g777(.A1(new_n499), .A2(new_n958), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n946), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(new_n561), .ZN(new_n981));
  XNOR2_X1  g780(.A(KEYINPUT124), .B(G197gat), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n759), .A2(new_n452), .A3(new_n272), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n984), .A2(KEYINPUT123), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(KEYINPUT123), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n985), .A2(new_n961), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n562), .A2(new_n982), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n983), .A2(new_n989), .ZN(G1352gat));
  NAND3_X1  g789(.A1(new_n987), .A2(new_n229), .A3(new_n691), .ZN(new_n991));
  XOR2_X1   g790(.A(new_n991), .B(KEYINPUT62), .Z(new_n992));
  NAND3_X1  g791(.A1(new_n946), .A2(new_n691), .A3(new_n979), .ZN(new_n993));
  INV_X1    g792(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n992), .B1(new_n229), .B2(new_n994), .ZN(G1353gat));
  OAI211_X1 g794(.A(new_n662), .B(new_n979), .C1(new_n924), .C2(new_n945), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(G211gat), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT63), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(KEYINPUT126), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT125), .ZN(new_n1001));
  NAND4_X1  g800(.A1(new_n996), .A2(new_n1001), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n1002));
  OAI21_X1  g801(.A(KEYINPUT125), .B1(new_n997), .B2(new_n998), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT126), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n997), .A2(new_n1004), .A3(new_n998), .ZN(new_n1005));
  NAND4_X1  g804(.A1(new_n1000), .A2(new_n1002), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1006));
  INV_X1    g805(.A(G211gat), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n987), .A2(new_n1007), .A3(new_n662), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1006), .A2(new_n1008), .ZN(G1354gat));
  INV_X1    g808(.A(G218gat), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n987), .A2(new_n1010), .A3(new_n599), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n980), .A2(new_n599), .ZN(new_n1012));
  INV_X1    g811(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1011), .B1(new_n1013), .B2(new_n1010), .ZN(G1355gat));
endmodule


