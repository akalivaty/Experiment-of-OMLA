//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n202), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  XOR2_X1   g0014(.A(KEYINPUT64), .B(G244), .Z(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G107), .A2(G264), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n205), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n208), .B(new_n214), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0025(.A(G226), .B(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT66), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G68), .B(G77), .ZN(new_n236));
  INV_X1    g0036(.A(G58), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT67), .B(G50), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  AND2_X1   g0044(.A1(G33), .A2(G41), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n245), .A2(new_n211), .ZN(new_n246));
  INV_X1    g0046(.A(G274), .ZN(new_n247));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n248), .B1(G41), .B2(G45), .ZN(new_n249));
  NOR3_X1   g0049(.A1(new_n246), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n249), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n250), .B1(G238), .B2(new_n252), .ZN(new_n253));
  AND2_X1   g0053(.A1(G1), .A2(G13), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  AND3_X1   g0055(.A1(new_n254), .A2(KEYINPUT68), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT68), .B1(new_n254), .B2(new_n255), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n260), .A2(new_n262), .A3(G226), .A4(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G97), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n264), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n260), .A2(new_n262), .ZN(new_n267));
  INV_X1    g0067(.A(G232), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n267), .A2(new_n268), .A3(new_n263), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n258), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT13), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n253), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n271), .B1(new_n253), .B2(new_n270), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G169), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT14), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT14), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n277), .B(G169), .C1(new_n272), .C2(new_n273), .ZN(new_n278));
  AOI21_X1  g0078(.A(KEYINPUT76), .B1(new_n274), .B2(G179), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT76), .ZN(new_n280));
  INV_X1    g0080(.A(G179), .ZN(new_n281));
  NOR4_X1   g0081(.A1(new_n272), .A2(new_n273), .A3(new_n280), .A4(new_n281), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n276), .B(new_n278), .C1(new_n279), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n248), .A2(G13), .A3(G20), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n284), .A2(G68), .B1(KEYINPUT75), .B2(KEYINPUT12), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT75), .A2(KEYINPUT12), .ZN(new_n286));
  OR2_X1    g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n286), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n211), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n284), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n248), .A2(G20), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G68), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n212), .A2(G33), .ZN(new_n296));
  OAI22_X1  g0096(.A1(new_n296), .A2(new_n216), .B1(new_n212), .B2(G68), .ZN(new_n297));
  INV_X1    g0097(.A(G50), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G20), .A2(G33), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n297), .A2(KEYINPUT74), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n297), .A2(KEYINPUT74), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n291), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT11), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n289), .B1(new_n293), .B2(new_n295), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n303), .A2(new_n304), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n283), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n274), .A2(G190), .ZN(new_n311));
  OAI21_X1  g0111(.A(G200), .B1(new_n272), .B2(new_n273), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(new_n307), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n294), .A2(G50), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n293), .A2(new_n316), .B1(G50), .B2(new_n284), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n317), .B(KEYINPUT70), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n212), .B1(new_n201), .B2(new_n298), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n319), .B(KEYINPUT69), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT8), .B(G58), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n296), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n322), .A2(new_n323), .B1(G150), .B2(new_n299), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n292), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n318), .A2(new_n325), .ZN(new_n326));
  OR2_X1    g0126(.A1(new_n326), .A2(KEYINPUT9), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT3), .B(G33), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(G222), .A3(new_n263), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(G1698), .ZN(new_n330));
  INV_X1    g0130(.A(G223), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n329), .B1(new_n216), .B2(new_n328), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n258), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n250), .B1(G226), .B2(new_n252), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(G190), .B1(KEYINPUT73), .B2(KEYINPUT10), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(G200), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n326), .A2(KEYINPUT9), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n327), .A2(new_n337), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT73), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT10), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n340), .B(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n326), .B1(new_n275), .B2(new_n335), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(G179), .B2(new_n335), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n322), .A2(new_n299), .B1(G20), .B2(G77), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT15), .B(G87), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n323), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n292), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n294), .A2(G77), .ZN(new_n352));
  OAI22_X1  g0152(.A1(new_n293), .A2(new_n352), .B1(G77), .B2(new_n284), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT72), .ZN(new_n355));
  INV_X1    g0155(.A(G238), .ZN(new_n356));
  XOR2_X1   g0156(.A(KEYINPUT71), .B(G107), .Z(new_n357));
  OAI22_X1  g0157(.A1(new_n330), .A2(new_n356), .B1(new_n357), .B2(new_n328), .ZN(new_n358));
  NOR3_X1   g0158(.A1(new_n267), .A2(new_n268), .A3(G1698), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n258), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n250), .ZN(new_n361));
  INV_X1    g0161(.A(new_n252), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n360), .B(new_n361), .C1(new_n215), .C2(new_n362), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n363), .A2(G179), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n275), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n355), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n363), .A2(G200), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n355), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n367), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n315), .A2(new_n344), .A3(new_n346), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n322), .A2(new_n294), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n374), .A2(new_n293), .B1(new_n284), .B2(new_n322), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT16), .ZN(new_n376));
  INV_X1    g0176(.A(G68), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n237), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(G20), .B1(new_n378), .B2(new_n201), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n299), .A2(G159), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT7), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n328), .B2(G20), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n267), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n377), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT77), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n382), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI211_X1 g0188(.A(KEYINPUT77), .B(new_n377), .C1(new_n384), .C2(new_n385), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n376), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n386), .A2(new_n381), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n292), .B1(new_n391), .B2(KEYINPUT16), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n375), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G200), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n256), .A2(new_n257), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n260), .A2(new_n262), .A3(G226), .A4(G1698), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT78), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT78), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n328), .A2(new_n398), .A3(G226), .A4(G1698), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n260), .A2(new_n262), .A3(G223), .A4(new_n263), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G87), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n395), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n361), .B1(new_n362), .B2(new_n268), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n394), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n250), .B1(G232), .B2(new_n252), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n403), .B1(new_n399), .B2(new_n397), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n408), .B(new_n369), .C1(new_n409), .C2(new_n395), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n393), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n412), .B(KEYINPUT17), .ZN(new_n413));
  INV_X1    g0213(.A(new_n375), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT7), .B1(new_n267), .B2(new_n212), .ZN(new_n415));
  AOI211_X1 g0215(.A(new_n383), .B(G20), .C1(new_n260), .C2(new_n262), .ZN(new_n416));
  OAI21_X1  g0216(.A(G68), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n381), .B1(new_n417), .B2(KEYINPUT77), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n386), .A2(new_n387), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT16), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n417), .A2(KEYINPUT16), .A3(new_n382), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n291), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n414), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(G169), .B1(new_n405), .B2(new_n406), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n408), .B(G179), .C1(new_n409), .C2(new_n395), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT18), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n424), .A2(new_n425), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT18), .B1(new_n393), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT79), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n431), .B1(new_n428), .B2(new_n430), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n413), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n373), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n260), .A2(new_n262), .A3(G257), .A4(G1698), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n260), .A2(new_n262), .A3(G250), .A4(new_n263), .ZN(new_n437));
  INV_X1    g0237(.A(G294), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n436), .B(new_n437), .C1(new_n259), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n258), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n248), .A2(G45), .ZN(new_n441));
  OR2_X1    g0241(.A1(KEYINPUT5), .A2(G41), .ZN(new_n442));
  NAND2_X1  g0242(.A1(KEYINPUT5), .A2(G41), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n247), .B1(new_n254), .B2(new_n255), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n444), .A2(new_n246), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G264), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n440), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(KEYINPUT84), .A3(G169), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n439), .A2(new_n258), .B1(new_n447), .B2(G264), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(G179), .A3(new_n446), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT84), .B1(new_n449), .B2(G169), .ZN(new_n454));
  INV_X1    g0254(.A(G107), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G20), .ZN(new_n456));
  INV_X1    g0256(.A(G116), .ZN(new_n457));
  OAI22_X1  g0257(.A1(KEYINPUT23), .A2(new_n456), .B1(new_n296), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n357), .A2(G20), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n458), .B1(new_n459), .B2(KEYINPUT23), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n260), .A2(new_n262), .A3(new_n212), .A4(G87), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT22), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT22), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n328), .A2(new_n463), .A3(new_n212), .A4(G87), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT24), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT24), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n460), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n292), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G13), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G1), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(G20), .A3(new_n455), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n473), .B(KEYINPUT25), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n248), .A2(G33), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n284), .A2(new_n475), .A3(new_n211), .A4(new_n290), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(new_n455), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n453), .A2(new_n454), .B1(new_n470), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n469), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n468), .B1(new_n460), .B2(new_n465), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n291), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n451), .A2(G190), .A3(new_n446), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n449), .A2(G200), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n483), .A2(new_n478), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n447), .A2(G270), .B1(new_n445), .B2(new_n444), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n260), .A2(new_n262), .A3(G264), .A4(G1698), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n260), .A2(new_n262), .A3(G257), .A4(new_n263), .ZN(new_n490));
  XOR2_X1   g0290(.A(KEYINPUT81), .B(G303), .Z(new_n491));
  OAI211_X1 g0291(.A(new_n489), .B(new_n490), .C1(new_n491), .C2(new_n328), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n258), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n476), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G116), .ZN(new_n496));
  INV_X1    g0296(.A(new_n284), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n457), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n290), .A2(new_n211), .B1(G20), .B2(new_n457), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G283), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n500), .B(new_n212), .C1(G33), .C2(new_n265), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n499), .A2(KEYINPUT20), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT20), .B1(new_n499), .B2(new_n501), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n496), .B(new_n498), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n494), .A2(G169), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT82), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(KEYINPUT21), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(G45), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(G1), .ZN(new_n510));
  INV_X1    g0310(.A(new_n443), .ZN(new_n511));
  NOR2_X1   g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n254), .A2(new_n255), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(G270), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n446), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n517), .B1(new_n258), .B2(new_n492), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(G179), .A3(new_n504), .ZN(new_n519));
  INV_X1    g0319(.A(new_n507), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n494), .A2(G169), .A3(new_n520), .A4(new_n504), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n508), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n518), .A2(G190), .ZN(new_n523));
  INV_X1    g0323(.A(new_n504), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n494), .A2(G200), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT83), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT83), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n523), .A2(new_n525), .A3(new_n528), .A4(new_n524), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n522), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n441), .A2(G250), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n514), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n445), .A2(new_n510), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n260), .A2(new_n262), .A3(G244), .A4(G1698), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n260), .A2(new_n262), .A3(G238), .A4(new_n263), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G116), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n258), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G200), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n349), .A2(new_n284), .ZN(new_n542));
  INV_X1    g0342(.A(G87), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n476), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n212), .ZN(new_n546));
  XNOR2_X1  g0346(.A(KEYINPUT71), .B(G107), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n543), .A2(new_n265), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n328), .A2(new_n212), .A3(G68), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT19), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n296), .B2(new_n265), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  AOI211_X1 g0353(.A(new_n542), .B(new_n544), .C1(new_n553), .C2(new_n291), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n534), .A2(new_n539), .A3(G190), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n541), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n540), .A2(new_n275), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n553), .A2(new_n291), .ZN(new_n558));
  INV_X1    g0358(.A(new_n542), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n495), .A2(new_n349), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n534), .A2(new_n539), .A3(new_n281), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n557), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n284), .A2(G97), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n495), .B2(G97), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n547), .B1(new_n415), .B2(new_n416), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT6), .ZN(new_n568));
  AND2_X1   g0368(.A1(G97), .A2(G107), .ZN(new_n569));
  NOR2_X1   g0369(.A1(G97), .A2(G107), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT80), .ZN(new_n572));
  NAND2_X1  g0372(.A1(KEYINPUT6), .A2(G97), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n572), .B1(new_n573), .B2(G107), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n455), .A2(KEYINPUT80), .A3(KEYINPUT6), .A4(G97), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n571), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(G20), .B1(G77), .B2(new_n299), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n567), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n566), .B1(new_n578), .B2(new_n292), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n260), .A2(new_n262), .A3(G250), .A4(G1698), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n260), .A2(new_n262), .A3(G244), .A4(new_n263), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT4), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n500), .B(new_n580), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n581), .A2(new_n582), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n258), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G257), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n446), .B1(new_n515), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n275), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n581), .A2(new_n582), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n328), .A2(KEYINPUT4), .A3(G244), .A4(new_n263), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(new_n500), .A4(new_n580), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n587), .B1(new_n258), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n281), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n579), .A2(new_n590), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n292), .B1(new_n567), .B2(new_n577), .ZN(new_n597));
  INV_X1    g0397(.A(new_n566), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n589), .A2(G200), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n594), .A2(G190), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n564), .A2(new_n596), .A3(new_n602), .ZN(new_n603));
  AND4_X1   g0403(.A1(new_n435), .A2(new_n487), .A3(new_n530), .A4(new_n603), .ZN(G372));
  INV_X1    g0404(.A(new_n563), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n564), .A2(new_n486), .A3(new_n596), .A4(new_n602), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n519), .A2(new_n521), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n275), .B1(new_n488), .B2(new_n493), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n520), .B1(new_n609), .B2(new_n504), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n480), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n605), .B1(new_n607), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT85), .ZN(new_n614));
  OAI22_X1  g0414(.A1(G179), .A2(new_n589), .B1(new_n597), .B2(new_n598), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n594), .A2(G169), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n579), .A2(KEYINPUT85), .A3(new_n590), .A4(new_n595), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(new_n564), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT26), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(KEYINPUT86), .A3(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n615), .A2(new_n616), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n564), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g0423(.A(KEYINPUT87), .B(KEYINPUT26), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT88), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT88), .ZN(new_n626));
  INV_X1    g0426(.A(new_n624), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n564), .A2(new_n622), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n621), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT86), .B1(new_n619), .B2(new_n620), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n613), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n435), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g0432(.A(new_n632), .B(KEYINPUT89), .Z(new_n633));
  INV_X1    g0433(.A(new_n346), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n393), .A2(new_n429), .A3(KEYINPUT18), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n427), .B1(new_n423), .B2(new_n426), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n310), .A2(new_n367), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n413), .A2(new_n313), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n634), .B1(new_n640), .B2(new_n344), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n633), .A2(new_n641), .ZN(G369));
  NAND2_X1  g0442(.A1(new_n472), .A2(new_n212), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(G213), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n504), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n530), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n611), .B2(new_n649), .ZN(new_n651));
  XNOR2_X1  g0451(.A(KEYINPUT90), .B(G330), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n483), .A2(new_n478), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n648), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n487), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n648), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n658), .B1(new_n480), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n454), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(new_n452), .A3(new_n450), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n663), .A2(new_n656), .A3(new_n659), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n611), .A2(new_n648), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n487), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n661), .A2(new_n664), .A3(new_n666), .ZN(G399));
  INV_X1    g0467(.A(new_n206), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(G41), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n547), .A2(G116), .A3(new_n548), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G1), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n209), .B2(new_n670), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT28), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n556), .A2(new_n563), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n624), .B1(new_n596), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT92), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n617), .A2(new_n564), .A3(KEYINPUT26), .A4(new_n618), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT92), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n679), .B(new_n624), .C1(new_n596), .C2(new_n675), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT93), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n522), .B1(new_n656), .B2(new_n663), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n682), .B1(new_n683), .B2(new_n606), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n603), .A2(new_n612), .A3(KEYINPUT93), .A4(new_n486), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n681), .A2(new_n684), .A3(new_n685), .A4(new_n563), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n686), .A2(KEYINPUT29), .A3(new_n659), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n619), .A2(new_n620), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT86), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n690), .A2(new_n621), .A3(new_n625), .A4(new_n628), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n648), .B1(new_n691), .B2(new_n613), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n687), .B1(new_n692), .B2(KEYINPUT29), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n589), .A2(new_n449), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n494), .A2(new_n281), .A3(new_n540), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n532), .A2(new_n533), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n258), .B2(new_n538), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n518), .A2(G179), .A3(new_n451), .A4(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT91), .B1(new_n699), .B2(new_n589), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n696), .B1(new_n700), .B2(KEYINPUT30), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  OAI211_X1 g0502(.A(KEYINPUT91), .B(new_n702), .C1(new_n699), .C2(new_n589), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n659), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT31), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n487), .A2(new_n603), .A3(new_n530), .A4(new_n659), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n704), .A2(KEYINPUT31), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n653), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n693), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n674), .B1(new_n711), .B2(G1), .ZN(G364));
  NOR2_X1   g0512(.A1(new_n471), .A2(G20), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n248), .B1(new_n713), .B2(G45), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n669), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n655), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n653), .B2(new_n651), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n328), .A2(new_n206), .ZN(new_n719));
  INV_X1    g0519(.A(G355), .ZN(new_n720));
  OAI22_X1  g0520(.A1(new_n719), .A2(new_n720), .B1(G116), .B2(new_n206), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n267), .A2(new_n206), .ZN(new_n722));
  XOR2_X1   g0522(.A(new_n722), .B(KEYINPUT94), .Z(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n724), .B1(new_n509), .B2(new_n210), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n240), .A2(G45), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n721), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G13), .A2(G33), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n211), .B1(G20), .B2(new_n275), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n716), .B1(new_n727), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n212), .A2(new_n281), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G200), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT95), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G190), .ZN(new_n738));
  XNOR2_X1  g0538(.A(KEYINPUT33), .B(G317), .ZN(new_n739));
  INV_X1    g0539(.A(new_n735), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n740), .A2(new_n369), .A3(G200), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n738), .A2(new_n739), .B1(G322), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT97), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n740), .A2(G190), .A3(G200), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n328), .B1(new_n744), .B2(G311), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n212), .A2(G179), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(G190), .A3(G200), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G303), .ZN(new_n749));
  INV_X1    g0549(.A(G283), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n746), .A2(new_n369), .A3(G200), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n745), .B(new_n749), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n281), .A2(new_n394), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT96), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n754), .A2(G20), .A3(new_n369), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n752), .B1(G329), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n737), .A2(new_n369), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n754), .A2(G190), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n758), .A2(G326), .B1(new_n760), .B2(G294), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n743), .A2(new_n757), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n756), .A2(G159), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(KEYINPUT32), .ZN(new_n764));
  INV_X1    g0564(.A(new_n744), .ZN(new_n765));
  INV_X1    g0565(.A(new_n741), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n328), .B1(new_n765), .B2(new_n216), .C1(new_n237), .C2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n747), .A2(new_n543), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n751), .A2(new_n455), .ZN(new_n769));
  NOR4_X1   g0569(.A1(new_n764), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n763), .A2(KEYINPUT32), .B1(G97), .B2(new_n760), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G50), .A2(new_n758), .B1(new_n738), .B2(G68), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n762), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n734), .B1(new_n774), .B2(new_n731), .ZN(new_n775));
  INV_X1    g0575(.A(new_n730), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n775), .B1(new_n651), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n718), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(G396));
  NAND2_X1  g0579(.A1(new_n367), .A2(new_n659), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n371), .A2(new_n368), .B1(new_n355), .B2(new_n648), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n780), .B1(new_n781), .B2(new_n367), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n692), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT100), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n372), .A2(new_n659), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n631), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n716), .B1(new_n789), .B2(new_n709), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(new_n709), .B2(new_n789), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n543), .A2(new_n751), .B1(new_n747), .B2(new_n455), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n267), .B1(new_n765), .B2(new_n457), .C1(new_n438), .C2(new_n766), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n792), .B(new_n793), .C1(G311), .C2(new_n756), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n758), .A2(G303), .B1(new_n760), .B2(G97), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n738), .A2(KEYINPUT98), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n738), .A2(KEYINPUT98), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n794), .B(new_n795), .C1(new_n799), .C2(new_n750), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G143), .A2(new_n741), .B1(new_n744), .B2(G159), .ZN(new_n801));
  INV_X1    g0601(.A(new_n738), .ZN(new_n802));
  INV_X1    g0602(.A(G150), .ZN(new_n803));
  INV_X1    g0603(.A(G137), .ZN(new_n804));
  INV_X1    g0604(.A(new_n758), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n801), .B1(new_n802), .B2(new_n803), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT34), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G132), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n328), .B1(new_n755), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(G58), .B2(new_n760), .ZN(new_n811));
  INV_X1    g0611(.A(new_n751), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G68), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n298), .B2(new_n747), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT99), .Z(new_n815));
  NAND3_X1  g0615(.A1(new_n808), .A2(new_n811), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n806), .A2(new_n807), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n800), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n731), .ZN(new_n819));
  INV_X1    g0619(.A(new_n716), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n731), .A2(new_n728), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n820), .B1(new_n216), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n819), .B(new_n822), .C1(new_n783), .C2(new_n729), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n791), .A2(new_n823), .ZN(G384));
  OR2_X1    g0624(.A1(new_n576), .A2(KEYINPUT35), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n576), .A2(KEYINPUT35), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n825), .A2(G116), .A3(new_n213), .A4(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT36), .Z(new_n828));
  OR3_X1    g0628(.A1(new_n209), .A2(new_n216), .A3(new_n378), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n298), .A2(G68), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n248), .B(G13), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT39), .ZN(new_n833));
  INV_X1    g0633(.A(new_n646), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n376), .B1(new_n386), .B2(new_n381), .ZN(new_n835));
  AND3_X1   g0635(.A1(new_n835), .A2(KEYINPUT101), .A3(new_n291), .ZN(new_n836));
  AOI21_X1  g0636(.A(KEYINPUT101), .B1(new_n835), .B2(new_n291), .ZN(new_n837));
  INV_X1    g0637(.A(new_n421), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n834), .B1(new_n839), .B2(new_n375), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT79), .B1(new_n635), .B2(new_n636), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n840), .B1(new_n843), .B2(new_n413), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n390), .A2(new_n392), .ZN(new_n845));
  AND3_X1   g0645(.A1(new_n845), .A2(new_n411), .A3(new_n414), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n845), .A2(new_n414), .B1(new_n424), .B2(new_n425), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT102), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n423), .A2(new_n834), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n848), .A2(new_n849), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n423), .A2(new_n426), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n853), .A2(new_n851), .A3(new_n850), .A4(new_n412), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT102), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n426), .B1(new_n839), .B2(new_n375), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n840), .A2(new_n856), .A3(new_n412), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n852), .A2(new_n855), .B1(KEYINPUT37), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT38), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n844), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n848), .A2(new_n851), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n854), .A2(KEYINPUT102), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n854), .A2(KEYINPUT102), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n851), .B1(new_n413), .B2(new_n637), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT38), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n833), .B1(new_n860), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n309), .A2(new_n648), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n859), .B1(new_n844), .B2(new_n858), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n857), .A2(KEYINPUT37), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n863), .B2(new_n864), .ZN(new_n873));
  INV_X1    g0673(.A(new_n840), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n434), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n873), .A2(new_n875), .A3(KEYINPUT38), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n871), .A2(new_n876), .A3(KEYINPUT39), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n869), .A2(new_n870), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n637), .A2(new_n834), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n308), .A2(new_n648), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n309), .A2(new_n313), .A3(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n308), .B(new_n648), .C1(new_n283), .C2(new_n314), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n788), .B2(new_n780), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n871), .A2(new_n876), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n879), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n878), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n435), .B(new_n687), .C1(KEYINPUT29), .C2(new_n692), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n641), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n887), .B(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT40), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT31), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n704), .B2(KEYINPUT103), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT103), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n894), .B(new_n659), .C1(new_n701), .C2(new_n703), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n705), .B(new_n706), .C1(new_n893), .C2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n782), .B1(new_n881), .B2(new_n882), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n885), .A2(new_n891), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n896), .A2(new_n897), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n852), .A2(new_n855), .B1(new_n861), .B2(KEYINPUT37), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n859), .B1(new_n901), .B2(new_n866), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n900), .B1(new_n876), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n899), .B1(new_n891), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n435), .A2(new_n896), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n904), .B(new_n905), .Z(new_n906));
  OAI21_X1  g0706(.A(new_n890), .B1(new_n906), .B2(new_n652), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n248), .B2(new_n713), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n906), .A2(new_n890), .A3(new_n652), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n832), .B1(new_n908), .B2(new_n909), .ZN(G367));
  NAND2_X1  g0710(.A1(new_n666), .A2(new_n664), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n596), .B(new_n602), .C1(new_n599), .C2(new_n659), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n622), .A2(new_n648), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT45), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n911), .A2(new_n915), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT105), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT44), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n919), .B2(new_n920), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n917), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(new_n661), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n666), .B1(new_n660), .B2(new_n665), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(new_n654), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n710), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n669), .B(KEYINPUT41), .Z(new_n930));
  OAI21_X1  g0730(.A(new_n714), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n659), .A2(new_n554), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n605), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n675), .B2(new_n932), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n914), .A2(new_n487), .A3(new_n665), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT42), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n596), .B1(new_n912), .B2(new_n480), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n659), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n936), .A2(KEYINPUT42), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n935), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT104), .Z(new_n944));
  XNOR2_X1  g0744(.A(new_n942), .B(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n661), .A2(new_n915), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n931), .A2(new_n948), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n723), .A2(new_n234), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n732), .B1(new_n206), .B2(new_n348), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n716), .B1(new_n950), .B2(new_n951), .C1(new_n934), .C2(new_n776), .ZN(new_n952));
  INV_X1    g0752(.A(new_n760), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(new_n377), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n328), .B1(new_n237), .B2(new_n747), .C1(new_n766), .C2(new_n803), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(G77), .B2(new_n812), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n804), .B2(new_n755), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n954), .B(new_n957), .C1(G143), .C2(new_n758), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n798), .A2(G159), .B1(G50), .B2(new_n744), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n959), .A2(KEYINPUT107), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(KEYINPUT107), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT108), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n747), .A2(new_n457), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(KEYINPUT46), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(KEYINPUT46), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n965), .B(new_n966), .C1(new_n799), .C2(new_n438), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n968), .A2(KEYINPUT106), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(KEYINPUT106), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n267), .B1(new_n765), .B2(new_n750), .C1(new_n491), .C2(new_n766), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n756), .A2(G317), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n751), .A2(new_n265), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n758), .A2(G311), .B1(new_n760), .B2(new_n547), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n969), .A2(new_n970), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n963), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT47), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n731), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(new_n979), .B2(new_n980), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n952), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n949), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(KEYINPUT109), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n985), .B1(new_n931), .B2(new_n948), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT109), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(G387));
  OR2_X1    g0793(.A1(new_n660), .A2(new_n776), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n671), .A2(new_n719), .B1(G107), .B2(new_n206), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT110), .Z(new_n996));
  NAND2_X1  g0796(.A1(new_n231), .A2(G45), .ZN(new_n997));
  INV_X1    g0797(.A(new_n671), .ZN(new_n998));
  AOI211_X1 g0798(.A(G45), .B(new_n998), .C1(G68), .C2(G77), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n321), .A2(G50), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT50), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n724), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n996), .B1(new_n997), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n716), .B1(new_n1003), .B2(new_n733), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n328), .B1(new_n765), .B2(new_n377), .C1(new_n298), .C2(new_n766), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n973), .B(new_n1005), .C1(G159), .C2(new_n758), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n747), .A2(new_n216), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(KEYINPUT111), .B(G150), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1007), .B1(new_n756), .B2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT112), .Z(new_n1010));
  NAND2_X1  g0810(.A1(new_n738), .A2(new_n322), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n760), .A2(new_n349), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1006), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n758), .A2(G322), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n741), .A2(G317), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(new_n491), .C2(new_n765), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n798), .B2(G311), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1017), .A2(KEYINPUT48), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n953), .A2(new_n750), .B1(new_n438), .B2(new_n747), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1017), .A2(KEYINPUT48), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1020), .A2(KEYINPUT49), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n756), .A2(G326), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n328), .B1(new_n812), .B2(G116), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT49), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1013), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1004), .B1(new_n1027), .B2(new_n731), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n928), .A2(new_n715), .B1(new_n994), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n711), .A2(new_n928), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n669), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n711), .A2(new_n928), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(G393));
  NAND2_X1  g0833(.A1(new_n925), .A2(new_n715), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n732), .B1(new_n265), .B2(new_n206), .C1(new_n724), .C2(new_n243), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n716), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n751), .A2(new_n543), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n328), .B1(new_n765), .B2(new_n321), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1037), .B(new_n1038), .C1(G68), .C2(new_n748), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n953), .A2(new_n216), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n756), .A2(G143), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n758), .A2(G150), .B1(G159), .B2(new_n741), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  XOR2_X1   g0845(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n1046));
  OAI22_X1  g0846(.A1(new_n799), .A2(new_n298), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1043), .B(new_n1047), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1049), .A2(KEYINPUT114), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(KEYINPUT114), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n758), .A2(G317), .B1(G311), .B2(new_n741), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT52), .Z(new_n1053));
  NAND2_X1  g0853(.A1(new_n756), .A2(G322), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n328), .B(new_n769), .C1(G294), .C2(new_n744), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n750), .C2(new_n747), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G116), .B2(new_n760), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1053), .B(new_n1057), .C1(new_n491), .C2(new_n799), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1050), .A2(new_n1051), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1036), .B1(new_n1059), .B2(new_n731), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n776), .B2(new_n914), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1034), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(KEYINPUT115), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT115), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1034), .A2(new_n1064), .A3(new_n1061), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1030), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n670), .B1(new_n925), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n1067), .B2(new_n925), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1066), .A2(new_n1069), .ZN(G390));
  NAND3_X1  g0870(.A1(new_n435), .A2(G330), .A3(new_n896), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n888), .A2(new_n641), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n883), .B1(new_n709), .B2(new_n782), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n896), .A2(G330), .A3(new_n897), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n786), .B1(new_n691), .B2(new_n613), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n780), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OR3_X1    g0878(.A1(new_n709), .A2(new_n782), .A3(new_n883), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n896), .A2(G330), .A3(new_n783), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n883), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n781), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n366), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n686), .A2(new_n659), .A3(new_n1083), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1079), .A2(new_n1081), .A3(new_n780), .A4(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1072), .B1(new_n1078), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT116), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1074), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n870), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n883), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n869), .A2(new_n877), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1084), .A2(new_n780), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n1091), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n870), .B1(new_n876), .B2(new_n902), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1088), .B(new_n1089), .C1(new_n1093), .C2(new_n1097), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n871), .A2(new_n876), .A3(KEYINPUT39), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT39), .B1(new_n876), .B2(new_n902), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1099), .A2(new_n1100), .B1(new_n870), .B2(new_n884), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1101), .A2(new_n1102), .A3(new_n1079), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1098), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1088), .B1(new_n1105), .B2(new_n1089), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1087), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1093), .A2(new_n1097), .ZN(new_n1108));
  OAI21_X1  g0908(.A(KEYINPUT116), .B1(new_n1108), .B2(new_n1074), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1109), .A2(new_n1103), .A3(new_n1098), .A4(new_n1086), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1107), .A2(new_n1110), .A3(new_n669), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n728), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n751), .A2(new_n298), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT54), .B(G143), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n328), .B1(new_n765), .B2(new_n1115), .C1(new_n809), .C2(new_n766), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1114), .B(new_n1116), .C1(G128), .C2(new_n758), .ZN(new_n1117));
  INV_X1    g0917(.A(G159), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1117), .B1(new_n1118), .B2(new_n953), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n748), .A2(new_n1008), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n756), .A2(G125), .B1(KEYINPUT53), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(KEYINPUT53), .B2(new_n1120), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n804), .B2(new_n799), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n813), .B1(new_n766), .B2(new_n457), .C1(new_n265), .C2(new_n765), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1125), .B(new_n1040), .C1(G294), .C2(new_n756), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n768), .A2(new_n328), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT117), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G283), .B2(new_n758), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1126), .B(new_n1129), .C1(new_n799), .C2(new_n357), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT118), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n983), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n1132), .B2(new_n1131), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n820), .B1(new_n321), .B2(new_n821), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1112), .A2(new_n715), .B1(new_n1113), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1111), .A2(new_n1137), .ZN(G378));
  NAND3_X1  g0938(.A1(new_n887), .A2(G330), .A3(new_n904), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n876), .A2(new_n902), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n891), .B1(new_n1140), .B2(new_n898), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n896), .A2(new_n891), .A3(new_n897), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n876), .B2(new_n871), .ZN(new_n1143));
  OAI21_X1  g0943(.A(G330), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(new_n878), .A3(new_n886), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n344), .A2(new_n346), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n326), .A2(new_n646), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT120), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1146), .B(new_n1148), .ZN(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1150));
  XNOR2_X1  g0950(.A(new_n1149), .B(new_n1150), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1139), .A2(new_n1145), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1151), .B1(new_n1139), .B2(new_n1145), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n715), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n328), .A2(G41), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n766), .B2(new_n455), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n349), .B2(new_n744), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n237), .B2(new_n751), .C1(new_n216), .C2(new_n747), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n954), .B1(G116), .B2(new_n758), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n265), .B2(new_n802), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1158), .B(new_n1160), .C1(G283), .C2(new_n756), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n298), .B1(G33), .B2(G41), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n1161), .A2(KEYINPUT58), .B1(new_n1155), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT119), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G128), .A2(new_n741), .B1(new_n744), .B2(G137), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n747), .B2(new_n1115), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G125), .B2(new_n758), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n809), .B2(new_n802), .C1(new_n803), .C2(new_n953), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1170));
  AOI211_X1 g0970(.A(G33), .B(G41), .C1(new_n812), .C2(G159), .ZN(new_n1171));
  INV_X1    g0971(.A(G124), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1171), .B1(new_n1172), .B2(new_n755), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n1169), .B2(KEYINPUT59), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1161), .A2(KEYINPUT58), .B1(new_n1170), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1165), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n731), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n820), .B1(new_n298), .B2(new_n821), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n1151), .B2(new_n728), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1154), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1078), .A2(new_n1085), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1072), .B1(new_n1112), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT57), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n669), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1072), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1110), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1139), .A2(new_n1145), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1151), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1139), .A2(new_n1145), .A3(new_n1151), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT57), .B1(new_n1190), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1184), .B1(new_n1188), .B2(new_n1196), .ZN(G375));
  NAND2_X1  g0997(.A1(new_n1185), .A2(new_n715), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1198), .A2(KEYINPUT121), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n820), .B1(new_n377), .B2(new_n821), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n216), .A2(new_n751), .B1(new_n747), .B2(new_n265), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n267), .B1(new_n765), .B2(new_n357), .C1(new_n750), .C2(new_n766), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(G303), .C2(new_n756), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n758), .A2(G294), .B1(new_n760), .B2(new_n349), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n799), .C2(new_n457), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT122), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n237), .A2(new_n751), .B1(new_n747), .B2(new_n1118), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n328), .B1(new_n765), .B2(new_n803), .C1(new_n804), .C2(new_n766), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(G128), .C2(new_n756), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n758), .A2(G132), .B1(new_n760), .B2(G50), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1210), .B(new_n1211), .C1(new_n799), .C2(new_n1115), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1207), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1200), .B1(new_n983), .B2(new_n1214), .C1(new_n1091), .C2(new_n729), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1198), .A2(KEYINPUT121), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1199), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT123), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1217), .B(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1185), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1072), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n930), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1087), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1220), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(G381));
  OR2_X1    g1026(.A1(G393), .A2(G396), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(G390), .A2(G384), .A3(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1225), .A2(new_n992), .A3(new_n1228), .ZN(new_n1229));
  OR3_X1    g1029(.A1(new_n1229), .A2(G378), .A3(G375), .ZN(G407));
  AND2_X1   g1030(.A1(new_n1111), .A2(new_n1137), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n647), .A2(G213), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  OAI211_X1 g1034(.A(G407), .B(G213), .C1(G375), .C2(new_n1234), .ZN(G409));
  NAND2_X1  g1035(.A1(G393), .A2(G396), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(G390), .A2(new_n989), .B1(new_n1227), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT125), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G390), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1066), .A2(new_n1069), .A3(KEYINPUT125), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1237), .B1(new_n1241), .B2(new_n992), .ZN(new_n1242));
  AND2_X1   g1042(.A1(G390), .A2(new_n989), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(G390), .A2(new_n989), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1227), .B(new_n1236), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT61), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(G378), .B(new_n1184), .C1(new_n1188), .C2(new_n1196), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1190), .A2(new_n1195), .A3(new_n1223), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1231), .B1(new_n1250), .B2(new_n1183), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1233), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT60), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1222), .B1(new_n1253), .B2(new_n1086), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1221), .A2(KEYINPUT60), .A3(new_n1072), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n669), .A3(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1216), .A2(new_n1215), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT123), .B1(new_n1258), .B2(new_n1199), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1256), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(new_n791), .A3(new_n823), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1219), .A2(G384), .A3(new_n1256), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT63), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1248), .B1(new_n1252), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT124), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1249), .A2(new_n1251), .A3(KEYINPUT124), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1269), .A2(new_n1232), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1264), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1269), .A2(new_n1232), .A3(new_n1271), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1233), .A2(G2897), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1263), .B(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1266), .B(new_n1273), .C1(new_n1274), .C2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1247), .B1(new_n1277), .B2(new_n1252), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1270), .A2(new_n1252), .A3(KEYINPUT62), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT62), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1272), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT126), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1280), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1272), .A2(KEYINPUT126), .A3(new_n1281), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1279), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1278), .B1(new_n1286), .B2(new_n1246), .ZN(G405));
  NAND2_X1  g1087(.A1(new_n1246), .A2(new_n1263), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1270), .A2(new_n1245), .A3(new_n1242), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(KEYINPUT127), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT127), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1288), .A2(new_n1292), .A3(new_n1289), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(G375), .B(G378), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1294), .B(new_n1295), .ZN(G402));
endmodule


