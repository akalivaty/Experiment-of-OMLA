//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977;
  OR3_X1    g000(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n202));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT15), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G29gat), .A2(G36gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT90), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI211_X1 g008(.A(KEYINPUT90), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT91), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n206), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT91), .B1(new_n209), .B2(new_n210), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n202), .B(new_n205), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n203), .A2(new_n204), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n211), .A2(new_n202), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n203), .A2(new_n204), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n216), .A2(new_n206), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT92), .B(KEYINPUT17), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT93), .ZN(new_n223));
  INV_X1    g022(.A(G22gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G15gat), .ZN(new_n225));
  INV_X1    g024(.A(G15gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G22gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n223), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n225), .A2(new_n227), .A3(new_n223), .ZN(new_n230));
  INV_X1    g029(.A(G1gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT16), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  AND3_X1   g032(.A1(new_n225), .A2(new_n227), .A3(new_n223), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n231), .B1(new_n234), .B2(new_n228), .ZN(new_n235));
  XOR2_X1   g034(.A(KEYINPUT94), .B(G8gat), .Z(new_n236));
  NAND3_X1  g035(.A1(new_n233), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n233), .A2(new_n235), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n237), .A2(KEYINPUT95), .B1(new_n238), .B2(G8gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n215), .A2(new_n219), .A3(KEYINPUT17), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT95), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n233), .A2(new_n235), .A3(new_n241), .A4(new_n236), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n222), .A2(new_n239), .A3(new_n240), .A4(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n237), .A2(KEYINPUT95), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n238), .A2(G8gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n246), .A3(new_n242), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n220), .ZN(new_n248));
  NAND2_X1  g047(.A1(G229gat), .A2(G233gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT18), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT96), .B1(new_n244), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT96), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n243), .A2(new_n254), .A3(new_n248), .A4(new_n251), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n249), .B(KEYINPUT13), .Z(new_n256));
  NOR2_X1   g055(.A1(new_n247), .A2(new_n220), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n239), .A2(new_n242), .B1(new_n215), .B2(new_n219), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n253), .A2(new_n255), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT97), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n253), .A2(KEYINPUT97), .A3(new_n255), .A4(new_n259), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n243), .A2(new_n248), .A3(new_n249), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT18), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n268));
  XNOR2_X1  g067(.A(G113gat), .B(G141gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G169gat), .B(G197gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(KEYINPUT12), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n273), .B(KEYINPUT89), .Z(new_n274));
  NAND2_X1  g073(.A1(new_n267), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n253), .A2(new_n255), .A3(new_n259), .A4(new_n273), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n266), .A2(KEYINPUT98), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT98), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n278), .B1(new_n264), .B2(new_n265), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n276), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n275), .A2(new_n281), .A3(KEYINPUT99), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT99), .ZN(new_n283));
  INV_X1    g082(.A(new_n274), .ZN(new_n284));
  INV_X1    g083(.A(new_n266), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n285), .B1(new_n260), .B2(new_n261), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n284), .B1(new_n286), .B2(new_n263), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n283), .B1(new_n287), .B2(new_n280), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G120gat), .ZN(new_n291));
  OR3_X1    g090(.A1(new_n291), .A2(KEYINPUT67), .A3(G113gat), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT67), .B1(new_n291), .B2(G113gat), .ZN(new_n293));
  INV_X1    g092(.A(G113gat), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n292), .B(new_n293), .C1(new_n294), .C2(G120gat), .ZN(new_n295));
  XOR2_X1   g094(.A(G127gat), .B(G134gat), .Z(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(KEYINPUT1), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n294), .A2(G120gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n291), .A2(G113gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n295), .A2(new_n297), .B1(new_n301), .B2(new_n296), .ZN(new_n302));
  AND2_X1   g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(G141gat), .A2(G148gat), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT73), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n308), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(new_n311), .A3(new_n306), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT2), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n303), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n309), .B(new_n312), .C1(new_n317), .C2(KEYINPUT75), .ZN(new_n318));
  NAND2_X1  g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319));
  AND2_X1   g118(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n320));
  NOR2_X1   g119(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n321));
  OAI211_X1 g120(.A(KEYINPUT75), .B(new_n319), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n305), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n304), .A2(new_n314), .ZN(new_n325));
  AOI211_X1 g124(.A(new_n308), .B(new_n307), .C1(new_n325), .C2(new_n319), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n302), .B1(new_n328), .B2(KEYINPUT3), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n332), .A2(new_n322), .A3(new_n309), .A4(new_n312), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n326), .B1(new_n333), .B2(new_n305), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n335), .B1(new_n334), .B2(new_n336), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n329), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT78), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n329), .B(new_n341), .C1(new_n337), .C2(new_n338), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n324), .A2(new_n327), .A3(new_n302), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT4), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT81), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT82), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n349), .B1(new_n334), .B2(new_n302), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT82), .B1(new_n350), .B2(KEYINPUT81), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n349), .A3(new_n302), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n348), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n352), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n347), .B1(new_n345), .B2(new_n346), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n350), .A2(KEYINPUT81), .A3(KEYINPUT82), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(KEYINPUT5), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n343), .A2(new_n353), .A3(new_n357), .A4(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT83), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n351), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n340), .A2(new_n342), .B1(new_n364), .B2(new_n354), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n365), .A2(KEYINPUT83), .A3(new_n353), .A4(new_n360), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n302), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n328), .A2(new_n368), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n369), .A2(new_n344), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT5), .B1(new_n370), .B2(new_n358), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n350), .B(KEYINPUT79), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n352), .B(KEYINPUT80), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n359), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n371), .B1(new_n374), .B2(new_n343), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n367), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT87), .ZN(new_n378));
  XNOR2_X1  g177(.A(G1gat), .B(G29gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT0), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(G57gat), .ZN(new_n381));
  INV_X1    g180(.A(G85gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n377), .A2(new_n378), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n375), .B1(new_n363), .B2(new_n366), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT87), .B1(new_n386), .B2(new_n383), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT6), .B1(new_n386), .B2(new_n383), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT6), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n386), .A2(new_n390), .A3(new_n383), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT85), .ZN(new_n394));
  XOR2_X1   g193(.A(KEYINPUT71), .B(KEYINPUT29), .Z(new_n395));
  OAI21_X1  g194(.A(new_n395), .B1(new_n337), .B2(new_n338), .ZN(new_n396));
  XNOR2_X1  g195(.A(G197gat), .B(G204gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT70), .B(G211gat), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n398), .A2(G218gat), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n397), .B1(new_n399), .B2(KEYINPUT22), .ZN(new_n400));
  XNOR2_X1  g199(.A(G211gat), .B(G218gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n395), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n336), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n396), .A2(new_n402), .B1(new_n404), .B2(new_n328), .ZN(new_n405));
  INV_X1    g204(.A(G228gat), .ZN(new_n406));
  INV_X1    g205(.A(G233gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT84), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n401), .ZN(new_n410));
  OR2_X1    g209(.A1(new_n400), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n400), .A2(new_n410), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n403), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n336), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n328), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT77), .B1(new_n328), .B2(new_n414), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n403), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n402), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n415), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT84), .ZN(new_n421));
  INV_X1    g220(.A(new_n408), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n396), .A2(new_n402), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT3), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(new_n402), .B2(KEYINPUT29), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n422), .B1(new_n426), .B2(new_n328), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n409), .A2(new_n423), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n394), .B1(new_n428), .B2(new_n224), .ZN(new_n429));
  XNOR2_X1  g228(.A(G78gat), .B(G106gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT31), .B(G50gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n424), .A2(new_n427), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n405), .A2(KEYINPUT84), .A3(new_n408), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n421), .B1(new_n420), .B2(new_n422), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G22gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n428), .A2(new_n224), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n433), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT85), .A4(new_n432), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G226gat), .A2(G233gat), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(G169gat), .A2(G176gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT23), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT23), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(G169gat), .B2(G176gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(G169gat), .A2(G176gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT24), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(G183gat), .A3(G190gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(G183gat), .B(G190gat), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n453), .B1(new_n454), .B2(new_n452), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n451), .B1(new_n455), .B2(KEYINPUT64), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT64), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n457), .B(new_n453), .C1(new_n454), .C2(new_n452), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT25), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n447), .A2(KEYINPUT25), .A3(new_n449), .A4(new_n450), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT65), .ZN(new_n463));
  OR3_X1    g262(.A1(new_n455), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n463), .B1(new_n455), .B2(new_n462), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT26), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n446), .A2(KEYINPUT66), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT66), .B1(new_n446), .B2(new_n468), .ZN(new_n470));
  OAI221_X1 g269(.A(new_n450), .B1(new_n468), .B2(new_n446), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(KEYINPUT27), .B(G183gat), .ZN(new_n472));
  INV_X1    g271(.A(G190gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n474), .A2(KEYINPUT28), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n474), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n471), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n467), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n445), .B1(new_n478), .B2(new_n395), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n459), .A2(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n480));
  INV_X1    g279(.A(new_n477), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(new_n444), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n402), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n444), .B1(new_n482), .B2(KEYINPUT29), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n478), .A2(new_n445), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n486), .A3(new_n419), .ZN(new_n487));
  XNOR2_X1  g286(.A(G8gat), .B(G36gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(G64gat), .ZN(new_n489));
  INV_X1    g288(.A(G92gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n484), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT30), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n491), .ZN(new_n495));
  INV_X1    g294(.A(new_n484), .ZN(new_n496));
  INV_X1    g295(.A(new_n487), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT72), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n492), .A2(new_n499), .A3(new_n493), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n499), .B1(new_n492), .B2(new_n493), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n494), .B(new_n498), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n467), .A2(new_n368), .A3(new_n477), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n302), .B1(new_n480), .B2(new_n481), .ZN(new_n504));
  NAND2_X1  g303(.A1(G227gat), .A2(G233gat), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT32), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT33), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g309(.A(G15gat), .B(G43gat), .Z(new_n511));
  XNOR2_X1  g310(.A(G71gat), .B(G99gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n508), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n513), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n507), .B(KEYINPUT32), .C1(new_n509), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n503), .A2(new_n504), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT34), .B1(new_n518), .B2(new_n505), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(KEYINPUT34), .A3(new_n505), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n517), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n521), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n514), .B(new_n516), .C1(new_n519), .C2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT35), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n502), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n393), .A2(new_n443), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n377), .A2(new_n384), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n388), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n502), .B1(new_n530), .B2(new_n392), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT68), .B1(new_n523), .B2(new_n519), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT68), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n520), .A2(new_n533), .A3(new_n521), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT69), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT69), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n517), .A2(new_n532), .A3(new_n534), .A4(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n538), .A3(new_n524), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n539), .B1(new_n441), .B2(new_n442), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n531), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n528), .B1(new_n541), .B2(new_n525), .ZN(new_n542));
  INV_X1    g341(.A(new_n443), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n391), .B1(new_n529), .B2(new_n388), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n543), .B1(new_n544), .B2(new_n502), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n522), .A2(new_n524), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(KEYINPUT36), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n547), .B1(new_n539), .B2(KEYINPUT36), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT38), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT37), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n484), .A2(new_n550), .A3(new_n487), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n495), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT37), .B1(new_n496), .B2(new_n497), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n485), .A2(new_n486), .A3(new_n402), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT37), .ZN(new_n557));
  INV_X1    g356(.A(new_n479), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n402), .B1(new_n558), .B2(new_n486), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n549), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n492), .B1(new_n560), .B2(new_n552), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n389), .A2(new_n392), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n358), .B1(new_n365), .B2(new_n353), .ZN(new_n564));
  INV_X1    g363(.A(new_n370), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT39), .B1(new_n565), .B2(new_n359), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n343), .A2(new_n353), .A3(new_n357), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT86), .B(KEYINPUT39), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n359), .A3(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n567), .A2(KEYINPUT40), .A3(new_n383), .A4(new_n570), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n570), .B(new_n383), .C1(new_n564), .C2(new_n566), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT40), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(new_n574), .A3(new_n502), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n385), .A2(new_n387), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n443), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n545), .B(new_n548), .C1(new_n563), .C2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n290), .B1(new_n542), .B2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G57gat), .B(G64gat), .Z(new_n580));
  INV_X1    g379(.A(KEYINPUT9), .ZN(new_n581));
  INV_X1    g380(.A(G71gat), .ZN(new_n582));
  INV_X1    g381(.A(G78gat), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G71gat), .B(G78gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n580), .A2(new_n586), .A3(new_n584), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n247), .B1(KEYINPUT21), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(G183gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(KEYINPUT100), .B(KEYINPUT21), .Z(new_n594));
  NOR2_X1   g393(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n593), .A2(new_n597), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G127gat), .B(G155gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n604), .B(G211gat), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n601), .B(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT8), .ZN(new_n607));
  NAND2_X1  g406(.A1(G99gat), .A2(G106gat), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n607), .B1(new_n608), .B2(KEYINPUT102), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT102), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n610), .A2(G99gat), .A3(G106gat), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n609), .A2(new_n611), .B1(new_n382), .B2(new_n490), .ZN(new_n612));
  XNOR2_X1  g411(.A(G99gat), .B(G106gat), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT7), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n614), .B(new_n615), .C1(new_n382), .C2(new_n490), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n614), .B1(new_n382), .B2(new_n490), .ZN(new_n617));
  NAND3_X1  g416(.A1(KEYINPUT101), .A2(G85gat), .A3(G92gat), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(KEYINPUT7), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n612), .A2(new_n613), .A3(new_n616), .A4(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n612), .A2(new_n616), .A3(new_n619), .ZN(new_n622));
  INV_X1    g421(.A(new_n613), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n222), .B(new_n240), .C1(new_n621), .C2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n621), .ZN(new_n626));
  AND2_X1   g425(.A1(G232gat), .A2(G233gat), .ZN(new_n627));
  AOI22_X1  g426(.A1(new_n626), .A2(new_n220), .B1(KEYINPUT41), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G190gat), .B(G218gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT103), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n629), .A2(new_n631), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G134gat), .B(G162gat), .Z(new_n635));
  NOR2_X1   g434(.A1(new_n627), .A2(KEYINPUT41), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(KEYINPUT104), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(KEYINPUT104), .Z(new_n639));
  OAI21_X1  g438(.A(new_n639), .B1(new_n632), .B2(new_n633), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n606), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(G230gat), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n643), .A2(new_n407), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n613), .A2(KEYINPUT105), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n588), .A2(new_n589), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n624), .B2(new_n621), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n622), .A2(new_n623), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n590), .A2(new_n620), .A3(new_n648), .A4(new_n645), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n647), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n626), .A2(KEYINPUT10), .A3(new_n590), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n644), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n647), .A2(new_n649), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n644), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G120gat), .B(G148gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G176gat), .ZN(new_n659));
  INV_X1    g458(.A(G204gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n654), .A2(new_n656), .A3(new_n661), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n642), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n579), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n544), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n668), .A2(KEYINPUT106), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(KEYINPUT106), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g473(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n675));
  NAND2_X1  g474(.A1(new_n667), .A2(new_n502), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT108), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT16), .B(G8gat), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n675), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n676), .A2(new_n680), .A3(new_n678), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n681), .B1(new_n677), .B2(G8gat), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n682), .ZN(G1325gat));
  INV_X1    g482(.A(new_n546), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n226), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n548), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n667), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n687), .B2(new_n226), .ZN(G1326gat));
  NAND2_X1  g487(.A1(new_n667), .A2(new_n543), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT43), .B(G22gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  INV_X1    g490(.A(new_n606), .ZN(new_n692));
  INV_X1    g491(.A(new_n641), .ZN(new_n693));
  INV_X1    g492(.A(new_n665), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT109), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n579), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(G29gat), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n699), .A3(new_n672), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT45), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n287), .A2(new_n280), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n563), .A2(new_n577), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n548), .B1(new_n531), .B2(new_n443), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n525), .B1(new_n531), .B2(new_n540), .ZN(new_n706));
  INV_X1    g505(.A(new_n442), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n429), .A2(new_n432), .B1(new_n438), .B2(new_n439), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n527), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n392), .B2(new_n389), .ZN(new_n710));
  OAI22_X1  g509(.A1(new_n704), .A2(new_n705), .B1(new_n706), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT111), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n542), .A2(new_n578), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n641), .A2(KEYINPUT44), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n711), .A2(new_n693), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT44), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n606), .B(KEYINPUT110), .Z(new_n720));
  AND4_X1   g519(.A1(new_n703), .A2(new_n719), .A3(new_n694), .A4(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n721), .A2(new_n672), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n701), .B1(new_n722), .B2(new_n699), .ZN(G1328gat));
  INV_X1    g522(.A(G36gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n698), .A2(new_n724), .A3(new_n502), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT46), .Z(new_n726));
  AND2_X1   g525(.A1(new_n721), .A2(new_n502), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(new_n724), .ZN(G1329gat));
  NOR3_X1   g527(.A1(new_n697), .A2(G43gat), .A3(new_n546), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n721), .A2(new_n686), .ZN(new_n731));
  INV_X1    g530(.A(G43gat), .ZN(new_n732));
  OAI211_X1 g531(.A(KEYINPUT47), .B(new_n730), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT47), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n732), .B1(new_n721), .B2(new_n686), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(new_n729), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n733), .A2(new_n736), .ZN(G1330gat));
  NOR3_X1   g536(.A1(new_n697), .A2(G50gat), .A3(new_n443), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n721), .A2(new_n543), .ZN(new_n740));
  INV_X1    g539(.A(G50gat), .ZN(new_n741));
  OAI211_X1 g540(.A(KEYINPUT48), .B(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n741), .B1(new_n721), .B2(new_n543), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(new_n738), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n745), .ZN(G1331gat));
  AND2_X1   g545(.A1(new_n712), .A2(new_n714), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n642), .A2(new_n703), .A3(new_n694), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n672), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g551(.A(new_n502), .B(KEYINPUT112), .Z(new_n753));
  AOI21_X1  g552(.A(new_n753), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT113), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n755), .A2(KEYINPUT113), .ZN(new_n758));
  OAI22_X1  g557(.A1(new_n757), .A2(new_n758), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n759));
  INV_X1    g558(.A(new_n758), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n760), .A2(new_n761), .A3(new_n756), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(G1333gat));
  XNOR2_X1  g562(.A(new_n546), .B(KEYINPUT114), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n582), .B1(new_n749), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n686), .A2(G71gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n749), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g567(.A1(new_n749), .A2(new_n443), .ZN(new_n769));
  XOR2_X1   g568(.A(KEYINPUT115), .B(G78gat), .Z(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1335gat));
  NOR2_X1   g570(.A1(new_n703), .A2(new_n606), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n711), .A2(new_n693), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n694), .B1(new_n773), .B2(KEYINPUT51), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n711), .A2(new_n775), .A3(new_n693), .A4(new_n772), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(new_n382), .A3(new_n672), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n772), .A2(new_n665), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n716), .B2(new_n718), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(new_n672), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n778), .B1(new_n781), .B2(new_n382), .ZN(G1336gat));
  INV_X1    g581(.A(KEYINPUT118), .ZN(new_n783));
  XNOR2_X1  g582(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n784));
  AOI211_X1 g583(.A(new_n753), .B(new_n779), .C1(new_n716), .C2(new_n718), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n785), .B2(new_n490), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n773), .A2(KEYINPUT51), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n753), .A2(G92gat), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n787), .A2(new_n665), .A3(new_n776), .A4(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n774), .A2(KEYINPUT116), .A3(new_n776), .A4(new_n788), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n786), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795));
  INV_X1    g594(.A(new_n779), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n719), .A2(new_n502), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G92gat), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n795), .B1(new_n798), .B2(new_n789), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n783), .B1(new_n794), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n490), .B1(new_n780), .B2(new_n502), .ZN(new_n801));
  INV_X1    g600(.A(new_n789), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT52), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n803), .B(KEYINPUT118), .C1(new_n786), .C2(new_n793), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n800), .A2(new_n804), .ZN(G1337gat));
  AOI21_X1  g604(.A(G99gat), .B1(new_n777), .B2(new_n684), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n686), .A2(G99gat), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n780), .B2(new_n807), .ZN(G1338gat));
  NAND2_X1  g607(.A1(new_n780), .A2(new_n543), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n443), .A2(G106gat), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n809), .A2(G106gat), .B1(new_n777), .B2(new_n810), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT53), .Z(G1339gat));
  NAND2_X1  g611(.A1(new_n672), .A2(new_n753), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n642), .A2(new_n703), .A3(new_n665), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n653), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n644), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n651), .A2(new_n652), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n820));
  AOI211_X1 g619(.A(new_n820), .B(new_n661), .C1(new_n653), .C2(new_n815), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(new_n815), .A3(new_n817), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT119), .B1(new_n822), .B2(new_n662), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n819), .B(KEYINPUT55), .C1(new_n821), .C2(new_n823), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n824), .A2(KEYINPUT120), .A3(new_n664), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT120), .B1(new_n824), .B2(new_n664), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n819), .B1(new_n821), .B2(new_n823), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n825), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  OR3_X1    g629(.A1(new_n257), .A2(new_n258), .A3(new_n256), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT121), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n244), .A2(new_n258), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(new_n249), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n831), .A2(new_n832), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n272), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n830), .A2(new_n281), .A3(new_n693), .A4(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n281), .A2(new_n665), .A3(new_n837), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n840), .B1(new_n830), .B2(new_n703), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n838), .B1(new_n841), .B2(new_n693), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n814), .B1(new_n842), .B2(new_n720), .ZN(new_n843));
  NOR4_X1   g642(.A1(new_n813), .A2(new_n843), .A3(new_n543), .A4(new_n546), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n290), .A2(new_n294), .ZN(new_n845));
  INV_X1    g644(.A(new_n540), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n843), .A2(new_n671), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n703), .A3(new_n753), .ZN(new_n848));
  AOI22_X1  g647(.A1(new_n844), .A2(new_n845), .B1(new_n294), .B2(new_n848), .ZN(G1340gat));
  NAND3_X1  g648(.A1(new_n844), .A2(G120gat), .A3(new_n665), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(new_n753), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n291), .B1(new_n851), .B2(new_n694), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT122), .ZN(G1341gat));
  INV_X1    g653(.A(G127gat), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n606), .B(KEYINPUT110), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n844), .B2(new_n856), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n851), .A2(G127gat), .A3(new_n692), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n857), .A2(new_n858), .ZN(G1342gat));
  OR2_X1    g658(.A1(new_n502), .A2(new_n641), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n860), .A2(G134gat), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n847), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT56), .Z(new_n863));
  NAND2_X1  g662(.A1(new_n844), .A2(new_n693), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n864), .A2(KEYINPUT123), .A3(G134gat), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT123), .B1(new_n864), .B2(G134gat), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n863), .B1(new_n865), .B2(new_n866), .ZN(G1343gat));
  NOR2_X1   g666(.A1(new_n813), .A2(new_n686), .ZN(new_n868));
  INV_X1    g667(.A(new_n843), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT57), .B1(new_n869), .B2(new_n543), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n443), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n824), .A2(new_n664), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n829), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT99), .B1(new_n275), .B2(new_n281), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n287), .A2(new_n283), .A3(new_n280), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n693), .B1(new_n878), .B2(new_n839), .ZN(new_n879));
  INV_X1    g678(.A(new_n838), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n692), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n814), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n873), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n868), .B1(new_n870), .B2(new_n883), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n884), .A2(new_n290), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(G141gat), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n843), .A2(new_n671), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n686), .A2(new_n443), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n753), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n891), .A2(G141gat), .A3(new_n290), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n892), .A2(KEYINPUT58), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n884), .A2(new_n702), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n892), .B1(new_n894), .B2(G141gat), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n886), .A2(new_n893), .B1(new_n895), .B2(new_n896), .ZN(G1344gat));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n898), .B(G148gat), .C1(new_n884), .C2(new_n694), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n666), .A2(new_n290), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n443), .B1(new_n881), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT125), .B1(new_n902), .B2(KEYINPUT57), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT124), .B1(new_n843), .B2(new_n873), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n826), .A2(new_n829), .ZN(new_n906));
  INV_X1    g705(.A(new_n825), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n839), .B1(new_n908), .B2(new_n702), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n641), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n856), .B1(new_n910), .B2(new_n838), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n905), .B(new_n872), .C1(new_n911), .C2(new_n814), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n904), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n840), .B1(new_n289), .B2(new_n875), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n838), .B1(new_n915), .B2(new_n693), .ZN(new_n916));
  AOI22_X1  g715(.A1(new_n916), .A2(new_n692), .B1(new_n290), .B2(new_n666), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n914), .B(new_n871), .C1(new_n917), .C2(new_n443), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n903), .A2(new_n913), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n665), .A3(new_n868), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(G148gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n900), .B1(new_n921), .B2(KEYINPUT59), .ZN(new_n922));
  AOI211_X1 g721(.A(KEYINPUT126), .B(new_n898), .C1(new_n920), .C2(G148gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n899), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OR3_X1    g723(.A1(new_n891), .A2(G148gat), .A3(new_n694), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1345gat));
  OAI21_X1  g725(.A(G155gat), .B1(new_n884), .B2(new_n720), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n692), .A2(G155gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n891), .B2(new_n928), .ZN(G1346gat));
  OAI21_X1  g728(.A(G162gat), .B1(new_n884), .B2(new_n641), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n860), .A2(G162gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n889), .B2(new_n931), .ZN(G1347gat));
  NAND2_X1  g731(.A1(new_n671), .A2(new_n502), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n933), .A2(new_n764), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n843), .A2(new_n543), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n937), .A2(G169gat), .A3(new_n289), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n672), .A2(new_n843), .ZN(new_n939));
  INV_X1    g738(.A(new_n753), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n540), .A3(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(G169gat), .B1(new_n942), .B2(new_n703), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n938), .A2(new_n943), .ZN(G1348gat));
  NAND3_X1  g743(.A1(new_n937), .A2(G176gat), .A3(new_n665), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  AOI21_X1  g747(.A(G176gat), .B1(new_n942), .B2(new_n665), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(G1349gat));
  OAI21_X1  g749(.A(G183gat), .B1(new_n936), .B2(new_n720), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n606), .A2(new_n472), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n941), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g753(.A1(new_n942), .A2(new_n473), .A3(new_n693), .ZN(new_n955));
  OAI21_X1  g754(.A(G190gat), .B1(new_n936), .B2(new_n641), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n956), .A2(KEYINPUT61), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n956), .A2(KEYINPUT61), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1351gat));
  NOR2_X1   g758(.A1(new_n933), .A2(new_n686), .ZN(new_n960));
  AND4_X1   g759(.A1(G197gat), .A2(new_n919), .A3(new_n289), .A4(new_n960), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n686), .A2(new_n753), .A3(new_n443), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n939), .A2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(G197gat), .B1(new_n964), .B2(new_n703), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n961), .A2(new_n965), .ZN(G1352gat));
  NOR3_X1   g765(.A1(new_n963), .A2(G204gat), .A3(new_n694), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n967), .B(KEYINPUT62), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n919), .A2(new_n665), .A3(new_n960), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n660), .B2(new_n969), .ZN(G1353gat));
  OR3_X1    g769(.A1(new_n963), .A2(new_n398), .A3(new_n692), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n919), .A2(new_n606), .A3(new_n960), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n972), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT63), .B1(new_n972), .B2(G211gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(G1354gat));
  AND4_X1   g774(.A1(G218gat), .A2(new_n919), .A3(new_n693), .A4(new_n960), .ZN(new_n976));
  AOI21_X1  g775(.A(G218gat), .B1(new_n964), .B2(new_n693), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n976), .A2(new_n977), .ZN(G1355gat));
endmodule


