

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590;

  XNOR2_X1 U321 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U322 ( .A(n424), .B(n423), .ZN(n537) );
  XNOR2_X1 U323 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n423) );
  NOR2_X1 U324 ( .A1(n422), .A2(n421), .ZN(n424) );
  XNOR2_X1 U325 ( .A(n388), .B(n387), .ZN(n565) );
  XOR2_X1 U326 ( .A(n353), .B(n309), .Z(n529) );
  NAND2_X1 U327 ( .A1(n529), .A2(n558), .ZN(n289) );
  INV_X1 U328 ( .A(KEYINPUT113), .ZN(n408) );
  XNOR2_X1 U329 ( .A(n408), .B(KEYINPUT45), .ZN(n409) );
  XNOR2_X1 U330 ( .A(n410), .B(n409), .ZN(n411) );
  INV_X1 U331 ( .A(KEYINPUT47), .ZN(n418) );
  XNOR2_X1 U332 ( .A(n418), .B(KEYINPUT112), .ZN(n419) );
  XNOR2_X1 U333 ( .A(n420), .B(n419), .ZN(n421) );
  INV_X1 U334 ( .A(G92GAT), .ZN(n375) );
  XNOR2_X1 U335 ( .A(n457), .B(n326), .ZN(n327) );
  NOR2_X1 U336 ( .A1(n524), .A2(n442), .ZN(n444) );
  XNOR2_X1 U337 ( .A(n328), .B(n327), .ZN(n334) );
  XNOR2_X1 U338 ( .A(n378), .B(n377), .ZN(n379) );
  NOR2_X1 U339 ( .A1(n538), .A2(n465), .ZN(n570) );
  XOR2_X1 U340 ( .A(n481), .B(KEYINPUT28), .Z(n539) );
  XNOR2_X1 U341 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n466) );
  XNOR2_X1 U342 ( .A(n467), .B(n466), .ZN(G1351GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT82), .B(G134GAT), .Z(n291) );
  XNOR2_X1 U344 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n290) );
  XNOR2_X1 U345 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U346 ( .A(G113GAT), .B(n292), .Z(n353) );
  XOR2_X1 U347 ( .A(G190GAT), .B(G99GAT), .Z(n294) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(G15GAT), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U350 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n296) );
  XNOR2_X1 U351 ( .A(G183GAT), .B(G176GAT), .ZN(n295) );
  XNOR2_X1 U352 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U353 ( .A(n298), .B(n297), .Z(n308) );
  XOR2_X1 U354 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n300) );
  XNOR2_X1 U355 ( .A(KEYINPUT85), .B(KEYINPUT20), .ZN(n299) );
  XNOR2_X1 U356 ( .A(n300), .B(n299), .ZN(n306) );
  XOR2_X1 U357 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n302) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n301) );
  XNOR2_X1 U359 ( .A(n302), .B(n301), .ZN(n436) );
  XOR2_X1 U360 ( .A(G120GAT), .B(G71GAT), .Z(n315) );
  XOR2_X1 U361 ( .A(n436), .B(n315), .Z(n304) );
  NAND2_X1 U362 ( .A1(G227GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U363 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U364 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U365 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U366 ( .A(KEYINPUT70), .B(KEYINPUT31), .Z(n314) );
  INV_X1 U367 ( .A(KEYINPUT13), .ZN(n310) );
  NAND2_X1 U368 ( .A1(G57GAT), .A2(n310), .ZN(n313) );
  INV_X1 U369 ( .A(G57GAT), .ZN(n311) );
  NAND2_X1 U370 ( .A1(n311), .A2(KEYINPUT13), .ZN(n312) );
  NAND2_X1 U371 ( .A1(n313), .A2(n312), .ZN(n395) );
  XNOR2_X1 U372 ( .A(n314), .B(n395), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n316), .B(n315), .ZN(n321) );
  INV_X1 U374 ( .A(n321), .ZN(n320) );
  XOR2_X1 U375 ( .A(KEYINPUT32), .B(KEYINPUT74), .Z(n318) );
  XNOR2_X1 U376 ( .A(KEYINPUT73), .B(KEYINPUT33), .ZN(n317) );
  XNOR2_X1 U377 ( .A(n318), .B(n317), .ZN(n322) );
  INV_X1 U378 ( .A(n322), .ZN(n319) );
  NAND2_X1 U379 ( .A1(n320), .A2(n319), .ZN(n324) );
  NAND2_X1 U380 ( .A1(n322), .A2(n321), .ZN(n323) );
  NAND2_X1 U381 ( .A1(n324), .A2(n323), .ZN(n328) );
  XNOR2_X1 U382 ( .A(G148GAT), .B(G106GAT), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n325), .B(G78GAT), .ZN(n457) );
  NAND2_X1 U384 ( .A1(G230GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U385 ( .A(G99GAT), .B(G85GAT), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n329), .B(KEYINPUT71), .ZN(n373) );
  XOR2_X1 U387 ( .A(G204GAT), .B(KEYINPUT72), .Z(n331) );
  XNOR2_X1 U388 ( .A(G92GAT), .B(G64GAT), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U390 ( .A(G176GAT), .B(n332), .Z(n435) );
  XNOR2_X1 U391 ( .A(n373), .B(n435), .ZN(n333) );
  XNOR2_X1 U392 ( .A(n334), .B(n333), .ZN(n372) );
  XOR2_X1 U393 ( .A(n372), .B(KEYINPUT41), .Z(n558) );
  XOR2_X1 U394 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n336) );
  XNOR2_X1 U395 ( .A(G57GAT), .B(KEYINPUT1), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U397 ( .A(G148GAT), .B(n337), .Z(n339) );
  NAND2_X1 U398 ( .A1(G225GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U400 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n341) );
  XNOR2_X1 U401 ( .A(KEYINPUT88), .B(G155GAT), .ZN(n340) );
  XNOR2_X1 U402 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U403 ( .A(KEYINPUT89), .B(n342), .Z(n458) );
  XOR2_X1 U404 ( .A(n343), .B(n458), .Z(n345) );
  XNOR2_X1 U405 ( .A(G1GAT), .B(G141GAT), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U407 ( .A(KEYINPUT5), .B(G85GAT), .Z(n347) );
  XNOR2_X1 U408 ( .A(G29GAT), .B(G162GAT), .ZN(n346) );
  XNOR2_X1 U409 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U410 ( .A(n349), .B(n348), .Z(n355) );
  XOR2_X1 U411 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n351) );
  XNOR2_X1 U412 ( .A(G120GAT), .B(KEYINPUT94), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U415 ( .A(n355), .B(n354), .Z(n479) );
  INV_X1 U416 ( .A(n479), .ZN(n524) );
  INV_X1 U417 ( .A(KEYINPUT54), .ZN(n441) );
  XNOR2_X1 U418 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n356) );
  XNOR2_X1 U419 ( .A(n356), .B(G15GAT), .ZN(n394) );
  XOR2_X1 U420 ( .A(G141GAT), .B(G22GAT), .Z(n448) );
  XOR2_X1 U421 ( .A(n394), .B(n448), .Z(n358) );
  NAND2_X1 U422 ( .A1(G229GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n359), .B(G197GAT), .ZN(n363) );
  XOR2_X1 U425 ( .A(G29GAT), .B(G43GAT), .Z(n361) );
  XNOR2_X1 U426 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n360) );
  XNOR2_X1 U427 ( .A(n361), .B(n360), .ZN(n378) );
  XOR2_X1 U428 ( .A(n378), .B(KEYINPUT67), .Z(n362) );
  XNOR2_X1 U429 ( .A(n363), .B(n362), .ZN(n371) );
  XOR2_X1 U430 ( .A(G8GAT), .B(G113GAT), .Z(n365) );
  XNOR2_X1 U431 ( .A(G50GAT), .B(G36GAT), .ZN(n364) );
  XNOR2_X1 U432 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U433 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n367) );
  XNOR2_X1 U434 ( .A(G169GAT), .B(KEYINPUT68), .ZN(n366) );
  XNOR2_X1 U435 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U436 ( .A(n369), .B(n368), .Z(n370) );
  XOR2_X1 U437 ( .A(n371), .B(n370), .Z(n574) );
  INV_X1 U438 ( .A(n574), .ZN(n568) );
  XOR2_X1 U439 ( .A(G50GAT), .B(G162GAT), .Z(n447) );
  XNOR2_X1 U440 ( .A(n447), .B(n373), .ZN(n374) );
  XOR2_X1 U441 ( .A(G36GAT), .B(G190GAT), .Z(n429) );
  XNOR2_X1 U442 ( .A(n374), .B(n429), .ZN(n380) );
  NAND2_X1 U443 ( .A1(G232GAT), .A2(G233GAT), .ZN(n376) );
  XOR2_X1 U444 ( .A(n380), .B(n379), .Z(n388) );
  XOR2_X1 U445 ( .A(KEYINPUT66), .B(KEYINPUT9), .Z(n382) );
  XNOR2_X1 U446 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n381) );
  XNOR2_X1 U447 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U448 ( .A(G106GAT), .B(KEYINPUT10), .Z(n384) );
  XNOR2_X1 U449 ( .A(G134GAT), .B(KEYINPUT76), .ZN(n383) );
  XNOR2_X1 U450 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U451 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U452 ( .A(KEYINPUT36), .B(n565), .ZN(n585) );
  XOR2_X1 U453 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n390) );
  XNOR2_X1 U454 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n389) );
  XNOR2_X1 U455 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U456 ( .A(G8GAT), .B(G183GAT), .Z(n428) );
  XOR2_X1 U457 ( .A(n391), .B(n428), .Z(n393) );
  XNOR2_X1 U458 ( .A(G127GAT), .B(G155GAT), .ZN(n392) );
  XNOR2_X1 U459 ( .A(n393), .B(n392), .ZN(n399) );
  XOR2_X1 U460 ( .A(n395), .B(n394), .Z(n397) );
  NAND2_X1 U461 ( .A1(G231GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U463 ( .A(n399), .B(n398), .Z(n407) );
  XOR2_X1 U464 ( .A(G211GAT), .B(KEYINPUT80), .Z(n401) );
  XNOR2_X1 U465 ( .A(KEYINPUT77), .B(KEYINPUT79), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U467 ( .A(G64GAT), .B(G78GAT), .Z(n403) );
  XNOR2_X1 U468 ( .A(G22GAT), .B(G71GAT), .ZN(n402) );
  XNOR2_X1 U469 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U470 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U471 ( .A(n407), .B(n406), .Z(n469) );
  INV_X1 U472 ( .A(n469), .ZN(n583) );
  NAND2_X1 U473 ( .A1(n585), .A2(n583), .ZN(n410) );
  NOR2_X1 U474 ( .A1(n372), .A2(n411), .ZN(n412) );
  XOR2_X1 U475 ( .A(KEYINPUT114), .B(n412), .Z(n413) );
  NOR2_X1 U476 ( .A1(n568), .A2(n413), .ZN(n422) );
  AND2_X1 U477 ( .A1(n568), .A2(n558), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n414), .B(KEYINPUT46), .ZN(n415) );
  NOR2_X1 U479 ( .A1(n415), .A2(n583), .ZN(n416) );
  XNOR2_X1 U480 ( .A(n416), .B(KEYINPUT111), .ZN(n417) );
  NOR2_X1 U481 ( .A1(n565), .A2(n417), .ZN(n420) );
  XOR2_X1 U482 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n426) );
  NAND2_X1 U483 ( .A1(G226GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U485 ( .A(n427), .B(KEYINPUT97), .Z(n431) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n434) );
  XOR2_X1 U488 ( .A(KEYINPUT21), .B(G211GAT), .Z(n433) );
  XNOR2_X1 U489 ( .A(G197GAT), .B(G218GAT), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n455) );
  XOR2_X1 U491 ( .A(n434), .B(n455), .Z(n438) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U493 ( .A(n438), .B(n437), .Z(n527) );
  INV_X1 U494 ( .A(n527), .ZN(n439) );
  NOR2_X1 U495 ( .A1(n537), .A2(n439), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n442) );
  INV_X1 U497 ( .A(KEYINPUT65), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n572) );
  XOR2_X1 U499 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n446) );
  XNOR2_X1 U500 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n445) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n452) );
  XOR2_X1 U502 ( .A(KEYINPUT23), .B(G204GAT), .Z(n450) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U505 ( .A(n452), .B(n451), .Z(n454) );
  NAND2_X1 U506 ( .A1(G228GAT), .A2(G233GAT), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n456) );
  XOR2_X1 U508 ( .A(n456), .B(n455), .Z(n460) );
  XNOR2_X1 U509 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U510 ( .A(n460), .B(n459), .ZN(n481) );
  AND2_X1 U511 ( .A1(n572), .A2(n481), .ZN(n461) );
  XNOR2_X1 U512 ( .A(n461), .B(KEYINPUT55), .ZN(n465) );
  OR2_X1 U513 ( .A1(n289), .A2(n465), .ZN(n464) );
  XOR2_X1 U514 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n462) );
  XNOR2_X1 U515 ( .A(n462), .B(G176GAT), .ZN(n463) );
  XNOR2_X1 U516 ( .A(n464), .B(n463), .ZN(G1349GAT) );
  INV_X1 U517 ( .A(n529), .ZN(n538) );
  NAND2_X1 U518 ( .A1(n570), .A2(n565), .ZN(n467) );
  XOR2_X1 U519 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n488) );
  NOR2_X1 U520 ( .A1(n574), .A2(n372), .ZN(n468) );
  XNOR2_X1 U521 ( .A(n468), .B(KEYINPUT75), .ZN(n499) );
  NOR2_X1 U522 ( .A1(n565), .A2(n469), .ZN(n470) );
  XOR2_X1 U523 ( .A(KEYINPUT16), .B(n470), .Z(n471) );
  XNOR2_X1 U524 ( .A(n471), .B(KEYINPUT81), .ZN(n486) );
  NAND2_X1 U525 ( .A1(n529), .A2(n527), .ZN(n472) );
  NAND2_X1 U526 ( .A1(n481), .A2(n472), .ZN(n473) );
  XOR2_X1 U527 ( .A(KEYINPUT25), .B(n473), .Z(n477) );
  XNOR2_X1 U528 ( .A(KEYINPUT98), .B(KEYINPUT26), .ZN(n475) );
  NOR2_X1 U529 ( .A1(n529), .A2(n481), .ZN(n474) );
  XNOR2_X1 U530 ( .A(n475), .B(n474), .ZN(n573) );
  XNOR2_X1 U531 ( .A(n527), .B(KEYINPUT27), .ZN(n482) );
  NAND2_X1 U532 ( .A1(n573), .A2(n482), .ZN(n476) );
  NAND2_X1 U533 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U534 ( .A1(n479), .A2(n478), .ZN(n480) );
  XOR2_X1 U535 ( .A(KEYINPUT99), .B(n480), .Z(n485) );
  NAND2_X1 U536 ( .A1(n524), .A2(n482), .ZN(n536) );
  NOR2_X1 U537 ( .A1(n539), .A2(n536), .ZN(n483) );
  NAND2_X1 U538 ( .A1(n483), .A2(n538), .ZN(n484) );
  NAND2_X1 U539 ( .A1(n485), .A2(n484), .ZN(n496) );
  NAND2_X1 U540 ( .A1(n486), .A2(n496), .ZN(n510) );
  NOR2_X1 U541 ( .A1(n499), .A2(n510), .ZN(n494) );
  NAND2_X1 U542 ( .A1(n494), .A2(n524), .ZN(n487) );
  XNOR2_X1 U543 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U544 ( .A(G1GAT), .B(n489), .Z(G1324GAT) );
  XOR2_X1 U545 ( .A(G8GAT), .B(KEYINPUT101), .Z(n491) );
  NAND2_X1 U546 ( .A1(n494), .A2(n527), .ZN(n490) );
  XNOR2_X1 U547 ( .A(n491), .B(n490), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(G15GAT), .B(KEYINPUT35), .Z(n493) );
  NAND2_X1 U549 ( .A1(n494), .A2(n529), .ZN(n492) );
  XNOR2_X1 U550 ( .A(n493), .B(n492), .ZN(G1326GAT) );
  NAND2_X1 U551 ( .A1(n494), .A2(n539), .ZN(n495) );
  XNOR2_X1 U552 ( .A(n495), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U553 ( .A1(n585), .A2(n496), .ZN(n497) );
  NOR2_X1 U554 ( .A1(n497), .A2(n583), .ZN(n498) );
  XNOR2_X1 U555 ( .A(n498), .B(KEYINPUT37), .ZN(n522) );
  NOR2_X1 U556 ( .A1(n522), .A2(n499), .ZN(n500) );
  XNOR2_X1 U557 ( .A(KEYINPUT38), .B(n500), .ZN(n508) );
  NAND2_X1 U558 ( .A1(n524), .A2(n508), .ZN(n502) );
  XOR2_X1 U559 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n501) );
  XNOR2_X1 U560 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(n503), .ZN(G1328GAT) );
  XOR2_X1 U562 ( .A(G36GAT), .B(KEYINPUT103), .Z(n505) );
  NAND2_X1 U563 ( .A1(n508), .A2(n527), .ZN(n504) );
  XNOR2_X1 U564 ( .A(n505), .B(n504), .ZN(G1329GAT) );
  NAND2_X1 U565 ( .A1(n508), .A2(n529), .ZN(n506) );
  XNOR2_X1 U566 ( .A(n506), .B(KEYINPUT40), .ZN(n507) );
  XNOR2_X1 U567 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  NAND2_X1 U568 ( .A1(n508), .A2(n539), .ZN(n509) );
  XNOR2_X1 U569 ( .A(n509), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n513) );
  NAND2_X1 U571 ( .A1(n574), .A2(n558), .ZN(n521) );
  NOR2_X1 U572 ( .A1(n510), .A2(n521), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n511), .B(KEYINPUT104), .ZN(n518) );
  NAND2_X1 U574 ( .A1(n524), .A2(n518), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(n514), .ZN(G1332GAT) );
  NAND2_X1 U577 ( .A1(n518), .A2(n527), .ZN(n515) );
  XNOR2_X1 U578 ( .A(n515), .B(KEYINPUT106), .ZN(n516) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(n516), .ZN(G1333GAT) );
  NAND2_X1 U580 ( .A1(n518), .A2(n529), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n517), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U583 ( .A1(n539), .A2(n518), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(KEYINPUT108), .ZN(n526) );
  NOR2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U587 ( .A(KEYINPUT107), .B(n523), .Z(n532) );
  NAND2_X1 U588 ( .A1(n524), .A2(n532), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n526), .B(n525), .ZN(G1336GAT) );
  NAND2_X1 U590 ( .A1(n527), .A2(n532), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U592 ( .A(G99GAT), .B(KEYINPUT109), .Z(n531) );
  NAND2_X1 U593 ( .A1(n532), .A2(n529), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n531), .B(n530), .ZN(G1338GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n534) );
  NAND2_X1 U596 ( .A1(n532), .A2(n539), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U598 ( .A(G106GAT), .B(n535), .Z(G1339GAT) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(KEYINPUT116), .ZN(n543) );
  NOR2_X1 U600 ( .A1(n537), .A2(n536), .ZN(n554) );
  NOR2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U602 ( .A1(n554), .A2(n540), .ZN(n541) );
  XNOR2_X1 U603 ( .A(KEYINPUT115), .B(n541), .ZN(n550) );
  NAND2_X1 U604 ( .A1(n550), .A2(n568), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n543), .B(n542), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n545) );
  NAND2_X1 U607 ( .A1(n550), .A2(n558), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U609 ( .A(n546), .B(G120GAT), .Z(G1341GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n548) );
  NAND2_X1 U611 ( .A1(n550), .A2(n583), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U613 ( .A(G127GAT), .B(n549), .Z(G1342GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n552) );
  NAND2_X1 U615 ( .A1(n550), .A2(n565), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U617 ( .A(G134GAT), .B(n553), .Z(G1343GAT) );
  XOR2_X1 U618 ( .A(G141GAT), .B(KEYINPUT121), .Z(n557) );
  NAND2_X1 U619 ( .A1(n554), .A2(n573), .ZN(n555) );
  XOR2_X1 U620 ( .A(KEYINPUT120), .B(n555), .Z(n566) );
  NAND2_X1 U621 ( .A1(n566), .A2(n568), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(G1344GAT) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT122), .ZN(n562) );
  XOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n560) );
  NAND2_X1 U625 ( .A1(n558), .A2(n566), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1345GAT) );
  XOR2_X1 U628 ( .A(G155GAT), .B(KEYINPUT123), .Z(n564) );
  NAND2_X1 U629 ( .A1(n583), .A2(n566), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1346GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n570), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n569), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U635 ( .A1(n570), .A2(n583), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U637 ( .A1(n572), .A2(n573), .ZN(n580) );
  NOR2_X1 U638 ( .A1(n574), .A2(n580), .ZN(n579) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n576) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(KEYINPUT59), .B(n577), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .Z(n582) );
  INV_X1 U645 ( .A(n580), .ZN(n586) );
  NAND2_X1 U646 ( .A1(n586), .A2(n372), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U648 ( .A1(n586), .A2(n583), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n590) );
  XOR2_X1 U651 ( .A(KEYINPUT127), .B(KEYINPUT126), .Z(n588) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(G1355GAT) );
endmodule

