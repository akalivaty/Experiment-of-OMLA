//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n613, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1120, new_n1121, new_n1122, new_n1123;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(KEYINPUT65), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n456), .A2(KEYINPUT65), .ZN(new_n458));
  NAND3_X1  g033(.A1(new_n455), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n463), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G137), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n466), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n468), .A2(G136), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT66), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n463), .A2(new_n466), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(G162));
  NAND2_X1  g055(.A1(new_n468), .A2(G138), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT4), .ZN(new_n482));
  NAND2_X1  g057(.A1(G114), .A2(G2104), .ZN(new_n483));
  INV_X1    g058(.A(G126), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n483), .B1(new_n463), .B2(new_n484), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n485), .A2(G2105), .B1(G102), .B2(new_n470), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G164));
  XNOR2_X1  g063(.A(KEYINPUT6), .B(G651), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G543), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G50), .ZN(new_n492));
  NAND2_X1  g067(.A1(G75), .A2(G543), .ZN(new_n493));
  INV_X1    g068(.A(G543), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT5), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G62), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n493), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n492), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT5), .B(G543), .ZN(new_n504));
  AND3_X1   g079(.A1(new_n489), .A2(new_n504), .A3(KEYINPUT67), .ZN(new_n505));
  AOI21_X1  g080(.A(KEYINPUT67), .B1(new_n489), .B2(new_n504), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n503), .B1(new_n507), .B2(G88), .ZN(G166));
  AND2_X1   g083(.A1(new_n507), .A2(G89), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT7), .ZN(new_n510));
  NAND2_X1  g085(.A1(G76), .A2(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(new_n502), .ZN(new_n512));
  XOR2_X1   g087(.A(KEYINPUT68), .B(G51), .Z(new_n513));
  NOR2_X1   g088(.A1(new_n511), .A2(new_n510), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n514), .B1(new_n504), .B2(G63), .ZN(new_n515));
  OAI221_X1 g090(.A(new_n512), .B1(new_n490), .B2(new_n513), .C1(new_n515), .C2(new_n502), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n509), .A2(new_n516), .ZN(G168));
  AOI22_X1  g092(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n520), .A2(new_n502), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n491), .A2(G52), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n502), .A2(KEYINPUT6), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT6), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G651), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n523), .A2(new_n525), .A3(new_n495), .A4(new_n497), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT67), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n489), .A2(new_n504), .A3(KEYINPUT67), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n522), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n521), .A2(new_n532), .ZN(G171));
  AOI22_X1  g108(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n502), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n491), .A2(G43), .ZN(new_n536));
  INV_X1    g111(.A(G81), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n538), .A2(new_n539), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n535), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G860), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n542), .A2(new_n543), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND3_X1  g120(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n546));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(KEYINPUT8), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n547), .A2(KEYINPUT8), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n546), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  XOR2_X1   g125(.A(new_n550), .B(KEYINPUT71), .Z(G188));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n552), .B1(new_n505), .B2(new_n506), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n528), .A2(KEYINPUT73), .A3(new_n529), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G91), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT72), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n491), .B2(G53), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n502), .ZN(new_n561));
  XOR2_X1   g136(.A(KEYINPUT72), .B(KEYINPUT9), .Z(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  NOR3_X1   g138(.A1(new_n490), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NOR3_X1   g139(.A1(new_n559), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n556), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  OAI21_X1  g144(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(new_n555), .B2(G87), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n491), .A2(G49), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT74), .ZN(new_n574));
  AND2_X1   g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G288));
  AOI22_X1  g151(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(G48), .B2(new_n491), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(G86), .B2(new_n555), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(new_n491), .A2(G47), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  OAI221_X1 g160(.A(new_n583), .B1(new_n502), .B2(new_n584), .C1(new_n530), .C2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT75), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n586), .B(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n528), .A2(KEYINPUT73), .A3(new_n529), .ZN(new_n590));
  AOI21_X1  g165(.A(KEYINPUT73), .B1(new_n528), .B2(new_n529), .ZN(new_n591));
  OAI21_X1  g166(.A(G92), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n498), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(G54), .A2(new_n491), .B1(new_n596), .B2(G651), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n555), .A2(new_n598), .A3(G92), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n593), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  XOR2_X1   g175(.A(new_n600), .B(KEYINPUT76), .Z(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n589), .B1(new_n602), .B2(G868), .ZN(G284));
  XOR2_X1   g178(.A(G284), .B(KEYINPUT77), .Z(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  XOR2_X1   g180(.A(G299), .B(KEYINPUT78), .Z(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G297));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(G148));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n542), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n601), .A2(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n611), .ZN(G323));
  XOR2_X1   g189(.A(G323), .B(KEYINPUT79), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n464), .A2(new_n470), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT82), .B(G2100), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT81), .B(KEYINPUT13), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n468), .A2(G135), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n478), .A2(G123), .ZN(new_n625));
  NOR2_X1   g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(new_n466), .B2(G111), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n624), .B(new_n625), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n623), .A2(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2435), .ZN(new_n632));
  XOR2_X1   g207(.A(G2427), .B(G2438), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(KEYINPUT14), .ZN(new_n635));
  XOR2_X1   g210(.A(G2443), .B(G2446), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n637), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n643), .A2(G14), .ZN(G401));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2067), .B(G2678), .Z(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n645), .B1(new_n649), .B2(KEYINPUT18), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2100), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(new_n648), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n649), .A2(new_n652), .A3(KEYINPUT17), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT18), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n651), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT84), .B(G2096), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G227));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  XOR2_X1   g235(.A(G1956), .B(G2474), .Z(new_n661));
  XOR2_X1   g236(.A(G1961), .B(G1966), .Z(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT20), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n661), .A2(new_n662), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n667), .A2(new_n660), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT85), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n667), .A2(new_n660), .A3(new_n663), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n665), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1991), .B(G1996), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT86), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G229));
  INV_X1    g253(.A(G29), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G26), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n478), .A2(G128), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT91), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n478), .A2(KEYINPUT91), .A3(G128), .ZN(new_n684));
  AOI22_X1  g259(.A1(new_n683), .A2(new_n684), .B1(G140), .B2(new_n468), .ZN(new_n685));
  OR2_X1    g260(.A1(G104), .A2(G2105), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n686), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n680), .B1(new_n689), .B2(new_n679), .ZN(new_n690));
  MUX2_X1   g265(.A(new_n680), .B(new_n690), .S(KEYINPUT28), .Z(new_n691));
  OR2_X1    g266(.A1(new_n691), .A2(G2067), .ZN(new_n692));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n575), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n693), .B2(G23), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT33), .Z(new_n696));
  INV_X1    g271(.A(G1976), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n695), .B(KEYINPUT33), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G1976), .ZN(new_n700));
  NOR2_X1   g275(.A1(G166), .A2(new_n693), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n693), .B2(G22), .ZN(new_n702));
  INV_X1    g277(.A(G1971), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n693), .A2(G6), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n581), .B2(new_n693), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT32), .B(G1981), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  NOR3_X1   g284(.A1(new_n704), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n702), .A2(new_n703), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n698), .A2(new_n700), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(KEYINPUT34), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT88), .ZN(new_n714));
  NOR2_X1   g289(.A1(G25), .A2(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n468), .A2(G131), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n478), .A2(G119), .ZN(new_n717));
  NOR2_X1   g292(.A1(G95), .A2(G2105), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(new_n466), .B2(G107), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n716), .B(new_n717), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT87), .Z(new_n721));
  AOI21_X1  g296(.A(new_n715), .B1(new_n721), .B2(G29), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT35), .B(G1991), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n722), .B(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n712), .A2(KEYINPUT34), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT89), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n693), .A2(G24), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n586), .B(KEYINPUT75), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n693), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1986), .ZN(new_n731));
  NOR3_X1   g306(.A1(new_n726), .A2(new_n727), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n714), .A2(new_n725), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT36), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n693), .A2(G21), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G168), .B2(new_n693), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT94), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(G1966), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n470), .A2(G103), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT25), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(new_n466), .ZN(new_n744));
  AOI211_X1 g319(.A(new_n742), .B(new_n744), .C1(G139), .C2(new_n468), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G29), .ZN(new_n746));
  OAI21_X1  g321(.A(KEYINPUT92), .B1(G29), .B2(G33), .ZN(new_n747));
  OR3_X1    g322(.A1(KEYINPUT92), .A2(G29), .A3(G33), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(G2072), .Z(new_n750));
  INV_X1    g325(.A(G2078), .ZN(new_n751));
  NOR2_X1   g326(.A1(G164), .A2(new_n679), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G27), .B2(new_n679), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n750), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  OR2_X1    g329(.A1(KEYINPUT24), .A2(G34), .ZN(new_n755));
  NAND2_X1  g330(.A1(KEYINPUT24), .A2(G34), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n755), .A2(new_n679), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G160), .B2(new_n679), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2084), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT27), .B(G1996), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT93), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n468), .A2(G141), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n478), .A2(G129), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n470), .A2(G105), .ZN(new_n764));
  NAND3_X1  g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT26), .Z(new_n766));
  NAND4_X1  g341(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n766), .ZN(new_n767));
  MUX2_X1   g342(.A(G32), .B(new_n767), .S(G29), .Z(new_n768));
  AOI21_X1  g343(.A(new_n759), .B1(new_n761), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n753), .A2(new_n751), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(G28), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(G28), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n772), .A2(new_n773), .A3(new_n679), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n774), .B1(new_n679), .B2(new_n628), .C1(new_n768), .C2(new_n761), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  AND4_X1   g351(.A1(new_n740), .A2(new_n754), .A3(new_n769), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n739), .A2(G1966), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT95), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT31), .B(G11), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n693), .A2(G5), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G171), .B2(new_n693), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT96), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1961), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n777), .A2(new_n779), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT97), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NOR2_X1   g363(.A1(G4), .A2(G16), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n602), .B2(G16), .ZN(new_n790));
  INV_X1    g365(.A(G1348), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n693), .A2(G19), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n542), .B2(G16), .ZN(new_n794));
  MUX2_X1   g369(.A(new_n793), .B(new_n794), .S(KEYINPUT90), .Z(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1341), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n679), .A2(G35), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G162), .B2(new_n679), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT29), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n799), .A2(G2090), .B1(new_n691), .B2(G2067), .ZN(new_n800));
  INV_X1    g375(.A(G299), .ZN(new_n801));
  OAI21_X1  g376(.A(KEYINPUT23), .B1(new_n801), .B2(new_n693), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n693), .A2(G20), .ZN(new_n803));
  MUX2_X1   g378(.A(new_n802), .B(KEYINPUT23), .S(new_n803), .Z(new_n804));
  OAI221_X1 g379(.A(new_n800), .B1(G1956), .B2(new_n804), .C1(G2090), .C2(new_n799), .ZN(new_n805));
  AOI211_X1 g380(.A(new_n796), .B(new_n805), .C1(G1956), .C2(new_n804), .ZN(new_n806));
  AND4_X1   g381(.A1(new_n787), .A2(new_n788), .A3(new_n792), .A4(new_n806), .ZN(new_n807));
  AND4_X1   g382(.A1(new_n692), .A2(new_n735), .A3(new_n736), .A4(new_n807), .ZN(G311));
  NAND4_X1  g383(.A1(new_n735), .A2(new_n692), .A3(new_n736), .A4(new_n807), .ZN(G150));
  NAND2_X1  g384(.A1(new_n491), .A2(G55), .ZN(new_n810));
  INV_X1    g385(.A(G93), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT99), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n504), .A2(G67), .ZN(new_n813));
  NAND2_X1  g388(.A1(G80), .A2(G543), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n812), .B1(new_n815), .B2(G651), .ZN(new_n816));
  AOI211_X1 g391(.A(KEYINPUT99), .B(new_n502), .C1(new_n813), .C2(new_n814), .ZN(new_n817));
  OAI221_X1 g392(.A(new_n810), .B1(new_n811), .B2(new_n530), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(G860), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT37), .Z(new_n820));
  INV_X1    g395(.A(KEYINPUT100), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n601), .A2(new_n609), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n818), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n542), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n818), .B(new_n535), .C1(new_n540), .C2(new_n541), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n824), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n821), .B1(new_n831), .B2(KEYINPUT39), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n830), .A2(KEYINPUT100), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n832), .A2(new_n543), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n830), .A2(new_n833), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n820), .B1(new_n835), .B2(new_n836), .ZN(G145));
  NAND2_X1  g412(.A1(new_n745), .A2(KEYINPUT101), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n688), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n720), .ZN(new_n840));
  XNOR2_X1  g415(.A(G160), .B(new_n628), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n619), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n840), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(G162), .B(new_n767), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n468), .A2(G142), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n478), .A2(G130), .ZN(new_n846));
  NOR2_X1   g421(.A1(G106), .A2(G2105), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(new_n466), .B2(G118), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n845), .B(new_n846), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n487), .B(new_n849), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n844), .B(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n843), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(G37), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT40), .Z(G395));
  NAND2_X1  g430(.A1(new_n818), .A2(new_n611), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n828), .B(KEYINPUT102), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(new_n613), .Z(new_n858));
  INV_X1    g433(.A(KEYINPUT104), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n598), .B1(new_n555), .B2(G92), .ZN(new_n860));
  INV_X1    g435(.A(G92), .ZN(new_n861));
  AOI211_X1 g436(.A(KEYINPUT10), .B(new_n861), .C1(new_n553), .C2(new_n554), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  OR3_X1    g438(.A1(new_n559), .A2(new_n561), .A3(new_n564), .ZN(new_n864));
  INV_X1    g439(.A(G91), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(new_n553), .B2(new_n554), .ZN(new_n866));
  OAI21_X1  g441(.A(KEYINPUT103), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n556), .A2(new_n868), .A3(new_n565), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n863), .A2(new_n867), .A3(new_n597), .A4(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n600), .A2(KEYINPUT103), .A3(G299), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT41), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT41), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n870), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n859), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT104), .B1(new_n872), .B2(KEYINPUT41), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n858), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n872), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n879), .B1(new_n880), .B2(new_n858), .ZN(new_n881));
  NAND2_X1  g456(.A1(G290), .A2(G166), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n729), .A2(G303), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n882), .A2(new_n883), .A3(G305), .ZN(new_n884));
  AOI21_X1  g459(.A(G305), .B1(new_n882), .B2(new_n883), .ZN(new_n885));
  OAI21_X1  g460(.A(G288), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(new_n883), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n581), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n882), .A2(new_n883), .A3(G305), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n575), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT42), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n881), .B(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n856), .B1(new_n893), .B2(new_n611), .ZN(G295));
  OAI21_X1  g469(.A(new_n856), .B1(new_n893), .B2(new_n611), .ZN(G331));
  XNOR2_X1  g470(.A(G171), .B(G168), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(new_n827), .A3(new_n826), .ZN(new_n897));
  XNOR2_X1  g472(.A(G286), .B(G171), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n828), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n876), .B2(new_n877), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n897), .A2(new_n899), .A3(KEYINPUT106), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(KEYINPUT106), .B2(new_n897), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n880), .ZN(new_n906));
  OAI211_X1 g481(.A(KEYINPUT105), .B(new_n900), .C1(new_n876), .C2(new_n877), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n903), .A2(KEYINPUT107), .A3(new_n906), .A4(new_n907), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n886), .A2(new_n890), .A3(KEYINPUT108), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT108), .B1(new_n886), .B2(new_n890), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n910), .A2(new_n911), .A3(new_n915), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n903), .A2(new_n891), .A3(new_n906), .A4(new_n907), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n853), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n921), .A3(KEYINPUT43), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n914), .B1(new_n908), .B2(new_n909), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n918), .B1(new_n923), .B2(new_n911), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT109), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n873), .A2(new_n875), .ZN(new_n927));
  OAI22_X1  g502(.A1(new_n905), .A2(new_n927), .B1(new_n872), .B2(new_n900), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n918), .B1(new_n915), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n925), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n922), .A2(new_n926), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(KEYINPUT43), .B2(new_n924), .ZN(new_n933));
  MUX2_X1   g508(.A(new_n931), .B(new_n933), .S(KEYINPUT44), .Z(G397));
  AOI21_X1  g509(.A(G1384), .B1(new_n482), .B2(new_n486), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n935), .A2(KEYINPUT45), .ZN(new_n936));
  AND2_X1   g511(.A1(G160), .A2(G40), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G1996), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT125), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT46), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n941), .B(new_n943), .Z(new_n944));
  INV_X1    g519(.A(G2067), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n688), .B(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n939), .B1(new_n947), .B2(new_n767), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT126), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n944), .B(new_n949), .C1(new_n942), .C2(KEYINPUT46), .ZN(new_n950));
  XOR2_X1   g525(.A(new_n950), .B(KEYINPUT47), .Z(new_n951));
  INV_X1    g526(.A(new_n939), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n952), .A2(G1986), .A3(G290), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT48), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n767), .B(G1996), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n947), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n720), .B(new_n724), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n954), .B1(new_n939), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n724), .A3(new_n721), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n689), .A2(new_n945), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n952), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n951), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n937), .A2(new_n935), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n964), .A2(G8), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n575), .A2(G1976), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n967), .A2(KEYINPUT112), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(KEYINPUT112), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n969), .A3(KEYINPUT52), .ZN(new_n970));
  OR2_X1    g545(.A1(G305), .A2(G1981), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n507), .A2(G86), .ZN(new_n972));
  OAI21_X1  g547(.A(G1981), .B1(new_n580), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT49), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n965), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n965), .A2(new_n977), .A3(new_n966), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT113), .B(G1976), .Z(new_n979));
  AND2_X1   g554(.A1(G288), .A2(new_n979), .ZN(new_n980));
  OR3_X1    g555(.A1(new_n978), .A2(KEYINPUT114), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT114), .B1(new_n978), .B2(new_n980), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n970), .A2(new_n976), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(G303), .A2(G8), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT55), .ZN(new_n986));
  XOR2_X1   g561(.A(new_n986), .B(KEYINPUT111), .Z(new_n987));
  NAND2_X1  g562(.A1(new_n935), .A2(KEYINPUT45), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n936), .A2(new_n937), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n703), .ZN(new_n990));
  INV_X1    g565(.A(G1384), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n487), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT50), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n938), .B1(new_n993), .B2(KEYINPUT110), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n935), .A2(new_n995), .ZN(new_n996));
  OR3_X1    g571(.A1(new_n935), .A2(KEYINPUT110), .A3(new_n995), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n990), .B1(new_n998), .B2(G2090), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n987), .A2(G8), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n993), .A2(new_n937), .A3(new_n996), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n990), .B1(G2090), .B2(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1002), .A2(KEYINPUT115), .ZN(new_n1003));
  OAI21_X1  g578(.A(G8), .B1(new_n1002), .B2(KEYINPUT115), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n986), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n984), .A2(new_n1000), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n989), .ZN(new_n1007));
  OAI22_X1  g582(.A1(new_n998), .A2(G2084), .B1(new_n1007), .B2(G1966), .ZN(new_n1008));
  OAI21_X1  g583(.A(G8), .B1(new_n1008), .B2(G286), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(KEYINPUT51), .B(G8), .C1(new_n1008), .C2(G286), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(KEYINPUT120), .A3(new_n1012), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1008), .A2(G8), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G286), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1009), .A2(new_n1016), .A3(new_n1010), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1013), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT62), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(KEYINPUT124), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1013), .A2(new_n1020), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1961), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n998), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n989), .A2(G2078), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT53), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n989), .B2(G2078), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G171), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(KEYINPUT124), .B2(new_n1019), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1024), .A2(new_n1033), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1025), .A2(new_n998), .B1(new_n1027), .B2(KEYINPUT53), .ZN(new_n1035));
  AOI21_X1  g610(.A(G301), .B1(new_n1035), .B2(new_n1030), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT122), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT54), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1031), .A2(new_n1037), .A3(G171), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1035), .A2(G301), .A3(new_n1030), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT123), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1038), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  AND4_X1   g618(.A1(G301), .A2(new_n1026), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1046), .B1(new_n1032), .B2(KEYINPUT122), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT123), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1043), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n998), .A2(new_n791), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n964), .B(KEYINPUT119), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n945), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n600), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT118), .B(G1956), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1001), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(G299), .B(KEYINPUT57), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT56), .B(G2072), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1007), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1057), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1053), .A2(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1007), .A2(new_n1060), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1058), .B1(new_n1064), .B2(new_n1056), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1050), .A2(new_n600), .A3(new_n1052), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT60), .B1(new_n1066), .B2(new_n1053), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT61), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1064), .A2(new_n1058), .A3(new_n1056), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1059), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1065), .A2(new_n1062), .A3(KEYINPUT61), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n600), .A2(KEYINPUT60), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1050), .A2(new_n1052), .A3(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1067), .A2(new_n1071), .A3(new_n1072), .A4(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT58), .B(G1341), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1051), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1007), .A2(new_n940), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n542), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n1079), .B(KEYINPUT59), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1063), .B(new_n1065), .C1(new_n1075), .C2(new_n1080), .ZN(new_n1081));
  XOR2_X1   g656(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(new_n1036), .B2(new_n1044), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1049), .A2(new_n1018), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1006), .B1(new_n1034), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT63), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1014), .A2(G168), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n1006), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n999), .A2(new_n1090), .A3(G8), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1090), .B1(new_n999), .B2(G8), .ZN(new_n1093));
  INV_X1    g668(.A(new_n986), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n970), .A2(new_n976), .A3(new_n983), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1089), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1087), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1093), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(new_n986), .A3(new_n1091), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1100), .A2(new_n984), .A3(KEYINPUT117), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1097), .A2(new_n1000), .A3(new_n1098), .A4(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1088), .B1(new_n1102), .B2(new_n1086), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n976), .A2(new_n697), .A3(new_n575), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n971), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n965), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1096), .A2(new_n1000), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1085), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n958), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n729), .B(G1986), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n952), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n963), .B1(new_n1109), .B2(new_n1112), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g688(.A1(G227), .A2(new_n459), .ZN(new_n1115));
  NOR4_X1   g689(.A1(new_n854), .A2(G401), .A3(G229), .A4(new_n1115), .ZN(new_n1116));
  AND3_X1   g690(.A1(new_n931), .A2(KEYINPUT127), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g691(.A(KEYINPUT127), .B1(new_n931), .B2(new_n1116), .ZN(new_n1118));
  NOR2_X1   g692(.A1(new_n1117), .A2(new_n1118), .ZN(G308));
  NAND2_X1  g693(.A1(new_n931), .A2(new_n1116), .ZN(new_n1120));
  INV_X1    g694(.A(KEYINPUT127), .ZN(new_n1121));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g696(.A1(new_n931), .A2(KEYINPUT127), .A3(new_n1116), .ZN(new_n1123));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n1123), .ZN(G225));
endmodule


