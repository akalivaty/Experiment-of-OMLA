//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967;
  INV_X1    g000(.A(G113gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G120gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n203), .B(KEYINPUT71), .Z(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT70), .B(G120gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G113gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G127gat), .B(G134gat), .Z(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n211));
  INV_X1    g010(.A(G120gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G113gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n203), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n211), .B1(new_n214), .B2(KEYINPUT68), .ZN(new_n215));
  XNOR2_X1  g014(.A(G113gat), .B(G120gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n208), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(KEYINPUT69), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT69), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT1), .B1(new_n216), .B2(new_n217), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n214), .A2(KEYINPUT68), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n221), .B1(new_n224), .B2(new_n208), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n210), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G148gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G141gat), .ZN(new_n228));
  INV_X1    g027(.A(G141gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G148gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT77), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT2), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n233), .A2(KEYINPUT78), .B1(G155gat), .B2(G162gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(KEYINPUT78), .B2(new_n233), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT77), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n228), .A2(new_n230), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  XOR2_X1   g037(.A(G155gat), .B(G162gat), .Z(new_n239));
  NAND2_X1  g038(.A1(new_n229), .A2(KEYINPUT79), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT79), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G141gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n242), .A3(G148gat), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n239), .B1(new_n228), .B2(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(KEYINPUT80), .B(G162gat), .Z(new_n245));
  INV_X1    g044(.A(G155gat), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT2), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n238), .A2(new_n239), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n226), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G225gat), .A2(G233gat), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n248), .B(new_n210), .C1(new_n220), .C2(new_n225), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT85), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n252), .A2(KEYINPUT4), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n239), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n244), .A2(new_n247), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n258), .B1(new_n256), .B2(new_n257), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n226), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n219), .A2(KEYINPUT69), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n224), .A2(new_n221), .A3(new_n208), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n264), .A2(new_n265), .B1(new_n207), .B2(new_n209), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n263), .B1(new_n266), .B2(new_n248), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n255), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n251), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n254), .A2(KEYINPUT39), .A3(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G1gat), .B(G29gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(KEYINPUT0), .ZN(new_n273));
  XNOR2_X1  g072(.A(G57gat), .B(G85gat), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n273), .B(new_n274), .Z(new_n275));
  OAI211_X1 g074(.A(new_n271), .B(new_n275), .C1(KEYINPUT39), .C2(new_n270), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT40), .ZN(new_n277));
  XOR2_X1   g076(.A(G8gat), .B(G36gat), .Z(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT75), .ZN(new_n279));
  XNOR2_X1  g078(.A(G64gat), .B(G92gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT25), .ZN(new_n283));
  INV_X1    g082(.A(G190gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(G183gat), .ZN(new_n285));
  INV_X1    g084(.A(G183gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(G190gat), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT24), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  OR3_X1    g087(.A1(new_n286), .A2(new_n284), .A3(KEYINPUT24), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT23), .ZN(new_n290));
  INV_X1    g089(.A(G169gat), .ZN(new_n291));
  INV_X1    g090(.A(G176gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n293), .A2(new_n294), .B1(G169gat), .B2(G176gat), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n288), .B(new_n289), .C1(new_n295), .C2(KEYINPUT64), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n295), .A2(KEYINPUT64), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n283), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT65), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT65), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n300), .B(new_n283), .C1(new_n296), .C2(new_n297), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n293), .A2(new_n294), .ZN(new_n302));
  NAND2_X1  g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT66), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n283), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n302), .B(new_n305), .C1(new_n304), .C2(new_n303), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n288), .A2(new_n289), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n299), .A2(new_n301), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT27), .B(G183gat), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT67), .B1(new_n311), .B2(new_n284), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n312), .A2(KEYINPUT28), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(KEYINPUT28), .ZN(new_n314));
  NOR3_X1   g113(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT26), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n303), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI22_X1  g117(.A1(new_n315), .A2(new_n318), .B1(new_n286), .B2(new_n284), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n313), .A2(new_n314), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n310), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(G226gat), .A3(G233gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(G226gat), .A2(G233gat), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n308), .B1(new_n298), .B2(KEYINPUT65), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n320), .B1(new_n325), .B2(new_n301), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n324), .B1(new_n326), .B2(KEYINPUT29), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G197gat), .ZN(new_n329));
  INV_X1    g128(.A(G204gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(G197gat), .A2(G204gat), .ZN(new_n332));
  AND2_X1   g131(.A1(G211gat), .A2(G218gat), .ZN(new_n333));
  OAI22_X1  g132(.A1(new_n331), .A2(new_n332), .B1(KEYINPUT22), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT74), .ZN(new_n335));
  NOR2_X1   g134(.A1(G211gat), .A2(G218gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n337), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n334), .A2(new_n339), .A3(KEYINPUT74), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n328), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n323), .A2(new_n327), .A3(new_n341), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n282), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT76), .B1(new_n345), .B2(KEYINPUT30), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n323), .A2(new_n327), .A3(new_n341), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n341), .B1(new_n323), .B2(new_n327), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n281), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT30), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g152(.A(KEYINPUT30), .B(new_n281), .C1(new_n347), .C2(new_n348), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n343), .A2(new_n282), .A3(new_n344), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n359), .B1(new_n268), .B2(new_n269), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n266), .A2(new_n263), .A3(new_n248), .ZN(new_n361));
  NOR3_X1   g160(.A1(new_n266), .A2(new_n259), .A3(new_n260), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n252), .A2(KEYINPUT4), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(KEYINPUT81), .A3(new_n251), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n266), .A2(new_n248), .ZN(new_n366));
  INV_X1    g165(.A(new_n252), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n269), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT82), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n369), .A3(KEYINPUT5), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n251), .B1(new_n250), .B2(new_n252), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT5), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT82), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n360), .A2(new_n365), .A3(new_n370), .A4(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n364), .A2(new_n372), .A3(new_n251), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n275), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n277), .A2(new_n358), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT84), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n341), .B1(new_n259), .B2(KEYINPUT29), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n334), .A2(new_n339), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT29), .B1(new_n334), .B2(new_n339), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(KEYINPUT83), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n258), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT83), .B1(new_n381), .B2(new_n382), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n249), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G228gat), .A2(G233gat), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n258), .B1(new_n341), .B2(KEYINPUT29), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n388), .B1(new_n389), .B2(new_n249), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n387), .A2(new_n388), .B1(new_n390), .B2(new_n380), .ZN(new_n391));
  XNOR2_X1  g190(.A(G78gat), .B(G106gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(KEYINPUT31), .B(G50gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n392), .B(new_n393), .Z(new_n394));
  OAI21_X1  g193(.A(new_n379), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(G22gat), .ZN(new_n396));
  INV_X1    g195(.A(G22gat), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n379), .B(new_n397), .C1(new_n391), .C2(new_n394), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n391), .A2(new_n394), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n396), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n396), .B2(new_n398), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n365), .A2(new_n370), .A3(new_n373), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT81), .B1(new_n364), .B2(new_n251), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n375), .B(new_n275), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT6), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(new_n376), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI211_X1 g208(.A(new_n406), .B(new_n275), .C1(new_n374), .C2(new_n375), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT37), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT37), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n414), .B1(new_n343), .B2(new_n344), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n282), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n345), .B1(new_n416), .B2(KEYINPUT38), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n417), .B1(KEYINPUT38), .B2(new_n416), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n378), .B(new_n402), .C1(new_n412), .C2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT72), .ZN(new_n420));
  XNOR2_X1  g219(.A(G15gat), .B(G43gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(G71gat), .B(G99gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n310), .A2(new_n226), .A3(new_n321), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n226), .B1(new_n310), .B2(new_n321), .ZN(new_n426));
  NAND2_X1  g225(.A1(G227gat), .A2(G233gat), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT32), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n424), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n428), .A2(KEYINPUT33), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n420), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n426), .ZN(new_n433));
  INV_X1    g232(.A(new_n427), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n326), .A2(new_n226), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT32), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT33), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n437), .A2(new_n439), .A3(KEYINPUT72), .A4(new_n424), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n432), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n423), .A2(new_n438), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n427), .B1(new_n425), .B2(new_n426), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT34), .B1(new_n434), .B2(KEYINPUT73), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n446), .B(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n449), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n441), .A2(new_n451), .A3(new_n444), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(KEYINPUT36), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT36), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n451), .B1(new_n441), .B2(new_n444), .ZN(new_n455));
  AOI211_X1 g254(.A(new_n443), .B(new_n449), .C1(new_n432), .C2(new_n440), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n356), .B1(new_n346), .B2(new_n352), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(new_n408), .B2(new_n410), .ZN(new_n460));
  INV_X1    g259(.A(new_n402), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n419), .A2(new_n458), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n450), .A2(new_n402), .A3(new_n452), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT35), .B1(new_n464), .B2(new_n460), .ZN(new_n465));
  NOR3_X1   g264(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT35), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n459), .B(new_n466), .C1(new_n408), .C2(new_n410), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n450), .A2(KEYINPUT86), .A3(new_n452), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT86), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n469), .B1(new_n455), .B2(new_n456), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n467), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n465), .B1(new_n471), .B2(KEYINPUT87), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT87), .ZN(new_n473));
  AOI211_X1 g272(.A(new_n473), .B(new_n467), .C1(new_n468), .C2(new_n470), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n463), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G113gat), .B(G141gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(G197gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT11), .B(G169gat), .ZN(new_n478));
  XOR2_X1   g277(.A(new_n477), .B(new_n478), .Z(new_n479));
  XNOR2_X1  g278(.A(new_n479), .B(KEYINPUT12), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G29gat), .ZN(new_n482));
  INV_X1    g281(.A(G36gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AND2_X1   g283(.A1(KEYINPUT88), .A2(KEYINPUT14), .ZN(new_n485));
  NOR2_X1   g284(.A1(KEYINPUT88), .A2(KEYINPUT14), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(KEYINPUT88), .A2(KEYINPUT14), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(new_n482), .A3(new_n483), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(G29gat), .A2(G36gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G50gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(G43gat), .ZN(new_n494));
  INV_X1    g293(.A(G43gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(G50gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n496), .A3(KEYINPUT15), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT91), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n487), .A2(new_n500), .A3(new_n489), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n500), .B1(new_n487), .B2(new_n489), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT90), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n493), .B2(G43gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n495), .A2(KEYINPUT90), .A3(G50gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n494), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n497), .A2(KEYINPUT89), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n494), .A2(new_n496), .A3(new_n511), .A4(KEYINPUT15), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n509), .A2(new_n491), .A3(new_n510), .A4(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n499), .B1(new_n503), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT92), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT17), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT92), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n517), .B(new_n499), .C1(new_n503), .C2(new_n513), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT93), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n515), .A2(KEYINPUT93), .A3(new_n516), .A4(new_n518), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n524), .A2(G1gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT16), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n524), .B1(new_n526), .B2(G1gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n527), .A3(KEYINPUT94), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n528), .B(G8gat), .C1(KEYINPUT94), .C2(new_n527), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n527), .A2(KEYINPUT95), .ZN(new_n530));
  INV_X1    g329(.A(G8gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n527), .A2(KEYINPUT95), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n525), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  OR3_X1    g333(.A1(new_n514), .A2(KEYINPUT96), .A3(new_n516), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT96), .B1(new_n514), .B2(new_n516), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n523), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n515), .A2(new_n534), .A3(new_n518), .ZN(new_n539));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT18), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n538), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n540), .B(KEYINPUT13), .Z(new_n545));
  INV_X1    g344(.A(new_n539), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n534), .B1(new_n515), .B2(new_n518), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n546), .B1(new_n523), .B2(new_n537), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT18), .B1(new_n550), .B2(new_n540), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n481), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n548), .A2(new_n480), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n544), .A2(new_n554), .ZN(new_n555));
  NOR3_X1   g354(.A1(new_n555), .A2(new_n551), .A3(KEYINPUT97), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n538), .A2(new_n540), .A3(new_n539), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(new_n542), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n553), .B1(new_n550), .B2(new_n543), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n552), .B1(new_n556), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n475), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT98), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT98), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n475), .A2(new_n565), .A3(new_n562), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT9), .ZN(new_n568));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n568), .B1(new_n569), .B2(KEYINPUT99), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n570), .B1(KEYINPUT99), .B2(new_n569), .ZN(new_n571));
  XOR2_X1   g370(.A(G71gat), .B(G78gat), .Z(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n569), .B(KEYINPUT100), .ZN(new_n574));
  INV_X1    g373(.A(G71gat), .ZN(new_n575));
  INV_X1    g374(.A(G78gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n576), .A3(KEYINPUT9), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n577), .B1(new_n575), .B2(new_n576), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n581), .A2(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(G127gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n534), .B1(KEYINPUT21), .B2(new_n581), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(G155gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(G183gat), .B(G211gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n588), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n596), .B(KEYINPUT101), .Z(new_n597));
  INV_X1    g396(.A(KEYINPUT41), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT102), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(G85gat), .A3(G92gat), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT7), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n602), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n605), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G99gat), .B(G106gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n515), .A2(new_n518), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(new_n598), .B2(new_n597), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n613), .B1(new_n535), .B2(new_n536), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n615), .B1(new_n523), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G190gat), .B(G218gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  AOI211_X1 g419(.A(new_n618), .B(new_n615), .C1(new_n523), .C2(new_n616), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n601), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT103), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI211_X1 g423(.A(KEYINPUT103), .B(new_n601), .C1(new_n620), .C2(new_n621), .ZN(new_n625));
  OR3_X1    g424(.A1(new_n617), .A2(KEYINPUT104), .A3(new_n619), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n621), .A2(new_n601), .ZN(new_n627));
  OAI21_X1  g426(.A(KEYINPUT104), .B1(new_n617), .B2(new_n619), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n624), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n595), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G120gat), .B(G148gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(G176gat), .B(G204gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n633), .B(new_n634), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n611), .B(new_n612), .Z(new_n637));
  NAND2_X1  g436(.A1(new_n580), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n613), .A2(new_n579), .A3(new_n573), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n581), .A2(KEYINPUT10), .A3(new_n613), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n644), .B1(new_n638), .B2(new_n640), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n636), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n636), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n645), .B(new_n650), .C1(new_n649), .C2(new_n647), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n632), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n412), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT106), .B1(new_n409), .B2(new_n411), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n567), .A2(new_n653), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G1gat), .ZN(G1324gat));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n475), .A2(new_n565), .A3(new_n562), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n565), .B1(new_n475), .B2(new_n562), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n358), .B(new_n653), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT16), .B(G8gat), .Z(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n660), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT107), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OR3_X1    g467(.A1(new_n663), .A2(new_n660), .A3(new_n665), .ZN(new_n669));
  OAI211_X1 g468(.A(KEYINPUT107), .B(new_n660), .C1(new_n663), .C2(new_n665), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n663), .A2(G8gat), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n668), .A2(new_n669), .A3(new_n670), .A4(new_n671), .ZN(G1325gat));
  NAND2_X1  g471(.A1(new_n567), .A2(new_n653), .ZN(new_n673));
  OAI21_X1  g472(.A(G15gat), .B1(new_n673), .B2(new_n458), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n468), .A2(new_n470), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n675), .A2(G15gat), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n674), .B1(new_n673), .B2(new_n676), .ZN(G1326gat));
  NAND3_X1  g476(.A1(new_n567), .A2(new_n461), .A3(new_n653), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT43), .B(G22gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  INV_X1    g479(.A(new_n595), .ZN(new_n681));
  INV_X1    g480(.A(new_n652), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n631), .ZN(new_n684));
  INV_X1    g483(.A(new_n657), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(G29gat), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n684), .B(new_n686), .C1(new_n661), .C2(new_n662), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT108), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT108), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n567), .A2(new_n689), .A3(new_n684), .A4(new_n686), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT45), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n691), .B1(new_n688), .B2(new_n690), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n475), .A2(new_n630), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n475), .A2(KEYINPUT44), .A3(new_n630), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n562), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT109), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n698), .A2(new_n657), .A3(new_n701), .ZN(new_n702));
  OAI22_X1  g501(.A1(new_n692), .A2(new_n693), .B1(new_n482), .B2(new_n702), .ZN(G1328gat));
  INV_X1    g502(.A(new_n684), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n704), .B1(new_n564), .B2(new_n566), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(new_n483), .A3(new_n358), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n706), .A2(KEYINPUT46), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n698), .A2(new_n358), .A3(new_n701), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G36gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n706), .A2(KEYINPUT46), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n707), .A2(new_n709), .A3(new_n710), .ZN(G1329gat));
  INV_X1    g510(.A(new_n675), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n712), .B(new_n684), .C1(new_n661), .C2(new_n662), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n495), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n458), .A2(new_n495), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n696), .A2(new_n697), .A3(new_n701), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT111), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n714), .A2(new_n716), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT47), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n714), .A2(new_n722), .A3(new_n716), .A4(new_n717), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n719), .A2(new_n721), .A3(new_n723), .ZN(G1330gat));
  NAND3_X1  g523(.A1(new_n705), .A2(new_n493), .A3(new_n461), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n696), .A2(new_n461), .A3(new_n697), .A4(new_n701), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G50gat), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n725), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n726), .B1(new_n725), .B2(new_n728), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(G1331gat));
  NOR3_X1   g530(.A1(new_n632), .A2(new_n562), .A3(new_n682), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n475), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n657), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n358), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT49), .B(G64gat), .Z(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT112), .ZN(G1333gat));
  NAND2_X1  g539(.A1(new_n733), .A2(new_n712), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n575), .ZN(new_n742));
  INV_X1    g541(.A(new_n458), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n733), .A2(G71gat), .A3(new_n743), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n744), .A2(KEYINPUT113), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(KEYINPUT113), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n742), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT50), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n749), .B(new_n742), .C1(new_n745), .C2(new_n746), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(G1334gat));
  NAND2_X1  g550(.A1(new_n733), .A2(new_n461), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G78gat), .ZN(G1335gat));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(KEYINPUT115), .ZN(new_n755));
  INV_X1    g554(.A(new_n694), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n681), .A2(new_n699), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT114), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n755), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n694), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n763), .A2(new_n607), .A3(new_n652), .A4(new_n657), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n758), .A2(new_n682), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n698), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G85gat), .B1(new_n766), .B2(new_n685), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n767), .ZN(G1336gat));
  NOR3_X1   g567(.A1(new_n459), .A2(G92gat), .A3(new_n682), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n760), .B2(new_n762), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n696), .A2(new_n358), .A3(new_n697), .A4(new_n765), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G92gat), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n770), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT52), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n770), .A2(new_n772), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(G1337gat));
  OAI21_X1  g577(.A(G99gat), .B1(new_n766), .B2(new_n458), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n675), .A2(G99gat), .A3(new_n682), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(G1338gat));
  NOR3_X1   g581(.A1(new_n402), .A2(G106gat), .A3(new_n682), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(new_n760), .B2(new_n762), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n696), .A2(new_n461), .A3(new_n697), .A4(new_n765), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G106gat), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT53), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n784), .A2(new_n786), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(G1339gat));
  NAND4_X1  g591(.A1(new_n595), .A2(new_n699), .A3(new_n631), .A4(new_n682), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n636), .B1(new_n645), .B2(KEYINPUT54), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n641), .A2(G230gat), .A3(G233gat), .A4(new_n642), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n645), .A2(KEYINPUT54), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT118), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n643), .B2(new_n644), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(KEYINPUT118), .A3(new_n795), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n794), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n651), .B1(new_n802), .B2(KEYINPUT55), .ZN(new_n803));
  INV_X1    g602(.A(new_n794), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n800), .A2(KEYINPUT118), .A3(new_n795), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT118), .B1(new_n800), .B2(new_n795), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n803), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n479), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n538), .A2(new_n539), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n541), .ZN(new_n813));
  OR3_X1    g612(.A1(new_n546), .A2(new_n547), .A3(new_n545), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n811), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT97), .B1(new_n555), .B2(new_n551), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n559), .A2(new_n557), .A3(new_n560), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n630), .A2(new_n810), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n813), .A2(new_n814), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n479), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n652), .B(new_n822), .C1(new_n556), .C2(new_n561), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n818), .A2(KEYINPUT119), .A3(new_n652), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n562), .A2(new_n810), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n820), .B1(new_n828), .B2(new_n631), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n793), .B1(new_n829), .B2(new_n595), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n830), .A2(new_n402), .A3(new_n712), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n459), .A3(new_n657), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n832), .A2(new_n202), .A3(new_n699), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n830), .A2(new_n657), .ZN(new_n834));
  INV_X1    g633(.A(new_n464), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n459), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n562), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n833), .B1(new_n838), .B2(new_n202), .ZN(G1340gat));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n205), .A3(new_n652), .ZN(new_n840));
  OAI21_X1  g639(.A(G120gat), .B1(new_n832), .B2(new_n682), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1341gat));
  NAND3_X1  g641(.A1(new_n837), .A2(new_n585), .A3(new_n595), .ZN(new_n843));
  OAI21_X1  g642(.A(G127gat), .B1(new_n832), .B2(new_n681), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(G1342gat));
  NOR3_X1   g644(.A1(new_n631), .A2(new_n358), .A3(G134gat), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n836), .A2(new_n846), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n847), .A2(KEYINPUT56), .ZN(new_n848));
  OAI21_X1  g647(.A(G134gat), .B1(new_n832), .B2(new_n631), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(KEYINPUT56), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(G1343gat));
  NAND4_X1  g650(.A1(new_n834), .A2(new_n461), .A3(new_n459), .A4(new_n458), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n229), .A3(new_n562), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n240), .A2(new_n242), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n830), .A2(new_n856), .A3(new_n461), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n685), .A2(new_n743), .A3(new_n358), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n807), .A2(new_n808), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n802), .A2(KEYINPUT55), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n860), .A3(new_n651), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n816), .A2(new_n817), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(new_n552), .ZN(new_n863));
  INV_X1    g662(.A(new_n823), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT120), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n827), .A2(new_n866), .A3(new_n823), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n630), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n681), .B1(new_n868), .B2(new_n820), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n402), .B1(new_n869), .B2(new_n793), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n857), .B(new_n858), .C1(new_n870), .C2(new_n856), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n855), .B1(new_n871), .B2(new_n699), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n854), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n227), .A2(KEYINPUT59), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n875), .B(new_n876), .C1(new_n871), .C2(new_n682), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n827), .A2(new_n866), .A3(new_n823), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n866), .B1(new_n827), .B2(new_n823), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n631), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n595), .B1(new_n881), .B2(new_n819), .ZN(new_n882));
  INV_X1    g681(.A(new_n793), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n461), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT57), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n885), .A2(new_n652), .A3(new_n857), .A4(new_n858), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n875), .B1(new_n886), .B2(new_n876), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n830), .A2(new_n461), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT57), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n402), .A2(KEYINPUT57), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n892), .B1(new_n631), .B2(new_n861), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n630), .A2(new_n810), .A3(KEYINPUT122), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(new_n818), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n595), .B1(new_n881), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n891), .B1(new_n896), .B2(new_n883), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n890), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n858), .A2(new_n652), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n227), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI22_X1  g699(.A1(new_n878), .A2(new_n887), .B1(new_n888), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n853), .A2(new_n227), .A3(new_n652), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1345gat));
  NAND3_X1  g702(.A1(new_n853), .A2(new_n246), .A3(new_n595), .ZN(new_n904));
  OAI21_X1  g703(.A(G155gat), .B1(new_n871), .B2(new_n681), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1346gat));
  OR3_X1    g705(.A1(new_n871), .A2(KEYINPUT123), .A3(new_n631), .ZN(new_n907));
  INV_X1    g706(.A(new_n245), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT123), .B1(new_n871), .B2(new_n631), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n853), .A2(new_n245), .A3(new_n630), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1347gat));
  NOR2_X1   g711(.A1(new_n657), .A2(new_n459), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n831), .A2(new_n913), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n914), .A2(new_n291), .A3(new_n699), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n830), .A2(new_n685), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n464), .A2(new_n459), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(new_n562), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n915), .B1(new_n291), .B2(new_n918), .ZN(G1348gat));
  OAI21_X1  g718(.A(G176gat), .B1(new_n914), .B2(new_n682), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n916), .A2(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n652), .A2(new_n292), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(G1349gat));
  OAI21_X1  g722(.A(G183gat), .B1(new_n914), .B2(new_n681), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n595), .A2(new_n311), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT60), .ZN(G1350gat));
  NOR3_X1   g726(.A1(new_n921), .A2(G190gat), .A3(new_n631), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n831), .A2(new_n630), .A3(new_n913), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n930), .B2(G190gat), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n930), .A2(new_n929), .A3(G190gat), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(G1351gat));
  NOR3_X1   g735(.A1(new_n743), .A2(new_n402), .A3(new_n459), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n916), .A2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(G197gat), .B1(new_n939), .B2(new_n562), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n657), .A2(new_n743), .A3(new_n459), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n890), .A2(new_n897), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n699), .A2(new_n329), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(G1352gat));
  NAND4_X1  g743(.A1(new_n916), .A2(new_n330), .A3(new_n652), .A4(new_n937), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n945), .B(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n942), .A2(new_n652), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n947), .B(new_n948), .C1(new_n949), .C2(new_n330), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n945), .B(KEYINPUT62), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n330), .B1(new_n942), .B2(new_n652), .ZN(new_n952));
  OAI21_X1  g751(.A(KEYINPUT125), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n950), .A2(new_n953), .ZN(G1353gat));
  INV_X1    g753(.A(G211gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n955), .A3(new_n595), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n890), .A2(new_n897), .A3(new_n595), .A4(new_n941), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n957), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT63), .B1(new_n957), .B2(G211gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(KEYINPUT126), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n962), .B(new_n956), .C1(new_n958), .C2(new_n959), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n961), .A2(new_n963), .ZN(G1354gat));
  AOI21_X1  g763(.A(G218gat), .B1(new_n939), .B2(new_n630), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n630), .A2(G218gat), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT127), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n965), .B1(new_n942), .B2(new_n967), .ZN(G1355gat));
endmodule


