//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT64), .Z(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT65), .Z(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n209), .B1(new_n213), .B2(new_n215), .C1(new_n222), .C2(KEYINPUT1), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0024(.A(G250), .B(G257), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT66), .ZN(new_n226));
  XOR2_X1   g0026(.A(G264), .B(G270), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n228), .B(new_n232), .Z(G358));
  XOR2_X1   g0033(.A(G87), .B(G97), .Z(new_n234));
  XNOR2_X1  g0034(.A(G107), .B(G116), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n202), .A2(G68), .ZN(new_n237));
  INV_X1    g0037(.A(G68), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G50), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n236), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G1), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n244), .A2(G13), .A3(G20), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n210), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n244), .A2(G20), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n249), .A2(G50), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n211), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G150), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n252), .A2(new_n253), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n257), .B1(G20), .B2(new_n203), .ZN(new_n258));
  INV_X1    g0058(.A(new_n248), .ZN(new_n259));
  OAI221_X1 g0059(.A(new_n251), .B1(G50), .B2(new_n245), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT9), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT68), .ZN(new_n262));
  AND2_X1   g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n262), .B1(new_n263), .B2(new_n210), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n265), .A2(KEYINPUT68), .A3(G1), .A4(G13), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(G274), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT67), .B(G41), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n244), .B1(new_n268), .B2(G45), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G222), .A2(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(G223), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n271), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n263), .A2(new_n210), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n275), .B(new_n276), .C1(G77), .C2(new_n271), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n264), .A2(new_n266), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n244), .B1(G41), .B2(G45), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G226), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n270), .B(new_n277), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G200), .ZN(new_n284));
  INV_X1    g0084(.A(G190), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n261), .B(new_n284), .C1(new_n285), .C2(new_n283), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n286), .B(KEYINPUT10), .ZN(new_n287));
  OR2_X1    g0087(.A1(new_n283), .A2(G179), .ZN(new_n288));
  INV_X1    g0088(.A(G169), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n288), .A2(new_n260), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n246), .A2(new_n238), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT12), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n255), .A2(G50), .B1(G20), .B2(new_n238), .ZN(new_n295));
  INV_X1    g0095(.A(G77), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n295), .B1(new_n296), .B2(new_n253), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(KEYINPUT11), .A3(new_n248), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n249), .A2(G68), .A3(new_n250), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n294), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(KEYINPUT11), .B1(new_n297), .B2(new_n248), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n276), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n271), .A2(G232), .A3(G1698), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT70), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n304), .B(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n282), .A2(G1698), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n271), .A2(new_n307), .B1(G33), .B2(G97), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n303), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G238), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n270), .B1(new_n281), .B2(new_n310), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n309), .A2(KEYINPUT13), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT13), .B1(new_n309), .B2(new_n311), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n302), .B1(new_n315), .B2(new_n285), .ZN(new_n316));
  INV_X1    g0116(.A(G200), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n313), .B2(new_n314), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n302), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT14), .ZN(new_n321));
  INV_X1    g0121(.A(new_n314), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n321), .B(G169), .C1(new_n322), .C2(new_n312), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n313), .A2(G179), .A3(new_n314), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n321), .B1(new_n315), .B2(G169), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n320), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n319), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT16), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT7), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n271), .B2(G20), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT3), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G33), .ZN(new_n333));
  INV_X1    g0133(.A(G33), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT3), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n238), .B1(new_n331), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G58), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(new_n238), .ZN(new_n340));
  OAI21_X1  g0140(.A(G20), .B1(new_n340), .B2(new_n201), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n255), .A2(G159), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n329), .B1(new_n338), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT72), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT71), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n333), .A2(new_n335), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n332), .A2(KEYINPUT71), .A3(G33), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n211), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT7), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n348), .A2(new_n330), .A3(new_n211), .A4(new_n349), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(G68), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n343), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(KEYINPUT16), .A3(new_n354), .ZN(new_n355));
  OAI211_X1 g0155(.A(KEYINPUT72), .B(new_n329), .C1(new_n338), .C2(new_n343), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n346), .A2(new_n248), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n249), .ZN(new_n358));
  INV_X1    g0158(.A(new_n252), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n250), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n358), .A2(new_n360), .B1(new_n245), .B2(new_n359), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n348), .A2(new_n349), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n282), .A2(G1698), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(G223), .B2(G1698), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G87), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n303), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n264), .A2(G232), .A3(new_n266), .A4(new_n280), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n267), .B2(new_n269), .ZN(new_n372));
  OAI21_X1  g0172(.A(G169), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n372), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n366), .B1(new_n349), .B2(new_n348), .ZN(new_n375));
  INV_X1    g0175(.A(new_n369), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n276), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n374), .A2(G179), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n363), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT18), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n317), .B1(new_n370), .B2(new_n372), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n377), .A2(new_n270), .A3(new_n285), .A4(new_n371), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n382), .A2(KEYINPUT73), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT73), .B1(new_n382), .B2(new_n383), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n362), .B(new_n357), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT17), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT18), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n363), .A2(new_n389), .A3(new_n379), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n336), .B2(new_n211), .ZN(new_n391));
  AOI211_X1 g0191(.A(new_n330), .B(G20), .C1(new_n333), .C2(new_n335), .ZN(new_n392));
  OAI21_X1  g0192(.A(G68), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n354), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT72), .B1(new_n394), .B2(new_n329), .ZN(new_n395));
  INV_X1    g0195(.A(new_n356), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n355), .A2(new_n248), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n361), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT73), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n370), .A2(G190), .A3(new_n372), .ZN(new_n401));
  AOI21_X1  g0201(.A(G200), .B1(new_n374), .B2(new_n377), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n382), .A2(KEYINPUT73), .A3(new_n383), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n399), .A2(KEYINPUT17), .A3(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n381), .A2(new_n388), .A3(new_n390), .A4(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n249), .A2(G77), .A3(new_n250), .ZN(new_n408));
  XNOR2_X1  g0208(.A(KEYINPUT15), .B(G87), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n409), .A2(new_n253), .B1(new_n211), .B2(new_n296), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n252), .B1(KEYINPUT69), .B2(new_n256), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n256), .A2(KEYINPUT69), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI221_X1 g0213(.A(new_n408), .B1(G77), .B2(new_n245), .C1(new_n413), .C2(new_n259), .ZN(new_n414));
  NOR2_X1   g0214(.A1(G232), .A2(G1698), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n273), .A2(G238), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n271), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n417), .B(new_n276), .C1(G107), .C2(new_n271), .ZN(new_n418));
  INV_X1    g0218(.A(G244), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n270), .B(new_n418), .C1(new_n281), .C2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n414), .B1(G200), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n285), .B2(new_n420), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n289), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n423), .B(new_n414), .C1(G179), .C2(new_n420), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NOR4_X1   g0225(.A1(new_n292), .A2(new_n328), .A3(new_n407), .A4(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n273), .A2(KEYINPUT4), .A3(G244), .ZN(new_n427));
  INV_X1    g0227(.A(G250), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n427), .B1(new_n428), .B2(new_n273), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n429), .A2(new_n271), .B1(G33), .B2(G283), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  AOI211_X1 g0231(.A(new_n419), .B(G1698), .C1(new_n348), .C2(new_n349), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT4), .B1(new_n432), .B2(KEYINPUT74), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n364), .A2(G244), .A3(new_n273), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT74), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n431), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT75), .B1(new_n437), .B2(new_n303), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT4), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n434), .B2(new_n435), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n432), .A2(KEYINPUT74), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n430), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT75), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n443), .A3(new_n276), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT5), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n244), .B(G45), .C1(new_n445), .C2(G41), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n446), .B1(new_n268), .B2(new_n445), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(new_n278), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G257), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n279), .A2(G274), .A3(new_n447), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G179), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n438), .A2(new_n444), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n451), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n437), .B2(new_n303), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n289), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT6), .ZN(new_n457));
  INV_X1    g0257(.A(G97), .ZN(new_n458));
  INV_X1    g0258(.A(G107), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(G97), .A2(G107), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n457), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n459), .A2(KEYINPUT6), .A3(G97), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n464), .A2(G20), .B1(G77), .B2(new_n255), .ZN(new_n465));
  OAI21_X1  g0265(.A(G107), .B1(new_n391), .B2(new_n392), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n259), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n246), .A2(new_n458), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n334), .A2(G1), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n246), .A2(new_n248), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n468), .B1(new_n471), .B2(new_n458), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n453), .A2(new_n456), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT76), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n453), .A2(new_n456), .A3(new_n474), .A4(KEYINPUT76), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n438), .A2(new_n444), .A3(new_n454), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G200), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n451), .B1(new_n442), .B2(new_n276), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n474), .B1(new_n481), .B2(G190), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n477), .A2(new_n478), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n268), .A2(new_n445), .ZN(new_n484));
  INV_X1    g0284(.A(new_n446), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(new_n267), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n487), .B1(G270), .B2(new_n448), .ZN(new_n488));
  OR2_X1    g0288(.A1(KEYINPUT77), .A2(G116), .ZN(new_n489));
  NAND2_X1  g0289(.A1(KEYINPUT77), .A2(G116), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n470), .A2(G116), .B1(new_n246), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n489), .A2(G20), .A3(new_n490), .ZN(new_n494));
  AOI21_X1  g0294(.A(G20), .B1(G33), .B2(G283), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(G33), .B2(new_n458), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n496), .A3(new_n248), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT20), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n497), .A2(new_n498), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n493), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G257), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n273), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(G264), .B2(new_n273), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(new_n349), .B2(new_n348), .ZN(new_n505));
  INV_X1    g0305(.A(G303), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n271), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n276), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n488), .A2(new_n501), .A3(G179), .A4(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n279), .A2(new_n486), .A3(G270), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n450), .A3(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n511), .A2(new_n501), .A3(KEYINPUT21), .A4(G169), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n501), .A3(G169), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT21), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n501), .B1(new_n511), .B2(G200), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT79), .ZN(new_n520));
  INV_X1    g0320(.A(new_n511), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n519), .A2(new_n520), .B1(G190), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n317), .B1(new_n488), .B2(new_n508), .ZN(new_n523));
  OAI21_X1  g0323(.A(KEYINPUT79), .B1(new_n523), .B2(new_n501), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT80), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n525), .B1(new_n522), .B2(new_n524), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n518), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT81), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT25), .ZN(new_n530));
  AOI211_X1 g0330(.A(G107), .B(new_n245), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n529), .A2(new_n530), .ZN(new_n532));
  XNOR2_X1  g0332(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n470), .A2(G107), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n364), .A2(KEYINPUT22), .A3(new_n211), .A4(G87), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n211), .A2(G107), .ZN(new_n538));
  XNOR2_X1  g0338(.A(new_n538), .B(KEYINPUT23), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT22), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n211), .A2(G87), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n540), .B1(new_n336), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n491), .A2(new_n211), .A3(G33), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT24), .B1(new_n537), .B2(new_n544), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n539), .A2(new_n543), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT24), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n546), .A2(new_n536), .A3(new_n547), .A4(new_n542), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n535), .B1(new_n549), .B2(new_n248), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n448), .A2(G264), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n502), .A2(G1698), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(G250), .B2(G1698), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n349), .B2(new_n348), .ZN(new_n554));
  INV_X1    g0354(.A(G294), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n334), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n276), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n551), .A2(new_n557), .A3(new_n450), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n317), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT83), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n557), .A2(KEYINPUT82), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT82), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n562), .B(new_n276), .C1(new_n554), .C2(new_n556), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n561), .A2(new_n450), .A3(new_n563), .A4(new_n551), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n560), .B1(G190), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n559), .A2(KEYINPUT83), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n550), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n419), .A2(new_n273), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n364), .A2(new_n568), .B1(G33), .B2(new_n491), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n364), .A2(G238), .A3(new_n273), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n276), .ZN(new_n572));
  INV_X1    g0372(.A(G45), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n428), .B1(new_n573), .B2(G1), .ZN(new_n574));
  OR3_X1    g0374(.A1(new_n573), .A2(G1), .A3(G274), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n279), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n572), .A2(G190), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n303), .B1(new_n569), .B2(new_n570), .ZN(new_n578));
  INV_X1    g0378(.A(new_n576), .ZN(new_n579));
  OAI21_X1  g0379(.A(G200), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n364), .A2(new_n211), .A3(G68), .ZN(new_n582));
  AOI21_X1  g0382(.A(G20), .B1(G33), .B2(G97), .ZN(new_n583));
  INV_X1    g0383(.A(G87), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n583), .B1(new_n584), .B2(new_n461), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT19), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n253), .A2(KEYINPUT19), .A3(new_n458), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n582), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n589), .A2(new_n248), .B1(new_n246), .B2(new_n409), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n470), .A2(G87), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(G179), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n578), .A2(new_n579), .ZN(new_n594));
  INV_X1    g0394(.A(new_n409), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n470), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g0396(.A(new_n596), .B(KEYINPUT78), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n593), .A2(new_n594), .B1(new_n590), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n572), .A2(new_n576), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n289), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n581), .A2(new_n592), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n558), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n564), .A2(G169), .B1(new_n602), .B2(G179), .ZN(new_n603));
  OR2_X1    g0403(.A1(new_n603), .A2(new_n550), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n567), .A2(new_n601), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n528), .A2(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n426), .A2(new_n483), .A3(new_n606), .ZN(G372));
  INV_X1    g0407(.A(KEYINPUT84), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n599), .A2(new_n608), .A3(new_n289), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT84), .B1(new_n594), .B2(G169), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n611), .A2(new_n598), .B1(new_n581), .B2(new_n592), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n513), .B(new_n516), .C1(new_n603), .C2(new_n550), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n612), .A2(new_n567), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n477), .A2(new_n478), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n480), .A2(new_n482), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n477), .A2(new_n478), .A3(new_n601), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT26), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n611), .A2(new_n598), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n453), .A2(new_n456), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n473), .B1(new_n621), .B2(KEYINPUT85), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT85), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n453), .A2(new_n624), .A3(new_n456), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n622), .A2(new_n623), .A3(new_n612), .A4(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n617), .A2(new_n619), .A3(new_n620), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n426), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n291), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n381), .A2(new_n390), .ZN(new_n630));
  XOR2_X1   g0430(.A(new_n424), .B(KEYINPUT86), .Z(new_n631));
  NAND2_X1  g0431(.A1(new_n315), .A2(G169), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT14), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n633), .A2(new_n324), .A3(new_n323), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n631), .B1(new_n634), .B2(new_n320), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n319), .A2(new_n388), .A3(new_n406), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n630), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n629), .B1(new_n637), .B2(new_n287), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n628), .A2(new_n638), .ZN(G369));
  NAND3_X1  g0439(.A1(new_n244), .A2(new_n211), .A3(G13), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(G213), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(G343), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n501), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n517), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n528), .B2(new_n646), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G330), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n567), .A2(new_n604), .ZN(new_n651));
  INV_X1    g0451(.A(new_n645), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n550), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n604), .B2(new_n652), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n518), .A2(new_n645), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n604), .B2(new_n645), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n655), .A2(new_n659), .ZN(G399));
  INV_X1    g0460(.A(new_n207), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(new_n268), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G116), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n461), .A2(new_n584), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n663), .A2(G1), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n214), .B2(new_n663), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT28), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT90), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT31), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n599), .A2(KEYINPUT87), .A3(new_n593), .A4(new_n511), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT87), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n511), .A2(new_n593), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n673), .B1(new_n674), .B2(new_n594), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n672), .A2(new_n675), .A3(new_n558), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n551), .A2(new_n557), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n677), .A2(new_n578), .A3(new_n579), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n511), .A2(new_n593), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT30), .B1(new_n680), .B2(new_n455), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT30), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n481), .A2(new_n682), .A3(new_n679), .A4(new_n678), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n676), .A2(new_n479), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n645), .B1(new_n684), .B2(KEYINPUT88), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n676), .A2(new_n479), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n681), .A2(new_n683), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n686), .A2(KEYINPUT88), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n671), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n606), .A2(new_n483), .A3(new_n652), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n686), .A2(new_n687), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n645), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT89), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n618), .A2(new_n623), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n622), .A2(KEYINPUT26), .A3(new_n612), .A4(new_n625), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n620), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n483), .B2(new_n614), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n696), .B1(new_n702), .B2(new_n652), .ZN(new_n703));
  AOI211_X1 g0503(.A(KEYINPUT89), .B(new_n645), .C1(new_n699), .C2(new_n701), .ZN(new_n704));
  OAI21_X1  g0504(.A(KEYINPUT29), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n627), .A2(new_n652), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI211_X1 g0508(.A(new_n670), .B(new_n695), .C1(new_n705), .C2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n705), .A2(new_n708), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n670), .B1(new_n711), .B2(new_n695), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n669), .B1(new_n713), .B2(G1), .ZN(G364));
  AND2_X1   g0514(.A1(new_n211), .A2(G13), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n244), .B1(new_n715), .B2(G45), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n662), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n650), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n648), .A2(G330), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G13), .A2(G33), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G20), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n648), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n718), .B(KEYINPUT91), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n271), .A2(new_n207), .ZN(new_n728));
  INV_X1    g0528(.A(G355), .ZN(new_n729));
  OAI22_X1  g0529(.A1(new_n728), .A2(new_n729), .B1(G116), .B2(new_n207), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT92), .Z(new_n731));
  NOR2_X1   g0531(.A1(new_n242), .A2(new_n573), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n364), .A2(new_n661), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(new_n215), .B2(G45), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n731), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n210), .B1(G20), .B2(new_n289), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n724), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n727), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n211), .A2(new_n285), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n317), .A2(G179), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n336), .B1(new_n743), .B2(new_n506), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n593), .A2(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n211), .A2(G190), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G179), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(G311), .A2(new_n748), .B1(new_n751), .B2(G329), .ZN(new_n752));
  INV_X1    g0552(.A(G322), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n741), .A2(new_n745), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n211), .B1(new_n749), .B2(G190), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n744), .B(new_n755), .C1(G294), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n746), .A2(new_n742), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT95), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G283), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n211), .A2(new_n593), .A3(new_n317), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT93), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n285), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT96), .B(G326), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n763), .A2(G190), .ZN(new_n767));
  XNOR2_X1  g0567(.A(KEYINPUT33), .B(G317), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n758), .A2(new_n761), .A3(new_n766), .A4(new_n769), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT97), .Z(new_n771));
  OAI22_X1  g0571(.A1(new_n754), .A2(new_n339), .B1(new_n747), .B2(new_n296), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n764), .B2(G50), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT94), .ZN(new_n774));
  INV_X1    g0574(.A(new_n760), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n459), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G159), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n750), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT32), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n781), .B(new_n271), .C1(new_n584), .C2(new_n743), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n756), .A2(new_n458), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n779), .A2(new_n780), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n767), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n777), .B(new_n785), .C1(new_n238), .C2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n771), .B1(new_n774), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n740), .B1(new_n788), .B2(new_n737), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n719), .A2(new_n721), .B1(new_n726), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(G396));
  NAND2_X1  g0591(.A1(new_n414), .A2(new_n645), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n425), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(new_n631), .B2(new_n793), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n706), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n795), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n627), .A2(new_n652), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n718), .B1(new_n799), .B2(new_n694), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n695), .A2(new_n796), .A3(new_n798), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n737), .A2(new_n722), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n727), .B1(G77), .B2(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G283), .A2(new_n767), .B1(new_n764), .B2(G303), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n760), .A2(G87), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n754), .A2(new_n555), .B1(new_n750), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(new_n491), .B2(new_n748), .ZN(new_n810));
  INV_X1    g0610(.A(new_n743), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n271), .B(new_n783), .C1(G107), .C2(new_n811), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n806), .A2(new_n807), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n754), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G143), .A2(new_n814), .B1(new_n748), .B2(G159), .ZN(new_n815));
  INV_X1    g0615(.A(new_n764), .ZN(new_n816));
  INV_X1    g0616(.A(G137), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n815), .B1(new_n816), .B2(new_n817), .C1(new_n254), .C2(new_n786), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT34), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n364), .B1(new_n821), .B2(new_n750), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT98), .Z(new_n823));
  NAND2_X1  g0623(.A1(new_n760), .A2(G68), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n811), .A2(G50), .B1(new_n757), .B2(G58), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n820), .A2(new_n823), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n818), .A2(new_n819), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n813), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n805), .B1(new_n828), .B2(new_n737), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n797), .B2(new_n723), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT99), .Z(new_n831));
  NOR2_X1   g0631(.A1(new_n802), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G384));
  AOI211_X1 g0633(.A(new_n664), .B(new_n213), .C1(new_n464), .C2(KEYINPUT35), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(KEYINPUT35), .B2(new_n464), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT36), .Z(new_n836));
  OR3_X1    g0636(.A1(new_n340), .A2(new_n214), .A3(new_n296), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n244), .B(G13), .C1(new_n837), .C2(new_n237), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n711), .A2(new_n426), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n638), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n316), .A2(new_n318), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n320), .B(new_n645), .C1(new_n634), .C2(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n319), .B(new_n327), .C1(new_n302), .C2(new_n652), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n424), .A2(new_n645), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT100), .Z(new_n848));
  AOI21_X1  g0648(.A(new_n846), .B1(new_n798), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n355), .A2(new_n248), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT16), .B1(new_n353), .B2(new_n354), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n362), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n373), .A2(new_n378), .A3(new_n643), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n399), .A2(new_n405), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT101), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n852), .A2(new_n853), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n386), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT101), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(new_n859), .A3(KEYINPUT37), .ZN(new_n860));
  INV_X1    g0660(.A(new_n643), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n363), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n380), .A2(new_n862), .A3(new_n386), .A4(new_n855), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n856), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n852), .A2(new_n861), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n407), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT38), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n864), .A2(KEYINPUT38), .A3(new_n866), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n849), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n630), .A2(new_n861), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n862), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n407), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n380), .A2(new_n862), .A3(new_n386), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n863), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT38), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n869), .B(new_n870), .C1(KEYINPUT102), .C2(new_n880), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n864), .A2(KEYINPUT38), .A3(new_n866), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n882), .A2(new_n880), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT39), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n884), .A2(KEYINPUT102), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n881), .A2(KEYINPUT39), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n634), .A2(new_n320), .A3(new_n652), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n872), .B(new_n874), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n841), .B(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT88), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n691), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n684), .A2(KEYINPUT88), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n891), .A2(KEYINPUT31), .A3(new_n892), .A4(new_n645), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n689), .A2(new_n690), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n795), .B1(new_n843), .B2(new_n844), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT40), .B1(new_n896), .B2(new_n883), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT40), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n871), .A2(new_n898), .A3(new_n894), .A4(new_n895), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n426), .A2(new_n894), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n901), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(G330), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n889), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n244), .B2(new_n715), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n889), .A2(new_n904), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n839), .B1(new_n906), .B2(new_n907), .ZN(G367));
  INV_X1    g0708(.A(new_n733), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n228), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n738), .B1(new_n207), .B2(new_n409), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n727), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI221_X1 g0712(.A(new_n271), .B1(new_n756), .B2(new_n238), .C1(new_n817), .C2(new_n750), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n339), .A2(new_n743), .B1(new_n754), .B2(new_n254), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n202), .A2(new_n747), .B1(new_n759), .B2(new_n296), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(G143), .ZN(new_n917));
  OAI221_X1 g0717(.A(new_n916), .B1(new_n816), .B2(new_n917), .C1(new_n778), .C2(new_n786), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT46), .B1(new_n811), .B2(new_n491), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(G107), .B2(new_n757), .ZN(new_n920));
  INV_X1    g0720(.A(new_n364), .ZN(new_n921));
  INV_X1    g0721(.A(G283), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n458), .A2(new_n759), .B1(new_n747), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(G303), .B2(new_n814), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n811), .A2(KEYINPUT46), .A3(G116), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(G317), .B2(new_n751), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n920), .A2(new_n921), .A3(new_n924), .A4(new_n926), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n555), .A2(new_n786), .B1(new_n816), .B2(new_n808), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n918), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT47), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n912), .B1(new_n930), .B2(new_n737), .ZN(new_n931));
  OR3_X1    g0731(.A1(new_n620), .A2(new_n592), .A3(new_n652), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n612), .B1(new_n592), .B2(new_n652), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(new_n724), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n483), .B1(new_n473), .B2(new_n652), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n622), .A2(new_n625), .A3(new_n645), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(new_n657), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT42), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT103), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n940), .A2(new_n941), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n615), .B1(new_n939), .B2(new_n604), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n944), .B1(new_n652), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n932), .A2(new_n933), .ZN(new_n948));
  OR3_X1    g0748(.A1(new_n947), .A2(KEYINPUT43), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n655), .A2(new_n939), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n947), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  AND3_X1   g0754(.A1(new_n949), .A2(new_n950), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n950), .B1(new_n949), .B2(new_n954), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n662), .B(KEYINPUT41), .Z(new_n958));
  XNOR2_X1  g0758(.A(new_n649), .B(KEYINPUT104), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n657), .B1(new_n654), .B2(new_n656), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n960), .B1(KEYINPUT104), .B2(new_n649), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n713), .A2(KEYINPUT105), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n705), .A2(new_n708), .ZN(new_n965));
  AOI21_X1  g0765(.A(KEYINPUT90), .B1(new_n965), .B2(new_n694), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n963), .B1(new_n966), .B2(new_n709), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT105), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n939), .A2(new_n658), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT44), .Z(new_n971));
  NOR2_X1   g0771(.A1(new_n939), .A2(new_n658), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT45), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(new_n655), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n964), .A2(new_n969), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n958), .B1(new_n976), .B2(new_n713), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n957), .B1(new_n977), .B2(new_n717), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT106), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n957), .B(KEYINPUT106), .C1(new_n977), .C2(new_n717), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n936), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n982), .A2(KEYINPUT107), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n982), .A2(KEYINPUT107), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(G387));
  OAI211_X1 g0785(.A(new_n710), .B(new_n712), .C1(new_n961), .C2(new_n962), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n986), .A2(new_n662), .A3(new_n967), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n654), .A2(new_n725), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n728), .A2(new_n666), .B1(G107), .B2(new_n207), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n909), .B1(new_n232), .B2(G45), .ZN(new_n990));
  XOR2_X1   g0790(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n252), .B2(G50), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n573), .B1(new_n238), .B2(new_n296), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(new_n665), .B2(KEYINPUT108), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n359), .A2(new_n991), .A3(new_n202), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n665), .A2(KEYINPUT108), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n993), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n989), .B1(new_n990), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n727), .B1(new_n999), .B2(new_n739), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G159), .A2(new_n764), .B1(new_n767), .B2(new_n359), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n760), .A2(G97), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n202), .A2(new_n754), .B1(new_n743), .B2(new_n296), .ZN(new_n1003));
  XOR2_X1   g0803(.A(KEYINPUT110), .B(G150), .Z(new_n1004));
  OAI22_X1  g0804(.A1(new_n1004), .A2(new_n750), .B1(new_n747), .B2(new_n238), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n756), .A2(new_n409), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n921), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1001), .A2(new_n1002), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n759), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n491), .A2(new_n1010), .B1(new_n751), .B2(new_n765), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n743), .A2(new_n555), .B1(new_n756), .B2(new_n922), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G317), .A2(new_n814), .B1(new_n748), .B2(G303), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n816), .B2(new_n753), .C1(new_n808), .C2(new_n786), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT48), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n1015), .B2(new_n1014), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT49), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n921), .B(new_n1011), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1009), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1000), .B1(new_n1021), .B2(new_n737), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n963), .A2(new_n717), .B1(new_n988), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(KEYINPUT111), .B1(new_n987), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n987), .A2(KEYINPUT111), .A3(new_n1023), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(G393));
  NAND2_X1  g0827(.A1(new_n975), .A2(new_n717), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n939), .A2(new_n724), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n738), .B1(new_n458), .B2(new_n207), .C1(new_n909), .C2(new_n236), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n727), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT112), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n767), .A2(G303), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n757), .A2(new_n491), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n743), .A2(new_n922), .B1(new_n747), .B2(new_n555), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n271), .B(new_n1035), .C1(G322), .C2(new_n751), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n777), .A2(new_n1033), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n764), .A2(G317), .B1(G311), .B2(new_n814), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT52), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n764), .A2(G150), .B1(G159), .B2(new_n814), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT51), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n767), .A2(G50), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n743), .A2(new_n238), .B1(new_n750), .B2(new_n917), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n359), .B2(new_n748), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n756), .A2(new_n296), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n921), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1042), .A2(new_n807), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n1037), .A2(new_n1039), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1032), .B1(new_n1048), .B2(new_n737), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1029), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1028), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n975), .B1(new_n713), .B2(new_n963), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1052), .A2(new_n663), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1051), .B1(new_n1053), .B2(new_n976), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(G390));
  NAND2_X1  g0855(.A1(new_n901), .A2(G330), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT114), .ZN(new_n1057));
  AND3_X1   g0857(.A1(new_n1057), .A2(new_n840), .A3(new_n638), .ZN(new_n1058));
  INV_X1    g0858(.A(G330), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n795), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n894), .A2(new_n845), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT113), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n693), .A2(new_n1060), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n846), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n798), .A2(new_n848), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1065), .A2(new_n846), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n845), .B1(new_n894), .B2(new_n1060), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n847), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n797), .B1(new_n703), .B2(new_n704), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1069), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1058), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n887), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n886), .B1(new_n849), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1070), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n846), .B1(new_n1074), .B2(new_n1073), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n887), .B1(new_n882), .B2(new_n880), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1079), .B(new_n1080), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1078), .B1(new_n1068), .B2(new_n845), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n883), .A2(new_n885), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n876), .A2(new_n879), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT102), .B1(new_n1086), .B2(new_n868), .ZN(new_n1087));
  AOI21_X1  g0887(.A(KEYINPUT38), .B1(new_n864), .B2(new_n866), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1087), .A2(new_n882), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1085), .B1(new_n1089), .B2(new_n884), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1084), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n702), .A2(new_n652), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(KEYINPUT89), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n702), .A2(new_n696), .A3(new_n652), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n795), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n845), .B1(new_n1095), .B2(new_n847), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1082), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1091), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1083), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n663), .B1(new_n1077), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1057), .A2(new_n840), .A3(new_n638), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1069), .A2(new_n1075), .ZN(new_n1103));
  OR3_X1    g0903(.A1(new_n1100), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n727), .B1(new_n359), .B2(new_n804), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1004), .A2(new_n743), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT53), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT54), .B(G143), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n271), .B1(new_n747), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(G125), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n754), .A2(new_n821), .B1(new_n750), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G50), .B2(new_n1010), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1107), .A2(new_n1108), .B1(G159), .B2(new_n757), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1112), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(G128), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1118), .A2(new_n816), .B1(new_n786), .B2(new_n817), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n459), .A2(new_n786), .B1(new_n816), .B2(new_n922), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n271), .B(new_n1045), .C1(G87), .C2(new_n811), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n747), .A2(new_n458), .B1(new_n750), .B2(new_n555), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G116), .B2(new_n814), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n824), .A3(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1117), .A2(new_n1119), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1106), .B1(new_n1125), .B2(new_n737), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n1090), .B2(new_n723), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n1100), .B2(new_n716), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT115), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1105), .B1(new_n1130), .B2(new_n1131), .ZN(G378));
  OAI21_X1  g0932(.A(new_n718), .B1(G50), .B2(new_n804), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n292), .B(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n260), .A2(new_n861), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT118), .Z(new_n1137));
  XOR2_X1   g0937(.A(new_n1135), .B(new_n1137), .Z(new_n1138));
  NOR2_X1   g0938(.A1(new_n1138), .A2(new_n723), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n759), .A2(new_n339), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(G77), .B2(new_n811), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n238), .B2(new_n756), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n814), .A2(G107), .B1(new_n748), .B2(new_n595), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n922), .B2(new_n750), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n364), .A2(new_n268), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n1142), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n458), .B2(new_n786), .C1(new_n664), .C2(new_n816), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT116), .Z(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(KEYINPUT58), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1145), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n754), .A2(new_n1118), .B1(new_n747), .B2(new_n817), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n743), .A2(new_n1110), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT117), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1152), .B(new_n1154), .C1(G150), .C2(new_n757), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1155), .B1(new_n1113), .B2(new_n816), .C1(new_n821), .C2(new_n786), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1010), .A2(G159), .ZN(new_n1159));
  AOI211_X1 g0959(.A(G33), .B(G41), .C1(new_n751), .C2(G124), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1151), .B1(KEYINPUT58), .B2(new_n1148), .C1(new_n1157), .C2(new_n1161), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1133), .B(new_n1139), .C1(new_n737), .C2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n900), .A2(G330), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n873), .B1(new_n1090), .B2(new_n1078), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1164), .A2(new_n1165), .A3(new_n872), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1059), .B1(new_n897), .B2(new_n899), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n888), .A2(new_n1167), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1166), .A2(new_n1168), .A3(new_n1138), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1138), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1163), .B1(new_n1171), .B2(new_n717), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1058), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1173), .A2(new_n1171), .A3(KEYINPUT57), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT57), .B1(new_n1173), .B2(new_n1171), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n662), .B(new_n1174), .C1(new_n1175), .C2(KEYINPUT119), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT119), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1177), .B(KEYINPUT57), .C1(new_n1173), .C2(new_n1171), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1172), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT120), .ZN(G375));
  NAND2_X1  g0980(.A1(new_n846), .A2(new_n722), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT121), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n803), .A2(new_n238), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n727), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1140), .B1(G150), .B2(new_n748), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1185), .B(new_n364), .C1(new_n202), .C2(new_n756), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G159), .A2(new_n811), .B1(new_n751), .B2(G128), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n817), .B2(new_n754), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n821), .A2(new_n816), .B1(new_n786), .B2(new_n1110), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n555), .A2(new_n816), .B1(new_n786), .B2(new_n492), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n271), .B(new_n1007), .C1(G107), .C2(new_n748), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n458), .A2(new_n743), .B1(new_n754), .B2(new_n922), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G303), .B2(new_n751), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1192), .B(new_n1194), .C1(new_n296), .C2(new_n775), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n1189), .A2(new_n1190), .B1(new_n1191), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1184), .B1(new_n1196), .B2(new_n737), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1076), .A2(new_n717), .B1(new_n1182), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n958), .B1(new_n1058), .B2(new_n1076), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1103), .A2(new_n1102), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(G381));
  INV_X1    g1003(.A(KEYINPUT124), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT120), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1179), .B(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT123), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1179), .A2(new_n1205), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1179), .A2(new_n1205), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1209), .A2(KEYINPUT123), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1208), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1128), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1054), .A2(new_n1202), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT122), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1025), .A2(new_n790), .A3(new_n1026), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1215), .B1(new_n1216), .B2(G384), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1026), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(new_n1218), .A2(G396), .A3(new_n1024), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1219), .A2(KEYINPUT122), .A3(new_n832), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1214), .A2(new_n1217), .A3(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n983), .B2(new_n984), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1204), .B1(new_n1212), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n980), .A2(new_n981), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n935), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT107), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n982), .A2(KEYINPUT107), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1221), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1230), .A2(KEYINPUT124), .A3(new_n1208), .A4(new_n1211), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1224), .A2(new_n1231), .ZN(G407));
  INV_X1    g1032(.A(G213), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1212), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(G343), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1213), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1233), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(G407), .A2(new_n1237), .ZN(G409));
  AOI21_X1  g1038(.A(new_n790), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1239));
  OAI21_X1  g1039(.A(KEYINPUT107), .B1(new_n1239), .B2(new_n1219), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1054), .ZN(new_n1241));
  OAI21_X1  g1041(.A(G390), .B1(new_n1239), .B2(new_n1219), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1226), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(G396), .B1(new_n1218), .B2(new_n1024), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1227), .B1(new_n1244), .B2(new_n1216), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1242), .B1(new_n1245), .B2(G390), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n982), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1243), .A2(new_n1247), .ZN(new_n1248));
  XOR2_X1   g1048(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1249));
  OAI211_X1 g1049(.A(G378), .B(new_n1172), .C1(new_n1176), .C2(new_n1178), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1173), .A2(new_n1171), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1172), .B1(new_n1251), .B2(new_n958), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1213), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1235), .B1(new_n1250), .B2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1103), .A2(new_n1102), .A3(KEYINPUT60), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n662), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1077), .A2(KEYINPUT60), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1256), .B1(new_n1257), .B2(new_n1201), .ZN(new_n1258));
  OR3_X1    g1058(.A1(new_n1258), .A2(new_n832), .A3(new_n1199), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n832), .B1(new_n1258), .B2(new_n1199), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1249), .B1(new_n1254), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT126), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1250), .A2(new_n1253), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1235), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1264), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  AOI211_X1 g1067(.A(KEYINPUT126), .B(new_n1235), .C1(new_n1250), .C2(new_n1253), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1262), .A2(KEYINPUT62), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1263), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1235), .A2(G2897), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1261), .B(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT61), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1248), .B1(new_n1271), .B2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1243), .A2(new_n1247), .A3(new_n1275), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1261), .A2(new_n1272), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1261), .A2(new_n1272), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1254), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1278), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT63), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1261), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1269), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1254), .A2(new_n1262), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1283), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(KEYINPUT125), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT125), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1286), .A2(new_n1289), .A3(new_n1283), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1282), .A2(new_n1285), .A3(new_n1288), .A4(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1277), .A2(new_n1291), .ZN(G405));
  NAND2_X1  g1092(.A1(G375), .A2(new_n1213), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1293), .A2(new_n1250), .A3(new_n1261), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1261), .B1(new_n1293), .B2(new_n1250), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1248), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1293), .A2(new_n1250), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1262), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1248), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1293), .A2(new_n1250), .A3(new_n1261), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1296), .A2(new_n1301), .ZN(G402));
endmodule


