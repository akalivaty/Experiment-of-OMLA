//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n449, new_n450, new_n453, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n582, new_n583, new_n584, new_n585, new_n587, new_n588, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1209, new_n1210;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n449));
  AND2_X1   g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  NAND2_X1  g026(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI22_X1  g036(.A1(new_n456), .A2(new_n460), .B1(new_n461), .B2(new_n457), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT68), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n471), .B2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n475));
  AND4_X1   g050(.A1(new_n469), .A2(new_n472), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G137), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n469), .A2(G101), .A3(G2104), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT70), .Z(new_n479));
  NAND3_X1  g054(.A1(new_n468), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n476), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n469), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n472), .A2(new_n475), .A3(G2105), .A4(new_n473), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT71), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n485), .B1(new_n487), .B2(G124), .ZN(G162));
  AND2_X1   g063(.A1(KEYINPUT4), .A2(G138), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n472), .A2(new_n475), .A3(new_n473), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(G102), .A2(G2104), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(new_n469), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n472), .A2(new_n475), .A3(G126), .A4(new_n473), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n469), .A2(G138), .ZN(new_n498));
  AOI21_X1  g073(.A(KEYINPUT4), .B1(new_n464), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n493), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT72), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n499), .B1(new_n496), .B2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(new_n493), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(KEYINPUT74), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT73), .B1(new_n517), .B2(G651), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(new_n515), .A3(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n517), .A2(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(new_n513), .A3(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT75), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n521), .A2(new_n513), .A3(KEYINPUT75), .A4(new_n522), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(G88), .A3(new_n526), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n521), .A2(G543), .A3(new_n522), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G50), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT76), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n527), .A2(new_n532), .A3(new_n529), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n516), .B1(new_n531), .B2(new_n533), .ZN(G166));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XOR2_X1   g110(.A(new_n535), .B(KEYINPUT7), .Z(new_n536));
  NAND2_X1  g111(.A1(new_n528), .A2(G51), .ZN(new_n537));
  AND2_X1   g112(.A1(G63), .A2(G651), .ZN(new_n538));
  AOI21_X1  g113(.A(KEYINPUT77), .B1(new_n513), .B2(new_n538), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n513), .A2(KEYINPUT77), .A3(new_n538), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n536), .B1(new_n541), .B2(KEYINPUT78), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT78), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n537), .B(new_n543), .C1(new_n539), .C2(new_n540), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n525), .A2(new_n526), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G89), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n542), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(G168));
  NAND2_X1  g123(.A1(new_n545), .A2(G90), .ZN(new_n549));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(new_n513), .ZN(new_n551));
  INV_X1    g126(.A(G64), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n553), .A2(G651), .B1(new_n528), .B2(G52), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n549), .A2(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  NAND2_X1  g131(.A1(new_n545), .A2(G81), .ZN(new_n557));
  NAND2_X1  g132(.A1(G68), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G56), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n551), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n560), .A2(G651), .B1(new_n528), .B2(G43), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(new_n564));
  XOR2_X1   g139(.A(new_n564), .B(KEYINPUT79), .Z(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  NAND2_X1  g144(.A1(new_n545), .A2(G91), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n521), .A2(G53), .A3(G543), .A4(new_n522), .ZN(new_n571));
  AND2_X1   g146(.A1(KEYINPUT80), .A2(KEYINPUT9), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n513), .A2(G65), .ZN(new_n575));
  INV_X1    g150(.A(G78), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT81), .B1(new_n576), .B2(new_n509), .ZN(new_n577));
  OR3_X1    g152(.A1(new_n576), .A2(new_n509), .A3(KEYINPUT81), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n573), .A2(new_n574), .B1(G651), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n570), .A2(new_n580), .ZN(G299));
  NOR2_X1   g156(.A1(new_n547), .A2(KEYINPUT82), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT82), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n546), .A2(new_n544), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(new_n542), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(G286));
  INV_X1    g161(.A(new_n533), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n532), .B1(new_n527), .B2(new_n529), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n587), .A2(new_n588), .B1(new_n515), .B2(new_n514), .ZN(G303));
  INV_X1    g164(.A(G74), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n515), .B1(new_n551), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n528), .B2(G49), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n525), .A2(G87), .A3(new_n526), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G288));
  NAND3_X1  g170(.A1(new_n525), .A2(G86), .A3(new_n526), .ZN(new_n596));
  INV_X1    g171(.A(G61), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(new_n510), .B2(new_n512), .ZN(new_n598));
  AND2_X1   g173(.A1(G73), .A2(G543), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n521), .A2(G48), .A3(G543), .A4(new_n522), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT83), .ZN(G305));
  NAND2_X1  g179(.A1(new_n545), .A2(G85), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(KEYINPUT84), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(KEYINPUT84), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n607), .A2(G651), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT85), .B(G47), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n528), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n605), .A2(new_n609), .A3(new_n611), .ZN(G290));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NOR2_X1   g188(.A1(G301), .A2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n615), .A2(new_n515), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n528), .A2(G54), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n545), .A2(KEYINPUT10), .A3(G92), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT10), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n525), .A2(new_n526), .ZN(new_n621));
  INV_X1    g196(.A(G92), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n618), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT86), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n614), .B1(new_n625), .B2(new_n613), .ZN(G284));
  AOI21_X1  g201(.A(new_n614), .B1(new_n625), .B2(new_n613), .ZN(G321));
  NOR2_X1   g202(.A1(G299), .A2(G868), .ZN(new_n628));
  INV_X1    g203(.A(G286), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(G297));
  AOI21_X1  g205(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n625), .B1(new_n632), .B2(G860), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT87), .Z(G148));
  NAND2_X1  g209(.A1(new_n625), .A2(new_n632), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(KEYINPUT88), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n635), .A2(KEYINPUT88), .ZN(new_n638));
  OAI21_X1  g213(.A(G868), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(G868), .B2(new_n563), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT89), .ZN(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  INV_X1    g218(.A(G111), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n643), .B1(new_n644), .B2(G2105), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(new_n476), .B2(G135), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n487), .B2(G123), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT90), .B(G2096), .Z(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n469), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT12), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT13), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2100), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n651), .A2(new_n652), .A3(new_n656), .ZN(G156));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2427), .B(G2430), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(KEYINPUT14), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT91), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(new_n659), .B2(new_n660), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2451), .B(G2454), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT16), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G14), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(new_n670), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(G401));
  XOR2_X1   g249(.A(KEYINPUT93), .B(KEYINPUT18), .Z(new_n675));
  XNOR2_X1  g250(.A(G2084), .B(G2090), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT92), .ZN(new_n677));
  XOR2_X1   g252(.A(G2067), .B(G2678), .Z(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT94), .B(KEYINPUT17), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n677), .A2(new_n678), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n675), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2072), .B(G2078), .Z(new_n684));
  NOR2_X1   g259(.A1(new_n682), .A2(new_n675), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(new_n683), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2096), .B(G2100), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT95), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n687), .B(new_n689), .ZN(G227));
  XNOR2_X1  g265(.A(G1971), .B(G1976), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT19), .Z(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1956), .B(G2474), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1961), .B(G1966), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT20), .Z(new_n699));
  OR2_X1    g274(.A1(new_n695), .A2(new_n696), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n693), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT96), .Z(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n697), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT97), .Z(new_n704));
  OAI211_X1 g279(.A(new_n699), .B(new_n702), .C1(new_n692), .C2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1991), .B(G1996), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1981), .B(G1986), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n709), .B(new_n710), .Z(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(G229));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G22), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G166), .B2(new_n713), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT98), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(G1971), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(G23), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n594), .B2(new_n713), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT33), .Z(new_n720));
  INV_X1    g295(.A(G1976), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n716), .A2(G1971), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n713), .A2(G6), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT83), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n603), .B(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n724), .B1(new_n726), .B2(new_n713), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT32), .B(G1981), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n717), .A2(new_n722), .A3(new_n723), .A4(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT34), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(KEYINPUT34), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n713), .A2(G24), .ZN(new_n733));
  INV_X1    g308(.A(G290), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(new_n713), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n735), .A2(G1986), .ZN(new_n736));
  INV_X1    g311(.A(G29), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G25), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n476), .A2(G131), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n469), .A2(G107), .ZN(new_n740));
  OAI21_X1  g315(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n487), .B2(G119), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n738), .B1(new_n743), .B2(new_n737), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT35), .B(G1991), .Z(new_n745));
  XOR2_X1   g320(.A(new_n744), .B(new_n745), .Z(new_n746));
  NOR2_X1   g321(.A1(new_n735), .A2(G1986), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n736), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n731), .A2(new_n732), .A3(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT36), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n713), .A2(G21), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G168), .B2(new_n713), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT101), .B(G1966), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G2078), .ZN(new_n756));
  NOR2_X1   g331(.A1(G164), .A2(new_n737), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G27), .B2(new_n737), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n755), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n625), .A2(new_n713), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G4), .B2(new_n713), .ZN(new_n761));
  INV_X1    g336(.A(G1348), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n759), .B(new_n763), .C1(new_n756), .C2(new_n758), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n713), .A2(G19), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n563), .B2(new_n713), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(G1341), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n713), .A2(G5), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G171), .B2(new_n713), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n737), .A2(G32), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n487), .A2(G129), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n476), .A2(G141), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT26), .Z(new_n774));
  NAND3_X1  g349(.A1(new_n469), .A2(G105), .A3(G2104), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n771), .A2(new_n772), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n770), .B1(new_n776), .B2(G29), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT27), .B(G1996), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n769), .A2(G1961), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G29), .A2(G35), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G162), .B2(G29), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT29), .B(G2090), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT30), .B(G28), .ZN(new_n784));
  OR2_X1    g359(.A1(KEYINPUT31), .A2(G11), .ZN(new_n785));
  NAND2_X1  g360(.A1(KEYINPUT31), .A2(G11), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n784), .A2(new_n737), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(G34), .ZN(new_n788));
  AOI21_X1  g363(.A(G29), .B1(new_n788), .B2(KEYINPUT24), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(KEYINPUT24), .B2(new_n788), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n480), .B2(new_n737), .ZN(new_n791));
  INV_X1    g366(.A(G2084), .ZN(new_n792));
  OAI221_X1 g367(.A(new_n787), .B1(new_n791), .B2(new_n792), .C1(new_n649), .C2(new_n737), .ZN(new_n793));
  INV_X1    g368(.A(G2072), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n737), .A2(G33), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n796), .A2(new_n469), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT99), .Z(new_n798));
  NAND3_X1  g373(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT25), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n476), .B2(G139), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n795), .B1(new_n802), .B2(G29), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n793), .B1(new_n794), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n767), .A2(new_n779), .A3(new_n783), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n803), .A2(new_n794), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT100), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n713), .A2(G20), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT23), .Z(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G299), .B2(G16), .ZN(new_n810));
  INV_X1    g385(.A(G1956), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n737), .A2(G26), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT28), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n487), .A2(G128), .ZN(new_n815));
  OAI21_X1  g390(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n816));
  INV_X1    g391(.A(G116), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(G2105), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n476), .B2(G140), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n814), .B1(new_n820), .B2(G29), .ZN(new_n821));
  INV_X1    g396(.A(G2067), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NOR4_X1   g398(.A1(new_n805), .A2(new_n807), .A3(new_n812), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n791), .A2(new_n792), .ZN(new_n825));
  OAI221_X1 g400(.A(new_n825), .B1(new_n777), .B2(new_n778), .C1(new_n769), .C2(G1961), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT102), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n761), .A2(new_n762), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n764), .A2(new_n824), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n751), .A2(new_n829), .ZN(G311));
  INV_X1    g405(.A(G311), .ZN(G150));
  XOR2_X1   g406(.A(KEYINPUT104), .B(G860), .Z(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(G80), .A2(G543), .ZN(new_n834));
  INV_X1    g409(.A(G67), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n551), .B2(new_n835), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n836), .A2(G651), .B1(new_n528), .B2(G55), .ZN(new_n837));
  INV_X1    g412(.A(G93), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n838), .B2(new_n621), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n562), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT103), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n839), .B(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n841), .B1(new_n843), .B2(new_n563), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n625), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n833), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n848), .B2(new_n847), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n843), .A2(new_n832), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT37), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(G145));
  XNOR2_X1  g428(.A(G162), .B(new_n648), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n480), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n776), .B(new_n820), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n802), .ZN(new_n857));
  AOI21_X1  g432(.A(G2105), .B1(new_n490), .B2(new_n491), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n469), .B1(new_n494), .B2(new_n495), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n858), .A2(new_n859), .A3(new_n499), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT105), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n857), .B(new_n861), .Z(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n476), .A2(G142), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n469), .A2(G118), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(G130), .B2(new_n487), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(new_n654), .Z(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(new_n743), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT106), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n855), .B1(new_n863), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n862), .A2(KEYINPUT106), .A3(new_n870), .ZN(new_n873));
  AOI21_X1  g448(.A(G37), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n862), .A2(new_n870), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n862), .A2(new_n870), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n855), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(G395));
  NAND2_X1  g455(.A1(new_n726), .A2(KEYINPUT108), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT108), .ZN(new_n882));
  NAND2_X1  g457(.A1(G305), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(G290), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(G166), .B(new_n594), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n881), .A2(new_n883), .A3(G290), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n886), .ZN(new_n889));
  INV_X1    g464(.A(new_n887), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n889), .B1(new_n890), .B2(new_n884), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n893));
  OR2_X1    g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(KEYINPUT109), .B2(KEYINPUT42), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(KEYINPUT110), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n624), .A2(new_n570), .A3(new_n580), .ZN(new_n897));
  INV_X1    g472(.A(new_n618), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT10), .B1(new_n545), .B2(G92), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n621), .A2(new_n620), .A3(new_n622), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(G299), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n839), .B(KEYINPUT103), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n840), .B1(new_n904), .B2(new_n562), .ZN(new_n905));
  INV_X1    g480(.A(new_n638), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n905), .B1(new_n906), .B2(new_n636), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n637), .A2(new_n638), .A3(new_n844), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n903), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n844), .B1(new_n637), .B2(new_n638), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n636), .A3(new_n905), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n897), .A2(new_n902), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n913), .B1(new_n897), .B2(new_n902), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n912), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(KEYINPUT107), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n910), .A2(new_n911), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n909), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT110), .B1(new_n894), .B2(new_n895), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n896), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n894), .A2(new_n895), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n925), .A2(KEYINPUT110), .A3(new_n921), .A4(new_n909), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(G868), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n843), .A2(G868), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(G295));
  INV_X1    g506(.A(KEYINPUT111), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n928), .A2(new_n932), .A3(new_n930), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n613), .B1(new_n924), .B2(new_n926), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT111), .B1(new_n934), .B2(new_n929), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(G331));
  AND2_X1   g511(.A1(new_n888), .A2(new_n891), .ZN(new_n937));
  OAI21_X1  g512(.A(G171), .B1(new_n582), .B2(new_n585), .ZN(new_n938));
  NOR2_X1   g513(.A1(G168), .A2(G171), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n940), .A3(new_n844), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n547), .A2(KEYINPUT82), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n584), .A2(new_n583), .A3(new_n542), .ZN(new_n943));
  AOI21_X1  g518(.A(G301), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n905), .B1(new_n944), .B2(new_n939), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n918), .B2(new_n917), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n903), .B1(new_n941), .B2(new_n945), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n937), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n948), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n950), .B(new_n892), .C1(new_n920), .C2(new_n946), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n952));
  INV_X1    g527(.A(G37), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n949), .A2(new_n951), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT112), .ZN(new_n955));
  INV_X1    g530(.A(new_n946), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n948), .B1(new_n956), .B2(new_n919), .ZN(new_n957));
  AOI21_X1  g532(.A(G37), .B1(new_n957), .B2(new_n892), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n958), .A2(new_n959), .A3(new_n952), .A4(new_n949), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n955), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n915), .A2(new_n916), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n946), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n937), .B1(new_n964), .B2(new_n948), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n958), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n962), .B1(new_n966), .B2(KEYINPUT43), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n961), .A2(KEYINPUT113), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT113), .B1(new_n961), .B2(new_n967), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n952), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n958), .A2(KEYINPUT43), .A3(new_n949), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI22_X1  g547(.A1(new_n968), .A2(new_n969), .B1(KEYINPUT44), .B2(new_n972), .ZN(G397));
  INV_X1    g548(.A(KEYINPUT125), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n468), .A2(G40), .A3(new_n477), .A4(new_n479), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT114), .B1(new_n860), .B2(G1384), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n977));
  INV_X1    g552(.A(G1384), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n501), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n975), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(G2078), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT116), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n506), .A2(new_n985), .A3(KEYINPUT45), .A4(new_n978), .ZN(new_n986));
  NOR4_X1   g561(.A1(new_n858), .A2(new_n859), .A3(KEYINPUT72), .A4(new_n499), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n504), .B1(new_n503), .B2(new_n493), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT45), .B(new_n978), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT116), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n982), .A2(new_n984), .A3(new_n986), .A4(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1961), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n976), .A2(new_n993), .A3(new_n979), .ZN(new_n994));
  INV_X1    g569(.A(new_n975), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(G1384), .B1(new_n502), .B2(new_n505), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n997), .A2(new_n993), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n992), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(G1384), .B1(new_n503), .B2(new_n493), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n975), .B1(new_n1000), .B2(KEYINPUT45), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n756), .B(new_n1001), .C1(new_n997), .C2(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n983), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n991), .A2(new_n999), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(G171), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1000), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n981), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1007), .A2(new_n1001), .A3(new_n984), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n999), .A2(new_n1003), .A3(G301), .A4(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT54), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT49), .ZN(new_n1011));
  INV_X1    g586(.A(G1981), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n596), .A2(new_n602), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1012), .B1(new_n596), .B2(new_n602), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1011), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n603), .A2(G1981), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1017), .A2(KEYINPUT49), .A3(new_n1013), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n976), .A2(new_n995), .A3(new_n979), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1016), .A2(new_n1018), .A3(G8), .A4(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1021), .B(new_n1022), .C1(new_n594), .C2(G1976), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1976), .B1(new_n592), .B2(new_n593), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT115), .B1(new_n1024), .B2(KEYINPUT52), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n594), .A2(G1976), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1019), .A2(new_n1027), .A3(G8), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1020), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1028), .A2(KEYINPUT52), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1001), .B1(new_n997), .B2(KEYINPUT45), .ZN(new_n1032));
  INV_X1    g607(.A(G1971), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n978), .B1(new_n987), .B2(new_n988), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT50), .ZN(new_n1036));
  INV_X1    g611(.A(G2090), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1036), .A2(new_n1037), .A3(new_n995), .A4(new_n994), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n1040));
  INV_X1    g615(.A(G8), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(G166), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1039), .A2(new_n1044), .A3(G8), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n975), .B1(new_n997), .B2(new_n993), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n980), .A2(KEYINPUT50), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(new_n1037), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1041), .B1(new_n1048), .B2(new_n1034), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1031), .B(new_n1045), .C1(new_n1044), .C2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1010), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1000), .A2(new_n977), .ZN(new_n1053));
  AOI211_X1 g628(.A(KEYINPUT114), .B(G1384), .C1(new_n503), .C2(new_n493), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n981), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n990), .A2(new_n986), .A3(new_n995), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n754), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1036), .A2(new_n792), .A3(new_n995), .A4(new_n994), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1041), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n547), .A2(G8), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1060), .B(KEYINPUT122), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1052), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n996), .A2(new_n998), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n754), .A2(new_n1056), .B1(new_n1064), .B2(new_n792), .ZN(new_n1065));
  OAI211_X1 g640(.A(KEYINPUT51), .B(new_n1061), .C1(new_n1065), .C2(new_n1041), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1062), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1063), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n991), .A2(new_n999), .A3(G301), .A4(new_n1003), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(KEYINPUT123), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n999), .A2(new_n1003), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT123), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1073), .A2(new_n1074), .A3(G301), .A4(new_n991), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n999), .A2(new_n1003), .A3(new_n1008), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT124), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1076), .A2(new_n1077), .A3(G171), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1077), .B1(new_n1076), .B2(G171), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1072), .B(new_n1075), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1051), .A2(new_n1069), .A3(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n995), .B1(new_n1035), .B2(KEYINPUT50), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n993), .B1(new_n976), .B2(new_n979), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n811), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n570), .A2(new_n580), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT56), .B(G2072), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1001), .B(new_n1090), .C1(new_n997), .C2(KEYINPUT45), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1084), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(G1956), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1091), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1088), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n762), .B1(new_n996), .B2(new_n998), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1019), .A2(G2067), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n901), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1092), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1095), .A2(KEYINPUT61), .A3(new_n1092), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT119), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1095), .A2(new_n1103), .A3(new_n1092), .A4(KEYINPUT61), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1106), .B1(new_n624), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1097), .A2(new_n1098), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n624), .A2(new_n1107), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1110), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1097), .A2(new_n1098), .A3(new_n1108), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1106), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT121), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1095), .A2(new_n1092), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1001), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1120), .B1(new_n981), .B2(new_n1035), .ZN(new_n1121));
  XOR2_X1   g696(.A(KEYINPUT118), .B(G1996), .Z(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT58), .B(G1341), .Z(new_n1124));
  NAND2_X1  g699(.A1(new_n1019), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1126), .A2(new_n1127), .A3(new_n563), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1121), .A2(new_n1122), .B1(new_n1019), .B2(new_n1124), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT59), .B1(new_n1129), .B2(new_n562), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1118), .A2(new_n1119), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1111), .A2(new_n1115), .A3(new_n1132), .A4(new_n1113), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1105), .A2(new_n1117), .A3(new_n1131), .A4(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1081), .B1(new_n1100), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(G288), .A2(G1976), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1014), .B1(new_n1020), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1019), .A2(G8), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1045), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1139), .B1(new_n1140), .B2(new_n1031), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1067), .A2(G8), .A3(new_n629), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT117), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT117), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1059), .A2(new_n1144), .A3(new_n629), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1031), .A2(new_n1045), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1049), .A2(new_n1044), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT63), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1039), .A2(G8), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1151), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1152), .A2(KEYINPUT63), .A3(new_n1045), .A4(new_n1031), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1153), .B1(new_n1145), .B2(new_n1143), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1141), .B1(new_n1150), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n974), .B1(new_n1135), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1134), .A2(new_n1100), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1051), .A2(new_n1080), .A3(new_n1069), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1141), .ZN(new_n1160));
  NOR4_X1   g735(.A1(new_n1065), .A2(KEYINPUT117), .A3(new_n1041), .A4(G286), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1144), .B1(new_n1059), .B2(new_n629), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1149), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT63), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1153), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n1146), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1160), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1159), .A2(KEYINPUT125), .A3(new_n1168), .ZN(new_n1169));
  AOI211_X1 g744(.A(new_n1050), .B(new_n1005), .C1(new_n1069), .C2(KEYINPUT62), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1170), .B1(KEYINPUT62), .B2(new_n1069), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1156), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1007), .A2(new_n975), .ZN(new_n1173));
  INV_X1    g748(.A(G1996), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n776), .B(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n820), .A2(G2067), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n815), .A2(new_n822), .A3(new_n819), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n743), .B(new_n745), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(G290), .B(G1986), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1173), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1172), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n743), .A2(new_n745), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1177), .B1(new_n1179), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(new_n1173), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1173), .ZN(new_n1189));
  NOR3_X1   g764(.A1(new_n1189), .A2(G1986), .A3(G290), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT127), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(KEYINPUT48), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1192), .B1(new_n1189), .B2(new_n1181), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1191), .A2(KEYINPUT48), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1188), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1178), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1173), .B1(new_n1196), .B2(new_n776), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT46), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1198), .B1(new_n1189), .B2(G1996), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1173), .A2(KEYINPUT46), .A3(new_n1174), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1197), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  XOR2_X1   g776(.A(new_n1201), .B(KEYINPUT47), .Z(new_n1202));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n1203));
  AND2_X1   g778(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1205));
  NOR3_X1   g780(.A1(new_n1195), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1185), .A2(new_n1206), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g782(.A1(G227), .A2(new_n462), .ZN(new_n1209));
  OAI211_X1 g783(.A(new_n711), .B(new_n1209), .C1(new_n673), .C2(new_n672), .ZN(new_n1210));
  NOR3_X1   g784(.A1(new_n1210), .A2(new_n878), .A3(new_n972), .ZN(G308));
  INV_X1    g785(.A(G308), .ZN(G225));
endmodule


