//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n450, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT64), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g024(.A(G2106), .ZN(new_n450));
  NOR2_X1   g025(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G325));
  XNOR2_X1  g033(.A(new_n457), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI22_X1  g035(.A1(new_n454), .A2(new_n450), .B1(new_n460), .B2(new_n456), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT68), .Z(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n465), .B1(new_n470), .B2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n466), .A2(new_n467), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n463), .A2(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n476), .A2(KEYINPUT69), .A3(G137), .A4(new_n463), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n473), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n473), .A2(new_n463), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(new_n491), .A3(G2104), .ZN(new_n492));
  AND2_X1   g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n466), .B2(new_n467), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n466), .B2(new_n467), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n497), .B(new_n500), .C1(new_n467), .C2(new_n466), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n495), .B1(new_n499), .B2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  XOR2_X1   g079(.A(new_n504), .B(KEYINPUT71), .Z(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G62), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n503), .B1(new_n505), .B2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n507), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  INV_X1    g091(.A(new_n509), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  XOR2_X1   g096(.A(KEYINPUT70), .B(G88), .Z(new_n522));
  OAI21_X1  g097(.A(new_n516), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n512), .A2(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(new_n515), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n510), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n513), .A2(new_n514), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G89), .ZN(new_n532));
  NAND2_X1  g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n529), .A2(new_n534), .ZN(G168));
  NAND2_X1  g110(.A1(new_n515), .A2(G52), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n537), .B2(new_n521), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n503), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n538), .A2(new_n540), .ZN(G171));
  NAND2_X1  g116(.A1(new_n515), .A2(G43), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n543), .B2(new_n521), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n503), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  INV_X1    g127(.A(G65), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n508), .B2(new_n509), .ZN(new_n554));
  AND2_X1   g129(.A1(G78), .A2(G543), .ZN(new_n555));
  OAI21_X1  g130(.A(G651), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n513), .A2(new_n514), .B1(new_n508), .B2(new_n509), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G91), .ZN(new_n558));
  OAI211_X1 g133(.A(G53), .B(G543), .C1(new_n519), .C2(new_n520), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n556), .B(new_n558), .C1(new_n560), .C2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  INV_X1    g138(.A(G168), .ZN(G286));
  INV_X1    g139(.A(G166), .ZN(G303));
  NAND2_X1  g140(.A1(new_n515), .A2(G49), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n557), .A2(G87), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(G288));
  NAND2_X1  g145(.A1(G73), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT72), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n508), .B2(new_n509), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n557), .A2(G86), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n515), .A2(G48), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  XOR2_X1   g154(.A(new_n579), .B(KEYINPUT73), .Z(G305));
  AOI22_X1  g155(.A1(new_n557), .A2(G85), .B1(new_n515), .B2(G47), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n503), .B2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  INV_X1    g159(.A(G92), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n521), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT10), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n530), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G54), .B2(new_n515), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n584), .B1(new_n592), .B2(G868), .ZN(G321));
  XOR2_X1   g168(.A(G321), .B(KEYINPUT74), .Z(G284));
  NAND2_X1  g169(.A1(G286), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(G299), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(G868), .B2(new_n596), .ZN(G297));
  OAI21_X1  g172(.A(new_n595), .B1(G868), .B2(new_n596), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n592), .B1(new_n599), .B2(G860), .ZN(G148));
  OAI21_X1  g175(.A(KEYINPUT75), .B1(new_n547), .B2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n592), .A2(new_n599), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  MUX2_X1   g178(.A(KEYINPUT75), .B(new_n601), .S(new_n603), .Z(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n481), .A2(G135), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT77), .ZN(new_n607));
  OAI21_X1  g182(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n608));
  INV_X1    g183(.A(G111), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G2105), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(new_n483), .B2(G123), .ZN(new_n611));
  AND2_X1   g186(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(G2096), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n476), .A2(new_n464), .ZN(new_n615));
  XOR2_X1   g190(.A(KEYINPUT76), .B(KEYINPUT12), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(G2100), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(G2100), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n613), .A2(G2096), .ZN(new_n622));
  NAND4_X1  g197(.A1(new_n614), .A2(new_n620), .A3(new_n621), .A4(new_n622), .ZN(G156));
  XOR2_X1   g198(.A(KEYINPUT15), .B(G2435), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2438), .ZN(new_n625));
  XOR2_X1   g200(.A(G2427), .B(G2430), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT79), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n625), .A2(new_n627), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n628), .A2(KEYINPUT14), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G1341), .B(G1348), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2443), .B(G2446), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n631), .B(new_n632), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n630), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(G14), .B1(new_n634), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n639), .B1(new_n638), .B2(new_n634), .ZN(G401));
  XOR2_X1   g215(.A(G2072), .B(G2078), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  NAND3_X1  g219(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT18), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT80), .B(KEYINPUT17), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n641), .B(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n644), .ZN(new_n649));
  NOR3_X1   g224(.A1(new_n648), .A2(new_n643), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n649), .B1(new_n642), .B2(new_n643), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n648), .B2(new_n643), .ZN(new_n652));
  NOR3_X1   g227(.A1(new_n646), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2096), .B(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(G227));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT19), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  AND2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n659), .A2(new_n660), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  MUX2_X1   g241(.A(new_n666), .B(new_n665), .S(new_n658), .Z(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G1981), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  INV_X1    g249(.A(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G229));
  NOR2_X1   g253(.A1(G5), .A2(G16), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT93), .ZN(new_n680));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n680), .B1(G301), .B2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(G1961), .ZN(new_n684));
  INV_X1    g259(.A(G29), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G27), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT94), .ZN(new_n687));
  OAI21_X1  g262(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  AOI22_X1  g264(.A1(new_n476), .A2(new_n493), .B1(new_n689), .B2(new_n491), .ZN(new_n690));
  INV_X1    g265(.A(new_n501), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n500), .B1(new_n476), .B2(new_n497), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n687), .B1(new_n693), .B2(G29), .ZN(new_n694));
  INV_X1    g269(.A(G2078), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n483), .A2(G129), .ZN(new_n697));
  NAND3_X1  g272(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT26), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n481), .A2(G141), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n464), .A2(G105), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n704), .A2(new_n685), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n685), .B2(G32), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT27), .B(G1996), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n683), .A2(G1961), .ZN(new_n709));
  NAND4_X1  g284(.A1(new_n684), .A2(new_n696), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n694), .A2(new_n695), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT30), .ZN(new_n712));
  AND3_X1   g287(.A1(new_n712), .A2(KEYINPUT92), .A3(G28), .ZN(new_n713));
  AOI21_X1  g288(.A(KEYINPUT92), .B1(new_n712), .B2(G28), .ZN(new_n714));
  OAI221_X1 g289(.A(new_n685), .B1(new_n712), .B2(G28), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT31), .B(G11), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n715), .B(new_n716), .C1(new_n613), .C2(new_n685), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n681), .A2(G19), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n547), .B2(new_n681), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G1341), .ZN(new_n720));
  NOR4_X1   g295(.A1(new_n710), .A2(new_n711), .A3(new_n717), .A4(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT24), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n722), .A2(G34), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(G34), .ZN(new_n724));
  AOI21_X1  g299(.A(G29), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n479), .B2(G29), .ZN(new_n726));
  INV_X1    g301(.A(G2084), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G4), .A2(G16), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n592), .B2(G16), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n681), .A2(G20), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT23), .Z(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G299), .B2(G16), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT96), .B(G1956), .ZN(new_n734));
  OAI22_X1  g309(.A1(new_n730), .A2(G1348), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AOI211_X1 g310(.A(new_n728), .B(new_n735), .C1(G1348), .C2(new_n730), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n721), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n685), .A2(G35), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G162), .B2(new_n685), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT29), .Z(new_n740));
  INV_X1    g315(.A(G2090), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n740), .A2(KEYINPUT95), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n685), .A2(G26), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT28), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n481), .A2(G140), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n483), .A2(G128), .ZN(new_n746));
  OR2_X1    g321(.A1(G104), .A2(G2105), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n747), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n744), .B1(new_n750), .B2(new_n685), .ZN(new_n751));
  INV_X1    g326(.A(G2067), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n734), .A2(new_n733), .B1(new_n726), .B2(new_n727), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n742), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(KEYINPUT95), .B1(new_n740), .B2(new_n741), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(G115), .A2(G2104), .ZN(new_n758));
  INV_X1    g333(.A(G127), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n473), .B2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT90), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n463), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n761), .B2(new_n760), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT25), .ZN(new_n764));
  NAND2_X1  g339(.A1(G103), .A2(G2104), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(G2105), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n463), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n481), .A2(G139), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n770), .A2(new_n685), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n685), .B2(G33), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT91), .B(G2072), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n681), .A2(G21), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G168), .B2(new_n681), .ZN(new_n776));
  INV_X1    g351(.A(G1966), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n774), .B(new_n778), .C1(new_n706), .C2(new_n707), .ZN(new_n779));
  OAI22_X1  g354(.A1(new_n740), .A2(new_n741), .B1(new_n772), .B2(new_n773), .ZN(new_n780));
  NOR4_X1   g355(.A1(new_n737), .A2(new_n757), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G25), .A2(G29), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n481), .A2(G131), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT83), .ZN(new_n786));
  OAI21_X1  g361(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n787));
  INV_X1    g362(.A(G107), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(G2105), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n483), .B2(G119), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(KEYINPUT84), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT84), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n786), .A2(new_n793), .A3(new_n790), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n784), .B1(new_n795), .B2(new_n685), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT35), .B(G1991), .Z(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n681), .A2(G24), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT85), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G290), .B2(G16), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT86), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(new_n675), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n796), .A2(new_n797), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n798), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n579), .B(KEYINPUT73), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(G16), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G6), .B2(G16), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT32), .B(G1981), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n809), .A2(new_n810), .ZN(new_n813));
  OAI21_X1  g388(.A(KEYINPUT87), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n809), .A2(new_n810), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT87), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n815), .A2(new_n816), .A3(new_n811), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n681), .A2(G23), .ZN(new_n818));
  INV_X1    g393(.A(G288), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n681), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT33), .B(G1976), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n681), .A2(G22), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G166), .B2(new_n681), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G1971), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n814), .A2(new_n817), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n806), .B1(new_n827), .B2(KEYINPUT34), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n827), .A2(KEYINPUT88), .A3(KEYINPUT34), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(KEYINPUT88), .B1(new_n827), .B2(KEYINPUT34), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n829), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT89), .B(KEYINPUT36), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n832), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(new_n830), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n838), .A2(new_n829), .A3(new_n834), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n782), .B1(new_n836), .B2(new_n839), .ZN(G311));
  AOI21_X1  g415(.A(new_n834), .B1(new_n838), .B2(new_n829), .ZN(new_n841));
  AOI211_X1 g416(.A(new_n835), .B(new_n828), .C1(new_n837), .C2(new_n830), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n781), .B1(new_n841), .B2(new_n842), .ZN(G150));
  XOR2_X1   g418(.A(KEYINPUT98), .B(G55), .Z(new_n844));
  INV_X1    g419(.A(G93), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n527), .A2(new_n844), .B1(new_n521), .B2(new_n845), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n847), .A2(new_n503), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(G860), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT37), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n547), .ZN(new_n855));
  OAI21_X1  g430(.A(KEYINPUT99), .B1(new_n848), .B2(new_n846), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n547), .A2(new_n849), .A3(new_n853), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n592), .A2(G559), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n850), .B1(new_n863), .B2(KEYINPUT39), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n852), .B1(new_n864), .B2(new_n865), .ZN(G145));
  INV_X1    g441(.A(KEYINPUT105), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n499), .A2(new_n501), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n869));
  NAND2_X1  g444(.A1(G126), .A2(G2105), .ZN(new_n870));
  INV_X1    g445(.A(new_n467), .ZN(new_n871));
  NAND2_X1  g446(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n463), .A2(G114), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n874), .A2(new_n688), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n869), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n492), .A2(new_n494), .A3(KEYINPUT101), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n868), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n749), .ZN(new_n879));
  INV_X1    g454(.A(new_n704), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n770), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n879), .A2(new_n704), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n879), .A2(new_n704), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n769), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n617), .B(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n786), .A2(new_n793), .A3(new_n790), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n793), .B1(new_n786), .B2(new_n790), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n792), .A2(new_n794), .A3(new_n889), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n481), .A2(G142), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n483), .A2(G130), .ZN(new_n897));
  OR2_X1    g472(.A1(G106), .A2(G2105), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n898), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n900), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n893), .A2(new_n894), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(KEYINPUT104), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n887), .A2(new_n904), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n893), .A2(new_n894), .A3(new_n902), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n902), .B1(new_n893), .B2(new_n894), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(new_n886), .A3(KEYINPUT104), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(G160), .A2(G162), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n479), .A2(new_n487), .ZN(new_n912));
  OR3_X1    g487(.A1(new_n911), .A2(KEYINPUT100), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT100), .B1(new_n911), .B2(new_n912), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n913), .A2(new_n612), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n612), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n867), .B1(new_n910), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n917), .ZN(new_n919));
  AOI211_X1 g494(.A(KEYINPUT105), .B(new_n919), .C1(new_n905), .C2(new_n909), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G37), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n901), .A2(new_n903), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n917), .B1(new_n887), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n908), .A2(new_n886), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n882), .B(new_n885), .C1(new_n906), .C2(new_n907), .ZN(new_n928));
  AND4_X1   g503(.A1(new_n923), .A2(new_n926), .A3(new_n919), .A4(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n922), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT40), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n921), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n904), .B(new_n886), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT105), .B1(new_n933), .B2(new_n919), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n910), .A2(new_n867), .A3(new_n917), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n925), .A2(new_n923), .A3(new_n926), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n926), .A2(new_n919), .A3(new_n928), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT103), .ZN(new_n939));
  AOI21_X1  g514(.A(G37), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT40), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n932), .A2(new_n941), .ZN(G395));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n602), .B(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(new_n859), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n587), .A2(new_n591), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(G299), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n946), .B(new_n596), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT41), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n947), .A2(KEYINPUT41), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n945), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n948), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(G305), .A2(G166), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n807), .A2(G303), .ZN(new_n957));
  OR2_X1    g532(.A1(G288), .A2(G290), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n959));
  NAND2_X1  g534(.A1(G288), .A2(G290), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n956), .A2(new_n957), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n959), .B1(new_n958), .B2(new_n960), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n963), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n965), .A2(new_n957), .A3(new_n956), .A4(new_n961), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(KEYINPUT108), .B(KEYINPUT42), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n967), .B(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n955), .A2(new_n970), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n948), .A2(new_n969), .A3(new_n954), .ZN(new_n972));
  OAI21_X1  g547(.A(G868), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(G868), .B2(new_n849), .ZN(G295));
  OAI21_X1  g549(.A(new_n973), .B1(G868), .B2(new_n849), .ZN(G331));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n976));
  XNOR2_X1  g551(.A(G171), .B(G168), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n978), .A2(new_n857), .A3(new_n858), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n859), .A2(new_n977), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n953), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n979), .A2(new_n949), .A3(new_n980), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n967), .ZN(new_n986));
  AOI21_X1  g561(.A(G37), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n983), .A2(KEYINPUT110), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT109), .ZN(new_n990));
  OR3_X1    g565(.A1(new_n949), .A2(KEYINPUT109), .A3(new_n950), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(new_n991), .A3(new_n981), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n983), .A2(KEYINPUT110), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(new_n967), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n976), .B1(new_n987), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n967), .B1(new_n982), .B2(new_n984), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n953), .A2(new_n981), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n986), .A2(new_n998), .A3(new_n983), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n997), .A2(new_n999), .A3(new_n976), .A4(new_n922), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT44), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT111), .B1(new_n996), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n967), .B1(new_n983), .B2(KEYINPUT110), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(new_n992), .B2(new_n989), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n999), .A2(new_n922), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT43), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1006), .A2(new_n1007), .A3(KEYINPUT44), .A4(new_n1000), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n987), .A2(new_n995), .A3(new_n976), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n997), .A2(new_n999), .A3(new_n922), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT43), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1009), .A2(new_n1015), .ZN(G397));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n1017));
  INV_X1    g592(.A(G1384), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n877), .B1(new_n691), .B2(new_n692), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n690), .A2(KEYINPUT101), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT45), .B(new_n1018), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n471), .A2(G40), .A3(new_n478), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(G164), .B2(G1384), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1971), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n471), .A2(G40), .A3(new_n478), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1028), .A2(G2090), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT50), .B1(new_n878), .B2(new_n1018), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n1032));
  NOR3_X1   g607(.A1(G164), .A2(new_n1032), .A3(G1384), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1029), .B(new_n1030), .C1(new_n1031), .C2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1027), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1384), .B1(new_n868), .B2(new_n690), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT50), .ZN(new_n1037));
  AOI22_X1  g612(.A1(KEYINPUT101), .A2(new_n690), .B1(new_n499), .B2(new_n501), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1384), .B1(new_n1038), .B2(new_n876), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1037), .B1(new_n1039), .B2(KEYINPUT50), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1030), .B1(new_n1040), .B2(new_n1029), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1017), .B1(new_n1035), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G303), .A2(G8), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  NAND4_X1  g622(.A1(G303), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1029), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT113), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1051), .A2(KEYINPUT114), .A3(new_n1027), .A4(new_n1034), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1042), .A2(G8), .A3(new_n1049), .A4(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G86), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n578), .B1(new_n521), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n510), .A2(G61), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n571), .B(KEYINPUT72), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n503), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(G1981), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1981), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n576), .A2(new_n577), .A3(new_n1060), .A4(new_n578), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT49), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1039), .A2(new_n1022), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1059), .A2(KEYINPUT49), .A3(new_n1061), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1064), .A2(new_n1065), .A3(G8), .A4(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1068));
  OAI21_X1  g643(.A(G8), .B1(new_n1068), .B2(new_n1028), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n569), .A2(G1976), .A3(new_n567), .A4(new_n566), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1070), .B(KEYINPUT116), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT52), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1070), .B(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1976), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT52), .B1(G288), .B2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1074), .A2(new_n1065), .A3(G8), .A4(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1067), .A2(new_n1072), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1049), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1027), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n693), .A2(new_n1032), .A3(new_n1018), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1022), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1032), .B1(new_n878), .B2(new_n1018), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1082), .A2(new_n1083), .A3(G2090), .ZN(new_n1084));
  OAI21_X1  g659(.A(G8), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1078), .B1(new_n1079), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n693), .A2(new_n1018), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1028), .B1(new_n1087), .B2(new_n1023), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1088), .A2(new_n695), .A3(new_n1021), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1022), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT123), .B(G1961), .Z(new_n1092));
  AOI22_X1  g667(.A1(new_n1089), .A2(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1028), .B1(KEYINPUT45), .B2(new_n1036), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1068), .A2(new_n1023), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1094), .A2(new_n1095), .A3(KEYINPUT53), .A4(new_n695), .ZN(new_n1096));
  AOI21_X1  g671(.A(G301), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1053), .A2(new_n1086), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(G1966), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n471), .A2(new_n478), .A3(G40), .A4(new_n727), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1068), .A2(new_n1032), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1100), .B1(new_n1101), .B2(new_n1037), .ZN(new_n1102));
  OAI21_X1  g677(.A(G8), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G8), .ZN(new_n1104));
  NOR2_X1   g679(.A1(G168), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1105), .A2(KEYINPUT51), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1103), .A2(KEYINPUT122), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n693), .A2(KEYINPUT45), .A3(new_n1018), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1022), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT45), .B1(new_n878), .B2(new_n1018), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n777), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n727), .B(new_n1022), .C1(new_n1031), .C2(new_n1033), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1104), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1106), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1108), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT121), .B(KEYINPUT51), .Z(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n1114), .B2(new_n1105), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1107), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1105), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1098), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT62), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT127), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT127), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1124), .A2(new_n1127), .A3(KEYINPUT62), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1123), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1053), .A2(new_n1086), .ZN(new_n1130));
  OAI211_X1 g705(.A(KEYINPUT124), .B(new_n1022), .C1(new_n1039), .C2(KEYINPUT45), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1111), .B2(new_n1028), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n695), .A2(KEYINPUT53), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1134), .B1(new_n1039), .B2(KEYINPUT45), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1131), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1090), .B1(new_n1025), .B2(G2078), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(G171), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT126), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1139), .A2(new_n1142), .A3(G171), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1138), .A2(new_n1137), .A3(G301), .A4(new_n1096), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1144), .A2(KEYINPUT54), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1141), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1130), .A2(new_n1146), .A3(new_n1124), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1068), .A2(G2067), .A3(new_n1028), .ZN(new_n1148));
  INV_X1    g723(.A(G1348), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1148), .B1(new_n1091), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1150), .A2(new_n946), .ZN(new_n1151));
  INV_X1    g726(.A(G1956), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT56), .B(G2072), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1088), .A2(new_n1021), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT118), .ZN(new_n1156));
  AND3_X1   g731(.A1(G299), .A2(new_n1156), .A3(KEYINPUT57), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT57), .B1(G299), .B2(new_n1156), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1153), .A2(new_n1155), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1151), .A2(new_n1160), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1028), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1068), .A2(KEYINPUT50), .ZN(new_n1164));
  AOI21_X1  g739(.A(G1956), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AND4_X1   g740(.A1(new_n1022), .A2(new_n1021), .A3(new_n1024), .A4(new_n1154), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1162), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1161), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT59), .ZN(new_n1169));
  INV_X1    g744(.A(G1996), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1021), .A2(new_n1024), .A3(new_n1022), .A4(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT119), .ZN(new_n1172));
  XOR2_X1   g747(.A(KEYINPUT58), .B(G1341), .Z(new_n1173));
  AOI22_X1  g748(.A1(new_n1171), .A2(new_n1172), .B1(new_n1065), .B2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1088), .A2(KEYINPUT119), .A3(new_n1170), .A4(new_n1021), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n1169), .B(new_n855), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1065), .A2(new_n1173), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1177), .A2(new_n1175), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(KEYINPUT59), .B1(new_n1179), .B2(new_n547), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1176), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1167), .A2(new_n1160), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT60), .ZN(new_n1184));
  AOI211_X1 g759(.A(new_n946), .B(new_n1148), .C1(new_n1091), .C2(new_n1149), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1182), .A2(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  OR2_X1    g761(.A1(new_n1150), .A2(new_n592), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1150), .A2(new_n592), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1187), .A2(KEYINPUT60), .A3(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1181), .A2(new_n1186), .A3(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1167), .A2(KEYINPUT61), .A3(new_n1160), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT120), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1167), .A2(KEYINPUT120), .A3(KEYINPUT61), .A4(new_n1160), .ZN(new_n1194));
  AND2_X1   g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1168), .B1(new_n1190), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT54), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1139), .A2(G171), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1197), .B1(new_n1198), .B2(new_n1097), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(KEYINPUT125), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n1201));
  OAI211_X1 g776(.A(new_n1201), .B(new_n1197), .C1(new_n1198), .C2(new_n1097), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1147), .A2(new_n1196), .A3(new_n1203), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1042), .A2(G8), .A3(new_n1052), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1205), .A2(new_n1079), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1114), .A2(G168), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT63), .ZN(new_n1208));
  NOR3_X1   g783(.A1(new_n1207), .A2(new_n1078), .A3(new_n1208), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1206), .A2(new_n1053), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT117), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1206), .A2(KEYINPUT117), .A3(new_n1053), .A4(new_n1209), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1053), .A2(new_n1086), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1208), .B1(new_n1214), .B2(new_n1207), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1212), .A2(new_n1213), .A3(new_n1215), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1053), .A2(new_n1078), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1067), .A2(new_n1075), .A3(new_n819), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1069), .B1(new_n1218), .B2(new_n1061), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  NAND4_X1  g795(.A1(new_n1129), .A2(new_n1204), .A3(new_n1216), .A4(new_n1220), .ZN(new_n1221));
  NOR2_X1   g796(.A1(new_n1095), .A2(new_n1028), .ZN(new_n1222));
  XNOR2_X1  g797(.A(new_n704), .B(G1996), .ZN(new_n1223));
  XNOR2_X1  g798(.A(new_n749), .B(new_n752), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g800(.A(new_n795), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1225), .B1(new_n1226), .B2(new_n797), .ZN(new_n1227));
  OAI21_X1  g802(.A(new_n1227), .B1(new_n1226), .B2(new_n797), .ZN(new_n1228));
  NOR2_X1   g803(.A1(G290), .A2(G1986), .ZN(new_n1229));
  NOR2_X1   g804(.A1(new_n1229), .A2(KEYINPUT112), .ZN(new_n1230));
  NAND2_X1  g805(.A1(G290), .A2(G1986), .ZN(new_n1231));
  XOR2_X1   g806(.A(new_n1230), .B(new_n1231), .Z(new_n1232));
  OAI21_X1  g807(.A(new_n1222), .B1(new_n1228), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1221), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1222), .A2(new_n1229), .ZN(new_n1235));
  XOR2_X1   g810(.A(new_n1235), .B(KEYINPUT48), .Z(new_n1236));
  AOI21_X1  g811(.A(new_n1236), .B1(new_n1222), .B2(new_n1228), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1222), .A2(new_n1170), .ZN(new_n1238));
  XNOR2_X1  g813(.A(new_n1238), .B(KEYINPUT46), .ZN(new_n1239));
  INV_X1    g814(.A(new_n1224), .ZN(new_n1240));
  OAI21_X1  g815(.A(new_n1222), .B1(new_n1240), .B2(new_n880), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  XOR2_X1   g817(.A(new_n1242), .B(KEYINPUT47), .Z(new_n1243));
  NAND2_X1  g818(.A1(new_n1226), .A2(new_n797), .ZN(new_n1244));
  OAI22_X1  g819(.A1(new_n1244), .A2(new_n1225), .B1(G2067), .B2(new_n749), .ZN(new_n1245));
  AOI211_X1 g820(.A(new_n1237), .B(new_n1243), .C1(new_n1222), .C2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n1234), .A2(new_n1246), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g822(.A(G319), .ZN(new_n1249));
  NOR3_X1   g823(.A1(G401), .A2(new_n1249), .A3(G227), .ZN(new_n1250));
  NAND2_X1  g824(.A1(new_n677), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g825(.A(new_n1251), .B1(new_n1012), .B2(new_n1010), .ZN(new_n1252));
  NAND2_X1  g826(.A1(new_n936), .A2(new_n940), .ZN(new_n1253));
  AND2_X1   g827(.A1(new_n1252), .A2(new_n1253), .ZN(G308));
  NAND2_X1  g828(.A1(new_n1252), .A2(new_n1253), .ZN(G225));
endmodule


