//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008;
  INV_X1    g000(.A(KEYINPUT34), .ZN(new_n202));
  OAI22_X1  g001(.A1(KEYINPUT65), .A2(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT66), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n205));
  OAI221_X1 g004(.A(new_n205), .B1(KEYINPUT65), .B2(KEYINPUT24), .C1(G183gat), .C2(G190gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n209), .B(KEYINPUT64), .ZN(new_n210));
  NOR2_X1   g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n208), .A2(new_n210), .A3(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n207), .B1(new_n204), .B2(new_n206), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT25), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT68), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT26), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n211), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n220), .A3(new_n210), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT28), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT27), .B(G183gat), .ZN(new_n226));
  INV_X1    g025(.A(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n222), .A2(new_n223), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n226), .A2(new_n227), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n224), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n221), .A2(new_n229), .A3(new_n207), .A4(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT24), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n207), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n234), .B(new_n235), .C1(G183gat), .C2(G190gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n213), .A2(new_n236), .A3(new_n210), .A4(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n216), .A2(new_n232), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G127gat), .ZN(new_n240));
  INV_X1    g039(.A(G134gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G127gat), .A2(G134gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(KEYINPUT1), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n247));
  INV_X1    g046(.A(G120gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n247), .B1(new_n248), .B2(G113gat), .ZN(new_n249));
  INV_X1    g048(.A(G113gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n249), .B(new_n251), .C1(new_n250), .C2(G120gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT1), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n250), .A2(G120gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n248), .A2(G113gat), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n246), .A2(new_n252), .B1(new_n256), .B2(new_n245), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n252), .A2(new_n253), .A3(new_n244), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n245), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n216), .A2(new_n232), .A3(new_n261), .A4(new_n238), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G227gat), .A2(G233gat), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n202), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n264), .ZN(new_n266));
  AOI211_X1 g065(.A(KEYINPUT34), .B(new_n266), .C1(new_n258), .C2(new_n262), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT71), .B(G71gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(G99gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(G15gat), .B(G43gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n258), .A2(new_n266), .A3(new_n262), .ZN(new_n273));
  XOR2_X1   g072(.A(KEYINPUT70), .B(KEYINPUT33), .Z(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n272), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n273), .A2(KEYINPUT32), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n273), .B(KEYINPUT32), .C1(new_n275), .C2(new_n272), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n268), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n268), .B1(new_n278), .B2(new_n279), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(G78gat), .B(G106gat), .Z(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT31), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n284), .B(G50gat), .Z(new_n285));
  INV_X1    g084(.A(KEYINPUT81), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n287), .B(KEYINPUT82), .Z(new_n288));
  INV_X1    g087(.A(G228gat), .ZN(new_n289));
  INV_X1    g088(.A(G233gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293));
  INV_X1    g092(.A(G155gat), .ZN(new_n294));
  INV_X1    g093(.A(G162gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n293), .B1(new_n296), .B2(KEYINPUT2), .ZN(new_n297));
  INV_X1    g096(.A(G148gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n298), .A2(G141gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n297), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n298), .A2(G141gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(KEYINPUT2), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT2), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(KEYINPUT75), .ZN(new_n310));
  OAI22_X1  g109(.A1(new_n304), .A2(new_n306), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n296), .A2(new_n293), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n305), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n315));
  AND2_X1   g114(.A1(G197gat), .A2(G204gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(G197gat), .A2(G204gat), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT22), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g117(.A1(G211gat), .A2(G218gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(G211gat), .A2(G218gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT22), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n323), .A2(G211gat), .A3(G218gat), .ZN(new_n324));
  OAI22_X1  g123(.A1(new_n324), .A2(new_n319), .B1(new_n317), .B2(new_n316), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT29), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT79), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n315), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G211gat), .ZN(new_n329));
  INV_X1    g128(.A(G218gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT22), .ZN(new_n331));
  NAND2_X1  g130(.A1(G211gat), .A2(G218gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G197gat), .B(G204gat), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n318), .A2(new_n321), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NOR3_X1   g134(.A1(new_n335), .A2(KEYINPUT79), .A3(KEYINPUT29), .ZN(new_n336));
  OAI211_X1 g135(.A(KEYINPUT80), .B(new_n314), .C1(new_n328), .C2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT79), .B1(new_n335), .B2(KEYINPUT29), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n325), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n327), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(new_n315), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT80), .B1(new_n343), .B2(new_n314), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n301), .ZN(new_n346));
  OAI21_X1  g145(.A(G148gat), .B1(new_n346), .B2(new_n299), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n303), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n348), .A2(new_n297), .B1(new_n311), .B2(new_n312), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT29), .B1(new_n349), .B2(new_n315), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n350), .A2(new_n340), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n292), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n292), .B1(new_n350), .B2(new_n340), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n322), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n318), .A2(KEYINPUT78), .A3(new_n321), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n356), .A3(new_n325), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n341), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n349), .B1(new_n358), .B2(new_n315), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(G22gat), .B1(new_n352), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n314), .B1(new_n328), .B2(new_n336), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(new_n351), .A3(new_n337), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n291), .ZN(new_n366));
  INV_X1    g165(.A(G22gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n360), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n361), .A2(new_n369), .ZN(new_n370));
  OR2_X1    g169(.A1(new_n285), .A2(new_n286), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n288), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n367), .B1(new_n366), .B2(new_n368), .ZN(new_n373));
  AOI211_X1 g172(.A(G22gat), .B(new_n360), .C1(new_n365), .C2(new_n291), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n371), .B(new_n288), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n282), .B1(new_n372), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT85), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G226gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(new_n290), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(KEYINPUT29), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n239), .A2(KEYINPUT73), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT73), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n216), .A2(new_n232), .A3(new_n385), .A4(new_n238), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n383), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n239), .A2(new_n380), .A3(new_n290), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n335), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390));
  INV_X1    g189(.A(G64gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G92gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n384), .A2(new_n381), .A3(new_n386), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n239), .A2(new_n382), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(new_n340), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n389), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n398), .A2(KEYINPUT74), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(KEYINPUT74), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT30), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n389), .A2(new_n397), .ZN(new_n402));
  INV_X1    g201(.A(new_n394), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI211_X1 g203(.A(KEYINPUT30), .B(new_n394), .C1(new_n389), .C2(new_n397), .ZN(new_n405));
  OAI22_X1  g204(.A1(new_n399), .A2(new_n400), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n407));
  XNOR2_X1  g206(.A(G1gat), .B(G29gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G57gat), .B(G85gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n314), .A2(KEYINPUT3), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n349), .A2(new_n315), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n413), .A3(new_n261), .ZN(new_n414));
  NAND2_X1  g213(.A1(G225gat), .A2(G233gat), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n314), .A2(new_n261), .A3(KEYINPUT4), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n417), .B1(new_n257), .B2(new_n349), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n414), .B(new_n415), .C1(new_n416), .C2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT5), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n415), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n257), .A2(new_n349), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n314), .A2(new_n261), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n411), .B(new_n421), .C1(new_n426), .C2(new_n420), .ZN(new_n427));
  INV_X1    g226(.A(new_n411), .ZN(new_n428));
  INV_X1    g227(.A(new_n421), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n420), .B1(new_n419), .B2(new_n425), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n427), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n429), .A2(new_n430), .A3(new_n428), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT6), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n406), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n439));
  INV_X1    g238(.A(new_n288), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n375), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(KEYINPUT85), .A3(new_n282), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n379), .A2(new_n438), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT35), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT72), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n280), .A2(new_n281), .A3(new_n446), .ZN(new_n447));
  AND4_X1   g246(.A1(new_n446), .A2(new_n268), .A3(new_n278), .A4(new_n279), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n442), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT84), .B1(new_n434), .B2(KEYINPUT6), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n452), .B1(new_n436), .B2(KEYINPUT84), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n453), .A2(new_n406), .A3(KEYINPUT35), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n445), .A2(new_n455), .ZN(new_n456));
  OR3_X1    g255(.A1(new_n423), .A2(new_n424), .A3(new_n422), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n424), .A2(new_n417), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT4), .B1(new_n314), .B2(new_n261), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n257), .B1(new_n314), .B2(KEYINPUT3), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n458), .A2(new_n459), .B1(new_n460), .B2(new_n413), .ZN(new_n461));
  OAI211_X1 g260(.A(KEYINPUT39), .B(new_n457), .C1(new_n461), .C2(new_n415), .ZN(new_n462));
  OR2_X1    g261(.A1(new_n461), .A2(new_n415), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n428), .B(new_n462), .C1(new_n463), .C2(KEYINPUT39), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(KEYINPUT40), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n406), .A2(new_n427), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT83), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n402), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n394), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n402), .A2(new_n468), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT38), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n402), .A2(new_n403), .ZN(new_n473));
  OR3_X1    g272(.A1(new_n387), .A2(new_n335), .A3(new_n388), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n395), .A2(new_n396), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n474), .B(KEYINPUT37), .C1(new_n475), .C2(new_n340), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT38), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n476), .A2(new_n469), .A3(new_n477), .A4(new_n394), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n453), .A2(new_n472), .A3(new_n473), .A4(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT83), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n406), .A2(new_n480), .A3(new_n465), .A4(new_n427), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n467), .A2(new_n442), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n375), .B(new_n441), .C1(new_n406), .C2(new_n437), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n447), .B2(new_n448), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT36), .B1(new_n280), .B2(new_n281), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n456), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G15gat), .B(G22gat), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT16), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n491), .A2(G1gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(G1gat), .B2(new_n490), .ZN(new_n494));
  INV_X1    g293(.A(G8gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G43gat), .B(G50gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(G29gat), .A2(G36gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT14), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(G29gat), .B2(G36gat), .ZN(new_n500));
  INV_X1    g299(.A(G29gat), .ZN(new_n501));
  INV_X1    g300(.A(G36gat), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT14), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT15), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(G29gat), .A2(G36gat), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n506), .B1(KEYINPUT14), .B2(new_n498), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n507), .A2(new_n508), .A3(new_n503), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n497), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n500), .A2(new_n504), .A3(KEYINPUT15), .ZN(new_n511));
  INV_X1    g310(.A(new_n497), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n496), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT17), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n510), .A2(new_n516), .A3(new_n513), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n508), .B1(new_n507), .B2(new_n503), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n512), .B1(new_n511), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n509), .A2(new_n497), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT17), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n517), .A2(new_n521), .A3(new_n496), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n515), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G229gat), .A2(G233gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(KEYINPUT18), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n496), .B(new_n514), .ZN(new_n526));
  XOR2_X1   g325(.A(new_n524), .B(KEYINPUT13), .Z(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n515), .A2(new_n524), .A3(new_n522), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT18), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n525), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G113gat), .B(G141gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(G197gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT11), .ZN(new_n535));
  INV_X1    g334(.A(G169gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT12), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n535), .B(G169gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT12), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n532), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n542), .A2(new_n528), .A3(new_n525), .A4(new_n531), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n489), .A2(KEYINPUT86), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT86), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n445), .A2(new_n455), .B1(new_n482), .B2(new_n487), .ZN(new_n549));
  INV_X1    g348(.A(new_n546), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G57gat), .B(G64gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(G71gat), .A2(G78gat), .ZN(new_n554));
  INV_X1    g353(.A(G71gat), .ZN(new_n555));
  INV_X1    g354(.A(G78gat), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT9), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n553), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n391), .A2(G57gat), .ZN(new_n559));
  INV_X1    g358(.A(G57gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(G64gat), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT87), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n553), .A2(KEYINPUT87), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT9), .ZN(new_n565));
  XOR2_X1   g364(.A(G71gat), .B(G78gat), .Z(new_n566));
  AOI21_X1  g365(.A(new_n558), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568));
  INV_X1    g367(.A(G85gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(KEYINPUT8), .A2(new_n568), .B1(new_n569), .B2(new_n393), .ZN(new_n570));
  NAND2_X1  g369(.A1(G85gat), .A2(G92gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT90), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT89), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT7), .ZN(new_n575));
  NAND3_X1  g374(.A1(KEYINPUT90), .A2(G85gat), .A3(G92gat), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n575), .B1(new_n573), .B2(new_n576), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n570), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT91), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(new_n582), .A3(new_n568), .ZN(new_n583));
  INV_X1    g382(.A(new_n568), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT91), .B1(new_n584), .B2(new_n580), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n579), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n568), .A2(KEYINPUT8), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n588), .B1(G85gat), .B2(G92gat), .ZN(new_n589));
  AND3_X1   g388(.A1(KEYINPUT90), .A2(G85gat), .A3(G92gat), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT90), .B1(G85gat), .B2(G92gat), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n574), .B(KEYINPUT7), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n589), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n583), .A2(new_n585), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n567), .B1(new_n587), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n595), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n579), .A2(new_n586), .ZN(new_n599));
  INV_X1    g398(.A(new_n566), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n559), .A2(new_n561), .A3(KEYINPUT87), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n601), .A2(new_n562), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n600), .B1(new_n602), .B2(KEYINPUT9), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n598), .B(new_n599), .C1(new_n603), .C2(new_n558), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT10), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n597), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT93), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n599), .A2(new_n598), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(KEYINPUT10), .A3(new_n567), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n597), .A2(new_n604), .A3(KEYINPUT93), .A4(new_n605), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n608), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n604), .ZN(new_n615));
  INV_X1    g414(.A(new_n613), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G120gat), .B(G148gat), .ZN(new_n619));
  INV_X1    g418(.A(G176gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n621), .B(G204gat), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n614), .A2(new_n617), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT94), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n623), .A2(KEYINPUT94), .A3(new_n625), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n567), .A2(KEYINPUT21), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n496), .ZN(new_n632));
  XOR2_X1   g431(.A(G127gat), .B(G155gat), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(G231gat), .A2(G233gat), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n567), .A2(KEYINPUT21), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n638), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G183gat), .B(G211gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT20), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n641), .A2(new_n645), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G190gat), .B(G218gat), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n594), .B(new_n586), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n521), .A2(new_n517), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n519), .A2(new_n520), .ZN(new_n656));
  AOI211_X1 g455(.A(KEYINPUT92), .B(new_n655), .C1(new_n656), .C2(new_n609), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT92), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n510), .B(new_n513), .C1(new_n587), .C2(new_n596), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n658), .B1(new_n659), .B2(new_n654), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n653), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n654), .B1(new_n652), .B2(new_n514), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT92), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n659), .A2(new_n658), .A3(new_n654), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n662), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(new_n668), .A3(new_n653), .ZN(new_n669));
  XNOR2_X1  g468(.A(G134gat), .B(G162gat), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n663), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n671), .B1(new_n663), .B2(new_n669), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n651), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n668), .B1(new_n667), .B2(new_n653), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n521), .A2(new_n517), .A3(new_n652), .ZN(new_n676));
  AOI211_X1 g475(.A(new_n662), .B(new_n676), .C1(new_n665), .C2(new_n666), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n670), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n663), .A2(new_n669), .A3(new_n671), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(new_n650), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n649), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n552), .A2(new_n630), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n436), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT95), .B(G1gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1324gat));
  AND2_X1   g485(.A1(new_n552), .A2(new_n682), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n491), .B1(KEYINPUT96), .B2(KEYINPUT42), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n687), .A2(new_n630), .A3(new_n406), .A4(new_n688), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n491), .A2(KEYINPUT96), .A3(KEYINPUT42), .ZN(new_n690));
  OAI21_X1  g489(.A(G8gat), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n406), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n683), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n690), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n693), .A2(new_n495), .A3(new_n694), .A4(new_n688), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n691), .B(new_n695), .C1(KEYINPUT42), .C2(new_n693), .ZN(G1325gat));
  INV_X1    g495(.A(G15gat), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n485), .A2(new_n486), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n683), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n697), .B1(new_n683), .B2(new_n449), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT97), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n699), .B1(new_n702), .B2(new_n703), .ZN(G1326gat));
  NOR2_X1   g503(.A1(new_n683), .A2(new_n442), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT43), .B(G22gat), .Z(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1327gat));
  INV_X1    g506(.A(new_n630), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n648), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n681), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT98), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n552), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n713), .A2(new_n501), .A3(new_n437), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(KEYINPUT45), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n716));
  INV_X1    g515(.A(new_n681), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT44), .B1(new_n549), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n482), .A2(new_n487), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n444), .A2(KEYINPUT35), .B1(new_n451), .B2(new_n454), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n719), .B(new_n681), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n723), .A2(new_n546), .A3(new_n709), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n437), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n716), .B1(new_n725), .B2(G29gat), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n715), .B1(new_n726), .B2(new_n714), .ZN(G1328gat));
  NAND3_X1  g526(.A1(new_n713), .A2(new_n502), .A3(new_n406), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n728), .A2(KEYINPUT46), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n723), .A2(new_n546), .A3(new_n709), .ZN(new_n730));
  OR3_X1    g529(.A1(new_n730), .A2(KEYINPUT99), .A3(new_n692), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT99), .B1(new_n730), .B2(new_n692), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n731), .A2(G36gat), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n728), .A2(KEYINPUT46), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n729), .A2(new_n733), .A3(new_n734), .ZN(G1329gat));
  NOR3_X1   g534(.A1(new_n712), .A2(G43gat), .A3(new_n449), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(G43gat), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n730), .A2(new_n698), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n737), .B(KEYINPUT47), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n739), .A2(new_n738), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n742), .B2(new_n736), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(G1330gat));
  INV_X1    g543(.A(KEYINPUT48), .ZN(new_n745));
  OAI21_X1  g544(.A(G50gat), .B1(new_n730), .B2(new_n442), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT100), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n442), .A2(G50gat), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT101), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n552), .A2(new_n711), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT102), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n552), .A2(KEYINPUT102), .A3(new_n711), .A4(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n745), .B1(new_n748), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n751), .A2(KEYINPUT103), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT103), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n552), .A2(new_n758), .A3(new_n711), .A4(new_n750), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n759), .A3(KEYINPUT48), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n760), .B(new_n746), .C1(new_n747), .C2(KEYINPUT48), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n756), .A2(new_n761), .ZN(G1331gat));
  NAND3_X1  g561(.A1(new_n648), .A2(new_n550), .A3(new_n717), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n549), .A2(new_n630), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n437), .ZN(new_n765));
  XNOR2_X1  g564(.A(KEYINPUT104), .B(G57gat), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(G1332gat));
  INV_X1    g566(.A(new_n764), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT49), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n391), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n406), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT105), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT105), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n771), .A2(new_n774), .A3(new_n406), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n773), .A2(new_n775), .A3(new_n769), .A4(new_n391), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(G1333gat));
  OAI21_X1  g578(.A(new_n555), .B1(new_n768), .B2(new_n449), .ZN(new_n780));
  INV_X1    g579(.A(new_n698), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n764), .A2(G71gat), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g583(.A1(new_n764), .A2(new_n450), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g585(.A1(new_n648), .A2(new_n546), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n489), .A2(new_n681), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n790), .A2(KEYINPUT106), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n489), .A2(KEYINPUT51), .A3(new_n681), .A4(new_n787), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT106), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n630), .A2(new_n436), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n569), .ZN(new_n796));
  INV_X1    g595(.A(new_n787), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n797), .B1(new_n718), .B2(new_n722), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n798), .A2(new_n795), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n794), .A2(new_n796), .B1(new_n569), .B2(new_n799), .ZN(G1336gat));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n708), .A3(new_n406), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT107), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n798), .A2(KEYINPUT107), .A3(new_n708), .A4(new_n406), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(G92gat), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n630), .A2(new_n692), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n393), .B(new_n806), .C1(new_n791), .C2(new_n793), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n801), .A2(G92gat), .ZN(new_n810));
  INV_X1    g609(.A(new_n806), .ZN(new_n811));
  AOI211_X1 g610(.A(G92gat), .B(new_n811), .C1(new_n790), .C2(new_n792), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT52), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n809), .A2(new_n813), .ZN(G1337gat));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n708), .A3(new_n781), .ZN(new_n815));
  XOR2_X1   g614(.A(KEYINPUT108), .B(G99gat), .Z(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI221_X1 g616(.A(new_n708), .B1(new_n448), .B2(new_n447), .C1(new_n791), .C2(new_n793), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n818), .B2(new_n816), .ZN(G1338gat));
  NAND4_X1  g618(.A1(new_n723), .A2(new_n708), .A3(new_n450), .A4(new_n787), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT53), .B1(new_n820), .B2(G106gat), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n630), .A2(G106gat), .A3(new_n442), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n794), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n820), .A2(new_n825), .A3(G106gat), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n820), .B2(G106gat), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n823), .B1(new_n790), .B2(new_n792), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n824), .B1(new_n829), .B2(new_n830), .ZN(G1339gat));
  NAND4_X1  g630(.A1(new_n648), .A2(new_n630), .A3(new_n550), .A4(new_n717), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n523), .A2(new_n524), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n526), .A2(new_n527), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n537), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n545), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n612), .A2(new_n837), .A3(new_n613), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n612), .A2(new_n613), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n608), .A2(new_n610), .A3(new_n616), .A4(new_n611), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT54), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n622), .B(new_n838), .C1(new_n839), .C2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843));
  AOI221_X4 g642(.A(new_n836), .B1(new_n842), .B2(new_n843), .C1(new_n674), .C2(new_n680), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT110), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n845), .B1(new_n842), .B2(new_n843), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n838), .A2(new_n622), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n614), .A2(KEYINPUT54), .A3(new_n840), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n847), .A2(KEYINPUT110), .A3(KEYINPUT55), .A4(new_n848), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n846), .A2(new_n625), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n844), .A2(new_n850), .A3(KEYINPUT111), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT111), .ZN(new_n852));
  INV_X1    g651(.A(new_n836), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n842), .A2(new_n843), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n681), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n846), .A2(new_n625), .A3(new_n849), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n852), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI22_X1  g656(.A1(new_n842), .A2(new_n843), .B1(new_n544), .B2(new_n545), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n858), .A2(new_n846), .A3(new_n625), .A4(new_n849), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n628), .A2(new_n629), .A3(new_n853), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI22_X1  g660(.A1(new_n851), .A2(new_n857), .B1(new_n717), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n832), .B1(new_n862), .B2(new_n648), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n406), .A2(new_n436), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n451), .ZN(new_n866));
  OAI21_X1  g665(.A(G113gat), .B1(new_n866), .B2(new_n550), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n379), .A2(new_n443), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n546), .A2(new_n250), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n867), .B1(new_n869), .B2(new_n870), .ZN(G1340gat));
  OAI21_X1  g670(.A(G120gat), .B1(new_n866), .B2(new_n630), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT112), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n708), .A2(new_n248), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n869), .B2(new_n874), .ZN(G1341gat));
  NOR3_X1   g674(.A1(new_n866), .A2(new_n240), .A3(new_n649), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n869), .A2(new_n649), .ZN(new_n877));
  XOR2_X1   g676(.A(new_n877), .B(KEYINPUT113), .Z(new_n878));
  AOI21_X1  g677(.A(new_n876), .B1(new_n878), .B2(new_n240), .ZN(G1342gat));
  NAND3_X1  g678(.A1(new_n692), .A2(KEYINPUT114), .A3(new_n681), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT114), .B1(new_n692), .B2(new_n681), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n881), .A2(new_n436), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n241), .A3(new_n868), .ZN(new_n884));
  XOR2_X1   g683(.A(new_n884), .B(KEYINPUT56), .Z(new_n885));
  OAI21_X1  g684(.A(G134gat), .B1(new_n866), .B2(new_n717), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1343gat));
  NAND2_X1  g686(.A1(new_n861), .A2(new_n717), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT111), .B1(new_n844), .B2(new_n850), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n855), .A2(new_n856), .A3(new_n852), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n649), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n442), .B1(new_n892), .B2(new_n832), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n698), .A2(new_n864), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OR3_X1    g694(.A1(new_n895), .A2(G141gat), .A3(new_n550), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n894), .B(KEYINPUT115), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n863), .A2(new_n450), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT57), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n851), .A2(new_n857), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n854), .A2(KEYINPUT116), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n842), .A2(new_n903), .A3(new_n843), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(new_n546), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n860), .B1(new_n905), .B2(new_n856), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n717), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n648), .B1(new_n901), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n832), .ZN(new_n909));
  OAI211_X1 g708(.A(KEYINPUT57), .B(new_n450), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n897), .B1(new_n900), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(new_n546), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n300), .A2(new_n301), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n896), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT58), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n916), .B(new_n896), .C1(new_n912), .C2(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1344gat));
  NAND2_X1  g717(.A1(new_n900), .A2(new_n910), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n897), .A2(new_n630), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n855), .A2(new_n856), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n923), .B1(new_n906), .B2(new_n717), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n832), .B1(new_n924), .B2(new_n648), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n925), .A2(new_n899), .A3(new_n450), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n899), .B1(new_n863), .B2(new_n450), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n921), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n930));
  INV_X1    g729(.A(new_n895), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n920), .B1(new_n931), .B2(new_n708), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n922), .B(new_n930), .C1(G148gat), .C2(new_n932), .ZN(G1345gat));
  NAND3_X1  g732(.A1(new_n911), .A2(G155gat), .A3(new_n648), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n294), .B1(new_n895), .B2(new_n649), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT117), .ZN(G1346gat));
  NAND4_X1  g736(.A1(new_n883), .A2(new_n295), .A3(new_n450), .A4(new_n698), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n911), .A2(new_n681), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(new_n295), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT118), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT118), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n942), .B(new_n938), .C1(new_n939), .C2(new_n295), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1347gat));
  AOI21_X1  g743(.A(new_n437), .B1(new_n892), .B2(new_n832), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n868), .A2(new_n406), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n946), .A2(KEYINPUT119), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(KEYINPUT119), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n536), .A3(new_n546), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n945), .A2(new_n406), .A3(new_n451), .ZN(new_n952));
  OAI21_X1  g751(.A(G169gat), .B1(new_n952), .B2(new_n550), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1348gat));
  AND4_X1   g753(.A1(G176gat), .A2(new_n945), .A3(new_n451), .A4(new_n806), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n950), .A2(new_n708), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n955), .B1(new_n956), .B2(new_n620), .ZN(G1349gat));
  NAND4_X1  g756(.A1(new_n948), .A2(new_n226), .A3(new_n648), .A4(new_n949), .ZN(new_n958));
  NAND2_X1  g757(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n959));
  OAI21_X1  g758(.A(G183gat), .B1(new_n952), .B2(new_n649), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g760(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT121), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n961), .B(new_n963), .Z(G1350gat));
  NAND3_X1  g763(.A1(new_n950), .A2(new_n227), .A3(new_n681), .ZN(new_n965));
  OAI21_X1  g764(.A(G190gat), .B1(new_n952), .B2(new_n717), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n966), .A2(KEYINPUT61), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n966), .A2(KEYINPUT61), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n965), .B1(new_n968), .B2(new_n969), .ZN(G1351gat));
  INV_X1    g769(.A(KEYINPUT122), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n971), .B1(new_n926), .B2(new_n927), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n781), .A2(new_n437), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(new_n406), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT123), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n925), .A2(new_n899), .A3(new_n450), .ZN(new_n976));
  OAI211_X1 g775(.A(KEYINPUT122), .B(new_n976), .C1(new_n893), .C2(new_n899), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n972), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g777(.A(G197gat), .B1(new_n978), .B2(new_n550), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n898), .A2(new_n974), .ZN(new_n980));
  INV_X1    g779(.A(G197gat), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n980), .A2(new_n981), .A3(new_n546), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n979), .A2(new_n982), .ZN(G1352gat));
  NAND4_X1  g782(.A1(new_n972), .A2(new_n708), .A3(new_n975), .A4(new_n977), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(G204gat), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n811), .A2(G204gat), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n893), .A2(new_n973), .A3(new_n986), .ZN(new_n987));
  XOR2_X1   g786(.A(new_n987), .B(KEYINPUT62), .Z(new_n988));
  NAND2_X1  g787(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(KEYINPUT124), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT124), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n985), .A2(new_n988), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n992), .ZN(G1353gat));
  NAND3_X1  g792(.A1(new_n928), .A2(new_n648), .A3(new_n975), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(KEYINPUT126), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT126), .ZN(new_n996));
  NAND4_X1  g795(.A1(new_n928), .A2(new_n996), .A3(new_n975), .A4(new_n648), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n995), .A2(G211gat), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(KEYINPUT63), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT63), .ZN(new_n1000));
  NAND4_X1  g799(.A1(new_n995), .A2(new_n997), .A3(new_n1000), .A4(G211gat), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n980), .A2(new_n329), .A3(new_n648), .ZN(new_n1002));
  XNOR2_X1  g801(.A(new_n1002), .B(KEYINPUT125), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .ZN(G1354gat));
  NAND2_X1  g803(.A1(new_n681), .A2(G218gat), .ZN(new_n1005));
  XNOR2_X1  g804(.A(new_n1005), .B(KEYINPUT127), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n978), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g806(.A(G218gat), .B1(new_n980), .B2(new_n681), .ZN(new_n1008));
  NOR2_X1   g807(.A1(new_n1007), .A2(new_n1008), .ZN(G1355gat));
endmodule


