//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n203), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n209), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n202), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n211), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT64), .Z(new_n234));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n217), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G50), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n255), .B1(new_n208), .B2(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n252), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n254), .A2(new_n256), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n259), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT66), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(new_n209), .A3(new_n260), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT66), .B1(G20), .B2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n264), .B1(G150), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n258), .B1(new_n269), .B2(new_n251), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT9), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n260), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(G222), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G77), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(G223), .ZN(new_n280));
  OAI221_X1 g0080(.A(new_n277), .B1(new_n278), .B2(new_n275), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G1), .A3(G13), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  INV_X1    g0086(.A(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n283), .A2(new_n208), .A3(G274), .A4(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n283), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n290), .B1(G226), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n285), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G190), .ZN(new_n297));
  XNOR2_X1  g0097(.A(KEYINPUT67), .B(G200), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n271), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT10), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT15), .B(G87), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n303), .A2(new_n262), .B1(new_n209), .B2(new_n278), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n263), .B1(new_n266), .B2(new_n267), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n250), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n208), .A2(G20), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G77), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n306), .B1(G77), .B2(new_n252), .C1(new_n253), .C2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n275), .A2(G232), .A3(new_n276), .ZN(new_n310));
  INV_X1    g0110(.A(G107), .ZN(new_n311));
  OAI221_X1 g0111(.A(new_n310), .B1(new_n311), .B2(new_n275), .C1(new_n279), .C2(new_n221), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n284), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n290), .B1(G244), .B2(new_n293), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n309), .B1(new_n315), .B2(G169), .ZN(new_n316));
  INV_X1    g0116(.A(G179), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(KEYINPUT68), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT68), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n313), .A2(new_n314), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(G179), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n316), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n315), .A2(G190), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n309), .B1(new_n320), .B2(new_n299), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n295), .A2(G179), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n327), .B(new_n270), .C1(G169), .C2(new_n296), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n302), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(KEYINPUT3), .A2(G33), .ZN(new_n330));
  NOR2_X1   g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  OAI211_X1 g0131(.A(G226), .B(new_n276), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT69), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n275), .A2(KEYINPUT69), .A3(G226), .A4(new_n276), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g0136(.A(G232), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n283), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n289), .B1(new_n221), .B2(new_n292), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT13), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n342), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT13), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n339), .B1(new_n334), .B2(new_n335), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n344), .B(new_n345), .C1(new_n346), .C2(new_n283), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n343), .A2(new_n347), .A3(KEYINPUT70), .ZN(new_n348));
  INV_X1    g0148(.A(new_n341), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT70), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n349), .A2(new_n350), .A3(new_n345), .A4(new_n344), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n348), .A2(new_n351), .A3(G169), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT14), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n348), .A2(new_n351), .A3(KEYINPUT14), .A4(G169), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n343), .A2(G179), .A3(new_n347), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT11), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n262), .A2(new_n278), .B1(new_n209), .B2(G68), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT71), .B1(new_n268), .B2(G50), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n268), .A2(KEYINPUT71), .A3(G50), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n359), .B1(new_n364), .B2(new_n251), .ZN(new_n365));
  INV_X1    g0165(.A(new_n363), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(new_n361), .ZN(new_n367));
  OAI211_X1 g0167(.A(KEYINPUT11), .B(new_n250), .C1(new_n367), .C2(new_n360), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n202), .B1(new_n208), .B2(G20), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT12), .B1(new_n252), .B2(G68), .ZN(new_n370));
  OR3_X1    g0170(.A1(new_n252), .A2(KEYINPUT12), .A3(G68), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n254), .A2(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n365), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n358), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT72), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n348), .A2(new_n351), .A3(G200), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n373), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n343), .A2(new_n347), .A3(G190), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n375), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n376), .A2(KEYINPUT72), .A3(new_n378), .A4(new_n379), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT74), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n330), .A2(new_n331), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT7), .B1(new_n385), .B2(new_n209), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT7), .ZN(new_n387));
  NOR4_X1   g0187(.A1(new_n330), .A2(new_n331), .A3(new_n387), .A4(G20), .ZN(new_n388));
  OAI21_X1  g0188(.A(G68), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT16), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G58), .A2(G68), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n203), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G20), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT73), .B1(new_n268), .B2(G159), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT73), .ZN(new_n395));
  INV_X1    g0195(.A(G159), .ZN(new_n396));
  AOI211_X1 g0196(.A(new_n395), .B(new_n396), .C1(new_n266), .C2(new_n267), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n393), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n250), .B1(new_n390), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n267), .ZN(new_n400));
  NOR3_X1   g0200(.A1(KEYINPUT66), .A2(G20), .A3(G33), .ZN(new_n401));
  OAI21_X1  g0201(.A(G159), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n395), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n268), .A2(KEYINPUT73), .A3(G159), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n403), .A2(new_n404), .B1(G20), .B2(new_n392), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT16), .B1(new_n405), .B2(new_n389), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n384), .B1(new_n399), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G200), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n280), .A2(new_n276), .ZN(new_n409));
  INV_X1    g0209(.A(G226), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G1698), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n409), .B(new_n411), .C1(new_n330), .C2(new_n331), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n284), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n283), .A2(G232), .A3(new_n291), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n289), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT76), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n283), .B1(new_n412), .B2(new_n413), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n289), .A2(new_n416), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT76), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n408), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n419), .A2(new_n420), .ZN(new_n424));
  INV_X1    g0224(.A(G190), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n405), .A2(KEYINPUT16), .A3(new_n389), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT16), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n387), .B1(new_n275), .B2(G20), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n385), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n202), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n429), .B1(new_n398), .B2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n428), .A2(new_n433), .A3(KEYINPUT74), .A4(new_n250), .ZN(new_n434));
  INV_X1    g0234(.A(new_n263), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n307), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n436), .A2(new_n253), .B1(new_n252), .B2(new_n435), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT75), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n407), .A2(new_n427), .A3(new_n434), .A4(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT17), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n428), .A2(new_n433), .A3(new_n250), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n438), .B1(new_n443), .B2(new_n384), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n444), .A2(KEYINPUT17), .A3(new_n427), .A4(new_n434), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n407), .A2(new_n434), .A3(new_n439), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n418), .A2(new_n422), .ZN(new_n448));
  INV_X1    g0248(.A(G169), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n448), .A2(new_n449), .B1(new_n317), .B2(new_n424), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT18), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n447), .A2(KEYINPUT18), .A3(new_n450), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n446), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n329), .A2(new_n374), .A3(new_n383), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n275), .A2(new_n209), .A3(G68), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT19), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n209), .B1(new_n338), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(G87), .B2(new_n206), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT79), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n261), .A2(G97), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(new_n459), .ZN(new_n464));
  AOI211_X1 g0264(.A(KEYINPUT79), .B(KEYINPUT19), .C1(new_n261), .C2(G97), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n458), .B(new_n461), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n250), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n208), .A2(G33), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n252), .A2(new_n468), .A3(new_n217), .A4(new_n249), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(new_n222), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT81), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n470), .B(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n303), .A2(new_n257), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n467), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(G244), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n475));
  OAI211_X1 g0275(.A(G238), .B(new_n276), .C1(new_n330), .C2(new_n331), .ZN(new_n476));
  INV_X1    g0276(.A(G116), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n475), .B(new_n476), .C1(new_n260), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n284), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT78), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n208), .A2(G45), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(new_n223), .ZN(new_n483));
  INV_X1    g0283(.A(G274), .ZN(new_n484));
  INV_X1    g0284(.A(new_n217), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n485), .B2(new_n282), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n483), .A2(new_n283), .B1(new_n486), .B2(new_n482), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n479), .A2(new_n480), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n480), .B1(new_n479), .B2(new_n487), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n488), .A2(new_n489), .A3(new_n425), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n474), .B1(new_n490), .B2(KEYINPUT82), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n479), .A2(new_n487), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT78), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n479), .A2(new_n480), .A3(new_n487), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(G190), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n298), .B1(new_n493), .B2(new_n494), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT82), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n488), .A2(new_n489), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n467), .A2(new_n473), .ZN(new_n500));
  XOR2_X1   g0300(.A(new_n303), .B(KEYINPUT80), .Z(new_n501));
  INV_X1    g0301(.A(new_n469), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n499), .A2(new_n317), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n493), .A2(new_n494), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n449), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n491), .A2(new_n498), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(G257), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n508));
  OAI211_X1 g0308(.A(G250), .B(new_n276), .C1(new_n330), .C2(new_n331), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G294), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n284), .ZN(new_n512));
  OR2_X1    g0312(.A1(KEYINPUT5), .A2(G41), .ZN(new_n513));
  NAND2_X1  g0313(.A1(KEYINPUT5), .A2(G41), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n481), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n486), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n513), .A2(new_n514), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n517), .A2(new_n482), .B1(new_n485), .B2(new_n282), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G264), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n512), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n449), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(G179), .B2(new_n520), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n275), .A2(new_n209), .A3(G87), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT85), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n524), .A2(KEYINPUT22), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n275), .A2(new_n209), .A3(G87), .A4(new_n525), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n524), .A2(KEYINPUT22), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT24), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT23), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n209), .B2(G107), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n311), .A2(KEYINPUT23), .A3(G20), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n533), .A2(new_n534), .B1(new_n261), .B2(G116), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n530), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n531), .B1(new_n530), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n250), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n257), .A2(KEYINPUT25), .A3(new_n311), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT86), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT25), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n252), .B2(G107), .ZN(new_n542));
  OR2_X1    g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n540), .A2(new_n542), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n543), .A2(new_n544), .B1(G107), .B2(new_n502), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n522), .B1(new_n538), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n530), .A2(new_n535), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT24), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n530), .A2(new_n531), .A3(new_n535), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n251), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n545), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n520), .A2(new_n408), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(G190), .B2(new_n520), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n546), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n518), .A2(G270), .B1(new_n486), .B2(new_n515), .ZN(new_n556));
  OAI211_X1 g0356(.A(G264), .B(G1698), .C1(new_n330), .C2(new_n331), .ZN(new_n557));
  OAI211_X1 g0357(.A(G257), .B(new_n276), .C1(new_n330), .C2(new_n331), .ZN(new_n558));
  XNOR2_X1  g0358(.A(KEYINPUT83), .B(G303), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n557), .B(new_n558), .C1(new_n275), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n284), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n502), .A2(G116), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n257), .A2(new_n477), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n249), .A2(new_n217), .B1(G20), .B2(new_n477), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G283), .ZN(new_n566));
  INV_X1    g0366(.A(G97), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n566), .B(new_n209), .C1(G33), .C2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(KEYINPUT20), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT20), .B1(new_n565), .B2(new_n568), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n563), .B(new_n564), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n562), .A2(new_n572), .A3(G169), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT21), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n556), .A2(new_n561), .A3(G179), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n572), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n562), .A2(new_n572), .A3(KEYINPUT21), .A4(G169), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT84), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n556), .A2(new_n561), .A3(G190), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n564), .B1(new_n469), .B2(new_n477), .ZN(new_n582));
  INV_X1    g0382(.A(new_n571), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n582), .B1(new_n583), .B2(new_n569), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n408), .B1(new_n556), .B2(new_n561), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n580), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n586), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n588), .A2(KEYINPUT84), .A3(new_n584), .A4(new_n581), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n311), .A2(KEYINPUT6), .A3(G97), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n567), .A2(new_n311), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n592), .A2(new_n205), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n591), .B1(new_n593), .B2(KEYINPUT6), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n594), .A2(G20), .B1(G77), .B2(new_n268), .ZN(new_n595));
  OAI21_X1  g0395(.A(G107), .B1(new_n386), .B2(new_n388), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n250), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n252), .A2(G97), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n502), .B2(G97), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n276), .B1(new_n273), .B2(new_n274), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n602), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n603));
  OAI211_X1 g0403(.A(G244), .B(new_n276), .C1(new_n330), .C2(new_n331), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT4), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(G1698), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n607), .B(G244), .C1(new_n331), .C2(new_n330), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(KEYINPUT77), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT77), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n275), .A2(new_n610), .A3(G244), .A4(new_n607), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n603), .A2(new_n606), .A3(new_n609), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n284), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n517), .A2(new_n482), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n614), .A2(G257), .A3(new_n283), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n516), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n449), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n616), .B1(new_n612), .B2(new_n284), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n317), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n601), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n618), .A2(G200), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n620), .A2(G190), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n623), .A2(new_n598), .A3(new_n600), .A4(new_n624), .ZN(new_n625));
  AND4_X1   g0425(.A1(new_n579), .A2(new_n590), .A3(new_n622), .A4(new_n625), .ZN(new_n626));
  AND4_X1   g0426(.A1(new_n457), .A2(new_n507), .A3(new_n555), .A4(new_n626), .ZN(G372));
  INV_X1    g0427(.A(new_n622), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n507), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT26), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n474), .B1(new_n299), .B2(new_n492), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n495), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n499), .A2(new_n317), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n500), .A2(new_n503), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n492), .A2(new_n449), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n538), .A2(new_n545), .A3(new_n554), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n625), .A2(new_n622), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n512), .A2(new_n516), .A3(new_n519), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n317), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n641), .B(new_n521), .C1(new_n550), .C2(new_n551), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n579), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n637), .A2(new_n638), .A3(new_n639), .A4(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n637), .A2(new_n645), .A3(new_n628), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n630), .A2(new_n644), .A3(new_n636), .A4(new_n646), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n457), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT87), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n447), .A2(new_n649), .A3(new_n450), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n649), .B1(new_n447), .B2(new_n450), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n452), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n451), .A2(KEYINPUT87), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n447), .A2(new_n649), .A3(new_n450), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(KEYINPUT18), .A3(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n442), .A2(new_n445), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n322), .B1(new_n377), .B2(new_n380), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n374), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n656), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n302), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n328), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n648), .A2(new_n662), .ZN(G369));
  NAND3_X1  g0463(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G213), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n579), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n555), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n669), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n546), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n642), .B(new_n638), .C1(new_n552), .C2(new_n672), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n642), .B2(new_n672), .ZN(new_n677));
  INV_X1    g0477(.A(G330), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n579), .B(new_n590), .C1(new_n584), .C2(new_n672), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(new_n572), .A3(new_n669), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n678), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n675), .A2(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n212), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G1), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n215), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT88), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n618), .A2(new_n692), .A3(new_n520), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT88), .B1(new_n620), .B2(new_n640), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n562), .A2(new_n492), .A3(new_n317), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n695), .A2(KEYINPUT90), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n512), .A2(new_n519), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n576), .A2(new_n620), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n699), .B1(new_n702), .B2(new_n505), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n562), .A2(new_n700), .A3(new_n317), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n499), .A2(new_n704), .A3(KEYINPUT30), .A4(new_n620), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n698), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n696), .B1(new_n693), .B2(new_n694), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(KEYINPUT90), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n669), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT31), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n626), .A2(new_n507), .A3(new_n555), .A4(new_n672), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n672), .A2(new_n710), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n499), .A2(new_n620), .A3(new_n704), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n707), .B1(new_n699), .B2(new_n716), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n717), .A2(KEYINPUT89), .ZN(new_n718));
  INV_X1    g0518(.A(new_n705), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n717), .B2(KEYINPUT89), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n715), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(G330), .B1(new_n713), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n507), .A2(new_n645), .A3(new_n628), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n632), .A2(new_n636), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT26), .B1(new_n724), .B2(new_n622), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n636), .B(KEYINPUT91), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n644), .A2(new_n723), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n672), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT29), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n647), .A2(new_n730), .A3(new_n672), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n722), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n691), .B1(new_n732), .B2(G1), .ZN(G364));
  INV_X1    g0533(.A(G13), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n208), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n686), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n682), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n679), .A2(new_n681), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n739), .B1(G330), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT92), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n685), .A2(new_n385), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G355), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(G116), .B2(new_n212), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n685), .A2(new_n275), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n287), .B2(new_n216), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n247), .A2(G45), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n745), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(G20), .B1(KEYINPUT93), .B2(G169), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(KEYINPUT93), .A2(G169), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n217), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G13), .A2(G33), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n738), .B1(new_n750), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n757), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n740), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n209), .A2(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n764), .A2(new_n317), .A3(G200), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT94), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT94), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n298), .A2(new_n764), .A3(G179), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n768), .A2(G311), .B1(G283), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G190), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  XOR2_X1   g0573(.A(KEYINPUT33), .B(G317), .Z(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G179), .A2(G200), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n209), .B1(new_n776), .B2(G190), .ZN(new_n777));
  INV_X1    g0577(.A(G294), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n209), .A2(new_n425), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(G179), .A3(new_n408), .ZN(new_n780));
  INV_X1    g0580(.A(G322), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n385), .B1(new_n777), .B2(new_n778), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n771), .A2(new_n425), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n775), .B(new_n782), .C1(G326), .C2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n299), .A2(new_n317), .A3(new_n779), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n763), .A2(new_n776), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT97), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G303), .A2(new_n786), .B1(new_n788), .B2(G329), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n770), .A2(new_n784), .A3(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n768), .A2(KEYINPUT95), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n768), .A2(KEYINPUT95), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n278), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n773), .A2(new_n202), .ZN(new_n795));
  INV_X1    g0595(.A(new_n787), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G159), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT96), .B(KEYINPUT32), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n797), .A2(new_n798), .B1(new_n567), .B2(new_n777), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n795), .B(new_n799), .C1(new_n797), .C2(new_n798), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n785), .A2(new_n222), .ZN(new_n801));
  INV_X1    g0601(.A(new_n783), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n275), .B1(new_n780), .B2(new_n201), .C1(new_n255), .C2(new_n802), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n801), .B(new_n803), .C1(G107), .C2(new_n769), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n790), .B1(new_n794), .B2(new_n805), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n760), .B(new_n762), .C1(new_n754), .C2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n742), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G396));
  NAND2_X1  g0609(.A1(new_n647), .A2(new_n672), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n309), .A2(new_n669), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n325), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n322), .A2(new_n309), .A3(new_n669), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n647), .A2(new_n672), .A3(new_n814), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n738), .B1(new_n818), .B2(new_n722), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n722), .B2(new_n818), .ZN(new_n820));
  INV_X1    g0620(.A(new_n738), .ZN(new_n821));
  INV_X1    g0621(.A(new_n754), .ZN(new_n822));
  INV_X1    g0622(.A(G150), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n773), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(G137), .ZN(new_n825));
  INV_X1    g0625(.A(G143), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n825), .A2(new_n802), .B1(new_n780), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n793), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n824), .B(new_n827), .C1(new_n828), .C2(G159), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n829), .A2(KEYINPUT34), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(KEYINPUT34), .ZN(new_n831));
  INV_X1    g0631(.A(new_n788), .ZN(new_n832));
  INV_X1    g0632(.A(G132), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n769), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n202), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n275), .B1(new_n777), .B2(new_n201), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n785), .A2(new_n255), .ZN(new_n838));
  NOR4_X1   g0638(.A1(new_n834), .A2(new_n836), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n830), .A2(new_n831), .A3(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(G283), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n773), .A2(new_n841), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n385), .B1(new_n777), .B2(new_n567), .C1(new_n780), .C2(new_n778), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n842), .B(new_n843), .C1(G303), .C2(new_n783), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n785), .A2(new_n311), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n835), .A2(new_n222), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n845), .B(new_n846), .C1(G311), .C2(new_n788), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n844), .B(new_n847), .C1(new_n793), .C2(new_n477), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n822), .B1(new_n840), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n754), .A2(new_n755), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n821), .B(new_n849), .C1(new_n278), .C2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n756), .B2(new_n814), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n820), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(G384));
  NOR2_X1   g0654(.A1(new_n735), .A2(new_n208), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT39), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT38), .ZN(new_n857));
  INV_X1    g0657(.A(new_n437), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n443), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n667), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n453), .A2(new_n454), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n861), .B1(new_n862), .B2(new_n657), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n450), .A2(new_n859), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n864), .A2(new_n440), .A3(new_n861), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT37), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n447), .B1(new_n450), .B2(new_n860), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(new_n868), .A3(new_n440), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n857), .B1(new_n863), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n866), .A2(new_n869), .ZN(new_n872));
  OAI211_X1 g0672(.A(KEYINPUT38), .B(new_n872), .C1(new_n455), .C2(new_n861), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n856), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n869), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n440), .B1(new_n650), .B2(new_n651), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT99), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n447), .A2(new_n860), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT99), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n879), .B(new_n440), .C1(new_n650), .C2(new_n651), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n875), .B1(new_n881), .B2(KEYINPUT37), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n652), .A2(new_n655), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n442), .A2(new_n445), .A3(KEYINPUT100), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT100), .B1(new_n442), .B2(new_n445), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n878), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n857), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n873), .A2(new_n856), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n874), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n374), .A2(new_n669), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT98), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n871), .A2(new_n894), .A3(new_n873), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n894), .B1(new_n871), .B2(new_n873), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n322), .A2(new_n672), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n817), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n373), .A2(new_n669), .ZN(new_n900));
  INV_X1    g0700(.A(new_n357), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n354), .B2(new_n355), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n900), .B1(new_n383), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n900), .B1(new_n377), .B2(new_n380), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n358), .B2(new_n373), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n899), .A2(new_n907), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n897), .A2(new_n908), .B1(new_n883), .B2(new_n860), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n893), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n456), .B1(new_n729), .B2(new_n731), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n911), .A2(new_n662), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT101), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n910), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n814), .B1(new_n903), .B2(new_n905), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n714), .B1(new_n706), .B2(new_n708), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT90), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n917), .B(new_n696), .C1(new_n693), .C2(new_n694), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n703), .A2(new_n705), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n707), .A2(KEYINPUT90), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n672), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n712), .B(new_n916), .C1(new_n922), .C2(KEYINPUT31), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT103), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT103), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n711), .A2(new_n925), .A3(new_n712), .A4(new_n916), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n915), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n895), .B2(new_n896), .ZN(new_n928));
  XNOR2_X1  g0728(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n888), .A2(new_n873), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n932), .B(new_n915), .C1(new_n926), .C2(new_n924), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n928), .A2(new_n930), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n456), .B1(new_n926), .B2(new_n924), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n678), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n934), .B2(new_n935), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n855), .B1(new_n914), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n914), .B2(new_n937), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n594), .A2(KEYINPUT35), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n594), .A2(KEYINPUT35), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n940), .A2(G116), .A3(new_n218), .A4(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT36), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n216), .A2(G77), .A3(new_n391), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(G50), .B2(new_n202), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(G1), .A3(new_n734), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n939), .A2(new_n943), .A3(new_n946), .ZN(G367));
  NAND2_X1  g0747(.A1(new_n601), .A2(new_n669), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n639), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n628), .A2(new_n669), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n951), .A2(new_n555), .A3(new_n670), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n952), .A2(KEYINPUT42), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n622), .B1(new_n949), .B2(new_n642), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n952), .A2(KEYINPUT42), .B1(new_n672), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n474), .A2(new_n669), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n637), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n636), .B2(new_n956), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n953), .A2(new_n955), .B1(KEYINPUT43), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n959), .B(new_n960), .Z(new_n961));
  INV_X1    g0761(.A(new_n951), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n683), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n961), .B(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n686), .B(KEYINPUT41), .Z(new_n965));
  OAI21_X1  g0765(.A(new_n671), .B1(new_n677), .B2(new_n670), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n682), .A2(KEYINPUT105), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n682), .B(KEYINPUT105), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n968), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n970), .A2(new_n729), .A3(new_n731), .A4(new_n722), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(KEYINPUT44), .B1(new_n962), .B2(new_n674), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n962), .A2(KEYINPUT44), .A3(new_n674), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n977));
  NAND3_X1  g0777(.A1(new_n675), .A2(new_n951), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n977), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n962), .B2(new_n674), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n976), .A2(new_n683), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n683), .ZN(new_n982));
  INV_X1    g0782(.A(new_n975), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(new_n973), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n978), .A2(new_n980), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n972), .A2(KEYINPUT106), .A3(new_n981), .A4(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT106), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n981), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n988), .B1(new_n989), .B2(new_n971), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n965), .B1(new_n991), .B2(new_n732), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n964), .B1(new_n992), .B2(new_n737), .ZN(new_n993));
  INV_X1    g0793(.A(new_n303), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n759), .B1(new_n685), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n746), .A2(new_n233), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n821), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n786), .A2(G116), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT46), .ZN(new_n999));
  INV_X1    g0799(.A(G317), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n385), .B1(new_n787), .B2(new_n1000), .C1(new_n780), .C2(new_n559), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n772), .A2(G294), .B1(new_n783), .B2(G311), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n311), .B2(new_n777), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1001), .B(new_n1003), .C1(G97), .C2(new_n769), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n999), .B(new_n1004), .C1(new_n793), .C2(new_n841), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n793), .A2(new_n255), .B1(new_n396), .B2(new_n773), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT108), .Z(new_n1007));
  OAI22_X1  g0807(.A1(new_n826), .A2(new_n802), .B1(new_n780), .B2(new_n823), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n777), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1008), .B1(G68), .B2(new_n1009), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1010), .A2(KEYINPUT107), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(KEYINPUT107), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n769), .A2(G77), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n275), .B1(new_n787), .B2(new_n825), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n786), .B2(G58), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1005), .B1(new_n1007), .B2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT47), .Z(new_n1018));
  OAI221_X1 g0818(.A(new_n997), .B1(new_n761), .B2(new_n958), .C1(new_n1018), .C2(new_n822), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n993), .A2(new_n1019), .ZN(G387));
  NOR2_X1   g0820(.A1(new_n972), .A2(new_n687), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n732), .B2(new_n970), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n970), .A2(new_n737), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n768), .A2(G68), .B1(G97), .B2(new_n769), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n275), .B1(new_n780), .B2(new_n255), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n396), .A2(new_n802), .B1(new_n773), .B2(new_n263), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(G150), .C2(new_n796), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n786), .A2(G77), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n501), .A2(new_n1009), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1024), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(G311), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n1031), .A2(new_n773), .B1(new_n780), .B2(new_n1000), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G322), .B2(new_n783), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n793), .B2(new_n559), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT48), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n785), .A2(new_n778), .B1(new_n841), .B2(new_n777), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(KEYINPUT49), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n275), .B1(new_n796), .B2(G326), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(new_n477), .C2(new_n835), .ZN(new_n1041));
  AOI21_X1  g0841(.A(KEYINPUT49), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1030), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n754), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n688), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n743), .A2(new_n1045), .B1(new_n311), .B2(new_n685), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n238), .A2(new_n287), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n435), .A2(new_n255), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT50), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n688), .B(new_n287), .C1(new_n202), .C2(new_n278), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n746), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1046), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n821), .B1(new_n1052), .B2(new_n758), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1044), .B(new_n1053), .C1(new_n677), .C2(new_n761), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1022), .A2(new_n1023), .A3(new_n1054), .ZN(G393));
  INV_X1    g0855(.A(KEYINPUT112), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT109), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n986), .B2(new_n981), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n981), .A2(new_n1057), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n1058), .A2(new_n1059), .A3(new_n736), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n962), .A2(new_n757), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n747), .A2(new_n242), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n758), .B1(new_n567), .B2(new_n212), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n738), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT110), .Z(new_n1065));
  AOI22_X1  g0865(.A1(new_n768), .A2(G294), .B1(G107), .B2(new_n769), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n1000), .A2(new_n802), .B1(new_n780), .B2(new_n1031), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT52), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n385), .B1(new_n787), .B2(new_n781), .C1(new_n773), .C2(new_n559), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G116), .B2(new_n1009), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n786), .A2(G283), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1066), .A2(new_n1068), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n275), .B1(new_n787), .B2(new_n826), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1073), .B(new_n846), .C1(G68), .C2(new_n786), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT111), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n823), .A2(new_n802), .B1(new_n780), .B2(new_n396), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT51), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1009), .A2(G77), .B1(G50), .B2(new_n772), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(new_n793), .C2(new_n263), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1072), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1065), .B1(new_n1080), .B2(new_n754), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1061), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1056), .B1(new_n1060), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n989), .A2(KEYINPUT109), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n981), .A2(new_n1057), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g0887(.A(KEYINPUT112), .B(new_n1082), .C1(new_n1087), .C2(new_n736), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n687), .B1(new_n1087), .B2(new_n971), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1084), .A2(new_n1088), .B1(new_n1089), .B2(new_n991), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(G390));
  NAND2_X1  g0891(.A1(new_n908), .A2(new_n892), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n890), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n727), .A2(new_n814), .A3(new_n672), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n898), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n891), .B1(new_n1095), .B2(new_n907), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n931), .A2(new_n1096), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n713), .A2(new_n721), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1098), .A2(new_n907), .A3(G330), .A4(new_n814), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1093), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n890), .A2(new_n1092), .B1(new_n931), .B2(new_n1096), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n678), .B1(new_n924), .B2(new_n926), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n915), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1100), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1102), .A2(new_n457), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n912), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n906), .B1(new_n722), .B2(new_n815), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n899), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1095), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n678), .B(new_n815), .C1(new_n924), .C2(new_n926), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1099), .B(new_n1111), .C1(new_n1112), .C2(new_n907), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1107), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1105), .A2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1114), .B(new_n1100), .C1(new_n1101), .C2(new_n1104), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n686), .A3(new_n1117), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1105), .A2(new_n736), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n890), .A2(new_n755), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n850), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n738), .B1(new_n1121), .B2(new_n435), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT113), .Z(new_n1123));
  OAI21_X1  g0923(.A(new_n385), .B1(new_n780), .B2(new_n477), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n773), .A2(new_n311), .B1(new_n802), .B2(new_n841), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1124), .B(new_n1125), .C1(G77), .C2(new_n1009), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n801), .B(new_n836), .C1(G294), .C2(new_n788), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1126), .B(new_n1127), .C1(new_n793), .C2(new_n567), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT54), .B(G143), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n793), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n785), .A2(new_n823), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT53), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n275), .B1(new_n780), .B2(new_n833), .ZN(new_n1133));
  INV_X1    g0933(.A(G128), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n773), .A2(new_n825), .B1(new_n802), .B2(new_n1134), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1133), .B(new_n1135), .C1(G159), .C2(new_n1009), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n788), .A2(G125), .B1(G50), .B2(new_n769), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1132), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1128), .B1(new_n1130), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1123), .B1(new_n1139), .B2(new_n754), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1120), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1118), .A2(new_n1119), .A3(new_n1141), .ZN(G378));
  INV_X1    g0942(.A(new_n910), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n678), .B1(new_n928), .B2(new_n930), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT118), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n931), .A2(new_n933), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1145), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n302), .A2(new_n328), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n270), .A2(new_n860), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1149), .B(new_n1150), .ZN(new_n1151));
  XOR2_X1   g0951(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1152));
  XNOR2_X1  g0952(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n1147), .A2(new_n1148), .A3(new_n1153), .ZN(new_n1154));
  AND4_X1   g0954(.A1(new_n1145), .A2(new_n1144), .A3(new_n1146), .A4(new_n1153), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1143), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1153), .B1(new_n1157), .B2(KEYINPUT118), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1155), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n910), .A3(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1156), .A2(new_n737), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1153), .A2(new_n755), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n738), .B1(new_n1121), .B2(G50), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n275), .A2(G41), .ZN(new_n1166));
  AOI211_X1 g0966(.A(G50), .B(new_n1166), .C1(new_n260), .C2(new_n286), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1166), .B1(new_n202), .B2(new_n777), .C1(new_n311), .C2(new_n780), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n769), .A2(G58), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1028), .B(new_n1169), .C1(new_n832), .C2(new_n841), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1168), .B(new_n1170), .C1(G116), .C2(new_n783), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n768), .A2(new_n501), .B1(G97), .B2(new_n772), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT114), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1171), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  XOR2_X1   g0976(.A(KEYINPUT115), .B(KEYINPUT58), .Z(new_n1177));
  AOI21_X1  g0977(.A(new_n1167), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n785), .A2(new_n1129), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT116), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n773), .A2(new_n833), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n780), .A2(new_n1134), .B1(new_n777), .B2(new_n823), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(G125), .C2(new_n783), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n768), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1180), .B(new_n1183), .C1(new_n825), .C2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1187));
  AOI211_X1 g0987(.A(G33), .B(G41), .C1(new_n796), .C2(G124), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n396), .B2(new_n835), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT117), .Z(new_n1190));
  NAND2_X1  g0990(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1178), .B1(new_n1186), .B2(new_n1191), .C1(new_n1177), .C2(new_n1176), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1165), .B1(new_n1192), .B2(new_n754), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1164), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1163), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT119), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1163), .A2(KEYINPUT119), .A3(new_n1194), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1107), .B(KEYINPUT120), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1117), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1156), .A2(new_n1162), .A3(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT57), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1203), .B1(new_n1117), .B2(new_n1200), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1156), .A2(new_n1162), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT121), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT121), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1156), .A2(new_n1205), .A3(new_n1162), .A4(new_n1208), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1204), .A2(new_n1207), .A3(new_n686), .A4(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1199), .A2(new_n1210), .ZN(G375));
  AOI21_X1  g1011(.A(new_n821), .B1(new_n850), .B2(new_n202), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n385), .B1(new_n780), .B2(new_n841), .C1(new_n778), .C2(new_n802), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G97), .A2(new_n786), .B1(new_n788), .B2(G303), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(new_n1013), .A3(new_n1029), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1213), .B(new_n1215), .C1(G116), .C2(new_n772), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n828), .A2(G107), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n275), .B1(new_n780), .B2(new_n825), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n833), .A2(new_n802), .B1(new_n773), .B2(new_n1129), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(G50), .C2(new_n1009), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n1184), .A2(new_n823), .B1(new_n396), .B2(new_n785), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1169), .B1(new_n832), .B2(new_n1134), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1216), .A2(new_n1217), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1212), .B1(new_n822), .B2(new_n1224), .C1(new_n907), .C2(new_n756), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1226), .B1(new_n1227), .B2(new_n737), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1114), .A2(new_n965), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1110), .A2(new_n1107), .A3(new_n1113), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1228), .B1(new_n1229), .B2(new_n1231), .ZN(G381));
  INV_X1    g1032(.A(G378), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1199), .A2(new_n1233), .A3(new_n1210), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n993), .A2(new_n1090), .A3(new_n1019), .ZN(new_n1236));
  NOR4_X1   g1036(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(G407));
  OAI211_X1 g1038(.A(G407), .B(G213), .C1(G343), .C2(new_n1234), .ZN(G409));
  XNOR2_X1  g1039(.A(G393), .B(new_n808), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1090), .B1(new_n993), .B2(new_n1019), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1241), .B1(new_n1236), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT125), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(KEYINPUT125), .B(new_n1241), .C1(new_n1236), .C2(new_n1242), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G387), .A2(G390), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n993), .A2(new_n1090), .A3(new_n1019), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n1249), .A3(new_n1240), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT124), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT124), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1248), .A2(new_n1252), .A3(new_n1249), .A4(new_n1240), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1247), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT61), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT126), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT126), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n1258), .B(KEYINPUT61), .C1(new_n1247), .C2(new_n1254), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n668), .A2(G213), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1210), .A2(G378), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1202), .A2(new_n965), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1233), .B1(new_n1264), .B2(new_n1195), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1262), .B1(new_n1263), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT122), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1230), .A2(new_n1267), .A3(KEYINPUT60), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT60), .B1(new_n1230), .B2(new_n1267), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n686), .B(new_n1115), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1228), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n853), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(G384), .A3(new_n1228), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1266), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1273), .B(new_n1274), .C1(KEYINPUT123), .C2(new_n1261), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1262), .A2(G2897), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1280), .B(new_n1281), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1266), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1266), .A2(KEYINPUT63), .A3(new_n1276), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1260), .A2(new_n1279), .A3(new_n1283), .A4(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1266), .A2(new_n1286), .A3(new_n1276), .ZN(new_n1287));
  XOR2_X1   g1087(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1288));
  OAI21_X1  g1088(.A(new_n1288), .B1(new_n1266), .B2(new_n1282), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1286), .B1(new_n1266), .B2(new_n1276), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1287), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1285), .B1(new_n1291), .B2(new_n1255), .ZN(G405));
  NAND2_X1  g1092(.A1(G375), .A2(new_n1233), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1263), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1276), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1255), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1293), .A2(new_n1263), .A3(new_n1275), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1296), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(G402));
endmodule


