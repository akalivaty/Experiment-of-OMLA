//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1328, new_n1329;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XOR2_X1   g0026(.A(G226), .B(G232), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n230), .B(new_n231), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT66), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n232), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  OR3_X1    g0046(.A1(new_n207), .A2(KEYINPUT68), .A3(G1), .ZN(new_n247));
  OAI21_X1  g0047(.A(KEYINPUT68), .B1(new_n207), .B2(G1), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n215), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n252), .A2(new_n257), .B1(new_n254), .B2(new_n251), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(KEYINPUT7), .B1(new_n261), .B2(new_n207), .ZN(new_n262));
  OR2_X1    g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  AND4_X1   g0064(.A1(KEYINPUT7), .A2(new_n263), .A3(new_n207), .A4(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(G68), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G159), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(G58), .A2(G68), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G58), .A2(G68), .ZN(new_n272));
  OAI21_X1  g0072(.A(G20), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT76), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI211_X1 g0075(.A(KEYINPUT76), .B(G20), .C1(new_n271), .C2(new_n272), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n270), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n266), .A2(new_n277), .A3(KEYINPUT16), .ZN(new_n278));
  AOI21_X1  g0078(.A(KEYINPUT16), .B1(new_n266), .B2(new_n277), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT77), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n256), .B(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n279), .A2(new_n280), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n258), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(G1), .A3(G13), .ZN(new_n285));
  INV_X1    g0085(.A(G226), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G1698), .ZN(new_n287));
  OAI221_X1 g0087(.A(new_n287), .B1(G223), .B2(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G87), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n285), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G41), .ZN(new_n291));
  INV_X1    g0091(.A(G45), .ZN(new_n292));
  AOI21_X1  g0092(.A(G1), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(new_n285), .A3(G274), .ZN(new_n294));
  INV_X1    g0094(.A(G232), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n285), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n294), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n290), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT78), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT78), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(new_n290), .B2(new_n298), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  INV_X1    g0104(.A(G179), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n303), .A2(new_n304), .B1(new_n305), .B2(new_n299), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n283), .A2(KEYINPUT18), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT79), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n283), .A2(KEYINPUT79), .A3(new_n306), .A4(KEYINPUT18), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n283), .A2(new_n306), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT18), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n309), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT17), .ZN(new_n315));
  INV_X1    g0115(.A(G200), .ZN(new_n316));
  INV_X1    g0116(.A(G190), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n303), .A2(new_n316), .B1(new_n317), .B2(new_n299), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n315), .B1(new_n283), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n302), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n290), .A2(new_n298), .A3(new_n301), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n316), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n299), .A2(new_n317), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n266), .A2(new_n277), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT16), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT77), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n278), .A2(new_n256), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n279), .A2(new_n280), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n324), .A2(new_n331), .A3(KEYINPUT17), .A4(new_n258), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n319), .A2(KEYINPUT80), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(KEYINPUT80), .B1(new_n319), .B2(new_n332), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n314), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n337));
  INV_X1    g0137(.A(G150), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n207), .A2(G33), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n337), .B1(new_n338), .B2(new_n268), .C1(new_n339), .C2(new_n251), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n340), .A2(new_n256), .B1(new_n201), .B2(new_n254), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT69), .B1(new_n250), .B2(new_n201), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n257), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n250), .A2(KEYINPUT69), .A3(new_n201), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n341), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT9), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n263), .A2(new_n264), .ZN(new_n348));
  INV_X1    g0148(.A(G1698), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(G222), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G77), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(G1698), .ZN(new_n352));
  INV_X1    g0152(.A(G223), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n350), .B1(new_n351), .B2(new_n348), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n294), .ZN(new_n357));
  INV_X1    g0157(.A(new_n297), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n357), .B1(G226), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G200), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n347), .B(new_n361), .C1(new_n317), .C2(new_n360), .ZN(new_n362));
  NAND2_X1  g0162(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n345), .B2(new_n346), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n360), .A2(new_n304), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n356), .A2(new_n305), .A3(new_n359), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(new_n345), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n348), .A2(G232), .A3(new_n349), .ZN(new_n371));
  INV_X1    g0171(.A(G107), .ZN(new_n372));
  INV_X1    g0172(.A(G238), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n371), .B1(new_n372), .B2(new_n348), .C1(new_n352), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n355), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n357), .B1(G244), .B2(new_n358), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n305), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n251), .A2(new_n268), .B1(new_n207), .B2(new_n351), .ZN(new_n380));
  XNOR2_X1  g0180(.A(KEYINPUT15), .B(G87), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(new_n339), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n256), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n250), .A2(new_n351), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n384), .A2(new_n257), .B1(new_n351), .B2(new_n254), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n377), .A2(new_n304), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n379), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT70), .B1(new_n378), .B2(new_n316), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n317), .B2(new_n377), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n385), .A2(new_n383), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n377), .A2(new_n317), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(KEYINPUT70), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n388), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n336), .A2(new_n367), .A3(new_n370), .A4(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n286), .A2(new_n349), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n295), .A2(G1698), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n397), .B(new_n398), .C1(new_n259), .C2(new_n260), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT72), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G97), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n400), .B1(new_n399), .B2(new_n401), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n403), .A2(new_n404), .A3(new_n285), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n357), .B1(G238), .B2(new_n358), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT13), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT13), .ZN(new_n409));
  OR2_X1    g0209(.A1(new_n404), .A2(new_n285), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n409), .B(new_n406), .C1(new_n410), .C2(new_n403), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n411), .A3(KEYINPUT73), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT73), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n413), .B(KEYINPUT13), .C1(new_n405), .C2(new_n407), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n412), .A2(G169), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT14), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT74), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n408), .A2(new_n411), .A3(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n405), .A2(new_n407), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(KEYINPUT74), .A3(new_n409), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G179), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT14), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n412), .A2(new_n423), .A3(G169), .A4(new_n414), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n416), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G68), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n254), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT12), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n267), .A2(G50), .B1(G20), .B2(new_n426), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n351), .B2(new_n339), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(KEYINPUT11), .A3(new_n256), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n257), .A2(new_n249), .A3(G68), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n428), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(KEYINPUT11), .B1(new_n430), .B2(new_n256), .ZN(new_n434));
  OR2_X1    g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n425), .A2(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n412), .A2(G200), .A3(new_n414), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n317), .B1(new_n418), .B2(new_n420), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n437), .A2(new_n438), .A3(new_n435), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n441), .A2(KEYINPUT75), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(KEYINPUT75), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n396), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  OAI211_X1 g0244(.A(G250), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT83), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT83), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n348), .A2(new_n447), .A3(G250), .A4(G1698), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(G244), .B(new_n349), .C1(new_n259), .C2(new_n260), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT4), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n348), .A2(KEYINPUT4), .A3(G244), .A4(new_n349), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G283), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT82), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT82), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(G33), .A3(G283), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n452), .A2(new_n453), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n355), .B1(new_n449), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n292), .A2(G1), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT5), .B(G41), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n355), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G257), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n462), .A2(G274), .A3(new_n285), .A4(new_n461), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n460), .A2(new_n467), .A3(G190), .ZN(new_n468));
  INV_X1    g0268(.A(G97), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n254), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G33), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G1), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n254), .A2(new_n256), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n470), .B1(new_n474), .B2(new_n469), .ZN(new_n475));
  OAI21_X1  g0275(.A(G107), .B1(new_n262), .B2(new_n265), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n469), .A2(new_n372), .A3(KEYINPUT6), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT6), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G97), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n372), .A2(KEYINPUT81), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT81), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G107), .ZN(new_n482));
  AND4_X1   g0282(.A1(new_n477), .A2(new_n479), .A3(new_n480), .A4(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n477), .A2(new_n479), .B1(new_n480), .B2(new_n482), .ZN(new_n484));
  OAI21_X1  g0284(.A(G20), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n267), .A2(G77), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n476), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n475), .B1(new_n487), .B2(new_n256), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n468), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n316), .B1(new_n460), .B2(new_n467), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT84), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n460), .A2(new_n467), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G200), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT84), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n493), .A2(new_n494), .A3(new_n488), .A4(new_n468), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT85), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n446), .A2(new_n448), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n498), .A2(new_n453), .A3(new_n458), .A4(new_n452), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n466), .B1(new_n499), .B2(new_n355), .ZN(new_n500));
  INV_X1    g0300(.A(new_n256), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n477), .A2(new_n479), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n480), .A2(new_n482), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n477), .A2(new_n479), .A3(new_n480), .A4(new_n482), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n506), .A2(G20), .B1(G77), .B2(new_n267), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n501), .B1(new_n507), .B2(new_n476), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n500), .A2(G169), .B1(new_n508), .B2(new_n475), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n492), .A2(G179), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n497), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n492), .A2(new_n304), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n500), .A2(new_n305), .ZN(new_n513));
  INV_X1    g0313(.A(new_n488), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n512), .A2(new_n513), .A3(new_n514), .A4(KEYINPUT85), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n496), .A2(new_n511), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n373), .A2(new_n349), .ZN(new_n517));
  INV_X1    g0317(.A(G244), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G1698), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n517), .B(new_n519), .C1(new_n259), .C2(new_n260), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G116), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT86), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n520), .A2(KEYINPUT86), .A3(new_n521), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n285), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n285), .A2(G274), .A3(new_n461), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n206), .A2(G45), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n285), .A2(G250), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(G169), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n348), .A2(new_n207), .A3(G68), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT19), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n207), .B1(new_n401), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(G87), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(new_n469), .A3(new_n372), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n534), .B1(new_n339), .B2(new_n469), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n533), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(new_n256), .B1(new_n254), .B2(new_n381), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n381), .B2(new_n474), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n520), .A2(KEYINPUT86), .A3(new_n521), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT86), .B1(new_n520), .B2(new_n521), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n355), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n530), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n305), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n532), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n545), .A2(new_n546), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G200), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n473), .A2(G87), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n541), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n545), .A2(G190), .A3(new_n546), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT87), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n545), .A2(KEYINPUT87), .A3(G190), .A4(new_n546), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT88), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n554), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n557), .A2(KEYINPUT88), .A3(new_n558), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n549), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n253), .A2(G116), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n473), .B2(G116), .ZN(new_n565));
  AOI21_X1  g0365(.A(G20), .B1(new_n471), .B2(G97), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n458), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G116), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n255), .A2(new_n215), .B1(G20), .B2(new_n568), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n567), .A2(new_n569), .A3(KEYINPUT20), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT20), .B1(new_n567), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n565), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT21), .ZN(new_n573));
  AND2_X1   g0373(.A1(KEYINPUT5), .A2(G41), .ZN(new_n574));
  NOR2_X1   g0374(.A1(KEYINPUT5), .A2(G41), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n461), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(G270), .A3(new_n285), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n577), .A2(new_n465), .ZN(new_n578));
  OAI211_X1 g0378(.A(G264), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n579));
  OAI211_X1 g0379(.A(G257), .B(new_n349), .C1(new_n259), .C2(new_n260), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n263), .A2(G303), .A3(new_n264), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n355), .ZN(new_n583));
  AOI211_X1 g0383(.A(new_n573), .B(new_n304), .C1(new_n578), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n578), .A2(new_n583), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n585), .A2(new_n305), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n572), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT89), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n304), .B1(new_n578), .B2(new_n583), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n572), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n588), .B1(new_n590), .B2(new_n573), .ZN(new_n591));
  AOI211_X1 g0391(.A(KEYINPUT89), .B(KEYINPUT21), .C1(new_n589), .C2(new_n572), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n348), .A2(G257), .A3(G1698), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n348), .A2(G250), .A3(new_n349), .ZN(new_n595));
  INV_X1    g0395(.A(G294), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n594), .B(new_n595), .C1(new_n471), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n355), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n463), .A2(G264), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n465), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n304), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n597), .A2(new_n355), .B1(G264), .B2(new_n463), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(new_n305), .A3(new_n465), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n521), .A2(G20), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT23), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n207), .B2(G107), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n372), .A2(KEYINPUT23), .A3(G20), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n207), .B(G87), .C1(new_n259), .C2(new_n260), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n609), .A2(KEYINPUT22), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n609), .A2(KEYINPUT22), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n608), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT24), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT24), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n614), .B(new_n608), .C1(new_n610), .C2(new_n611), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n501), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT25), .B1(new_n254), .B2(new_n372), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n254), .A2(KEYINPUT25), .A3(new_n372), .ZN(new_n618));
  OAI22_X1  g0418(.A1(new_n474), .A2(new_n372), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n601), .B(new_n603), .C1(new_n616), .C2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n593), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n316), .B1(new_n578), .B2(new_n583), .ZN(new_n623));
  INV_X1    g0423(.A(new_n585), .ZN(new_n624));
  AOI211_X1 g0424(.A(new_n572), .B(new_n623), .C1(G190), .C2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n600), .A2(new_n317), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(G200), .B2(new_n600), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n616), .A2(new_n619), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n563), .A2(new_n622), .A3(new_n629), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n444), .A2(new_n516), .A3(new_n630), .ZN(G372));
  INV_X1    g0431(.A(new_n444), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n511), .A2(new_n515), .ZN(new_n633));
  INV_X1    g0433(.A(new_n549), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n559), .A2(new_n560), .ZN(new_n635));
  INV_X1    g0435(.A(new_n554), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n562), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n633), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT26), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n530), .A2(KEYINPUT90), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT90), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n527), .A2(new_n529), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n304), .B1(new_n526), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n644), .A2(new_n542), .A3(new_n547), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n541), .A2(new_n552), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n647), .B1(new_n557), .B2(new_n558), .ZN(new_n648));
  OAI21_X1  g0448(.A(G200), .B1(new_n526), .B2(new_n643), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT91), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n545), .A2(new_n640), .A3(new_n642), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(KEYINPUT91), .A3(G200), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n646), .B1(new_n648), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT26), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n509), .A2(new_n510), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n639), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n620), .B(new_n587), .C1(new_n591), .C2(new_n592), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n627), .A2(new_n628), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(new_n655), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n645), .B1(new_n663), .B2(new_n516), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n632), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n370), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n440), .A2(new_n388), .B1(new_n425), .B2(new_n435), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n333), .A2(new_n334), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n283), .A2(KEYINPUT18), .A3(new_n306), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT18), .B1(new_n283), .B2(new_n306), .ZN(new_n672));
  OAI22_X1  g0472(.A1(new_n669), .A2(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n668), .B1(new_n673), .B2(new_n367), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n667), .A2(new_n674), .ZN(G369));
  NAND3_X1  g0475(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT92), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n677), .B(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G213), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n676), .B2(KEYINPUT27), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G343), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT93), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n572), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(new_n593), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(new_n625), .ZN(new_n687));
  INV_X1    g0487(.A(G330), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n684), .B1(new_n616), .B2(new_n619), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n621), .B1(new_n690), .B2(new_n662), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n684), .A2(new_n620), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n684), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n593), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT94), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n692), .B1(new_n697), .B2(new_n693), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n694), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n210), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n537), .A2(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n213), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n648), .A2(new_n654), .ZN(new_n707));
  AND4_X1   g0507(.A1(KEYINPUT26), .A2(new_n707), .A3(new_n657), .A4(new_n645), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n656), .B2(new_n638), .ZN(new_n709));
  OAI211_X1 g0509(.A(KEYINPUT29), .B(new_n695), .C1(new_n709), .C2(new_n664), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n684), .B1(new_n660), .B2(new_n665), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n710), .B1(new_n711), .B2(KEYINPUT29), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n563), .A2(new_n629), .ZN(new_n713));
  INV_X1    g0513(.A(new_n516), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n713), .A2(new_n714), .A3(new_n622), .A4(new_n695), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n500), .A2(new_n586), .A3(new_n531), .A4(new_n602), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n602), .A2(new_n546), .A3(new_n545), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n720), .A2(KEYINPUT30), .A3(new_n500), .A4(new_n586), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n624), .A2(G179), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n722), .A2(new_n652), .A3(new_n492), .A4(new_n600), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n719), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n716), .B1(new_n724), .B2(new_n684), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n724), .A2(new_n716), .A3(new_n684), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n688), .B1(new_n715), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n712), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n706), .B1(new_n732), .B2(G1), .ZN(G364));
  NOR2_X1   g0533(.A1(G13), .A2(G33), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n687), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n215), .B1(G20), .B2(new_n304), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n207), .A2(new_n317), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n305), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n207), .A2(G190), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI22_X1  g0546(.A1(G58), .A2(new_n743), .B1(new_n746), .B2(G77), .ZN(new_n747));
  NAND3_X1  g0547(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n317), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n747), .B1(new_n201), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT95), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n316), .A2(G179), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n744), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n372), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n740), .A2(new_n753), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n261), .B(new_n755), .C1(G87), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G179), .A2(G200), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n207), .B1(new_n759), .B2(G190), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n469), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n748), .A2(G190), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n761), .B1(new_n762), .B2(G68), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n744), .A2(new_n759), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n269), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT32), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n752), .A2(new_n758), .A3(new_n763), .A4(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G322), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n261), .B1(new_n742), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n760), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n769), .B1(G294), .B2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n764), .ZN(new_n772));
  AOI22_X1  g0572(.A1(G311), .A2(new_n746), .B1(new_n772), .B2(G329), .ZN(new_n773));
  INV_X1    g0573(.A(new_n754), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G303), .A2(new_n757), .B1(new_n774), .B2(G283), .ZN(new_n775));
  XOR2_X1   g0575(.A(KEYINPUT96), .B(G326), .Z(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(KEYINPUT33), .B(G317), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n777), .A2(new_n749), .B1(new_n762), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n771), .A2(new_n773), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n739), .B1(new_n767), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G13), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n206), .B1(new_n783), .B2(G45), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n701), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n210), .A2(new_n348), .ZN(new_n787));
  INV_X1    g0587(.A(G355), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n787), .A2(new_n788), .B1(G116), .B2(new_n210), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n242), .A2(new_n292), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n700), .A2(new_n348), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(new_n292), .B2(new_n214), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n789), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n736), .A2(new_n738), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n786), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  OR3_X1    g0597(.A1(new_n737), .A2(new_n781), .A3(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n689), .ZN(new_n799));
  INV_X1    g0599(.A(new_n786), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n687), .A2(new_n688), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(G396));
  AOI22_X1  g0604(.A1(new_n390), .A2(new_n393), .B1(new_n391), .B2(new_n684), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n388), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n387), .A2(new_n684), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n711), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n808), .B(new_n695), .C1(new_n659), .C2(new_n664), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n786), .B1(new_n811), .B2(new_n730), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n730), .B2(new_n811), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n738), .A2(new_n734), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n800), .B1(new_n351), .B2(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G143), .A2(new_n743), .B1(new_n746), .B2(G159), .ZN(new_n816));
  INV_X1    g0616(.A(G137), .ZN(new_n817));
  INV_X1    g0617(.A(new_n762), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n816), .B1(new_n750), .B2(new_n817), .C1(new_n338), .C2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT34), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n348), .B1(new_n754), .B2(new_n426), .ZN(new_n823));
  INV_X1    g0623(.A(G132), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n756), .A2(new_n201), .B1(new_n764), .B2(new_n824), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n823), .B(new_n825), .C1(G58), .C2(new_n770), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n821), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n261), .B1(new_n756), .B2(new_n372), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n761), .B(new_n828), .C1(G303), .C2(new_n749), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n742), .A2(new_n596), .B1(new_n745), .B2(new_n568), .ZN(new_n830));
  INV_X1    g0630(.A(G311), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n754), .A2(new_n536), .B1(new_n764), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G283), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n818), .A2(KEYINPUT97), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n818), .A2(KEYINPUT97), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n829), .B(new_n833), .C1(new_n834), .C2(new_n837), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n827), .A2(new_n838), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n815), .B1(new_n739), .B2(new_n839), .C1(new_n808), .C2(new_n735), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n813), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G384));
  NOR2_X1   g0642(.A1(new_n783), .A2(new_n206), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n684), .A2(new_n435), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n436), .A2(new_n440), .A3(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n435), .B(new_n684), .C1(new_n439), .C2(new_n425), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n807), .B(new_n806), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n715), .A2(new_n728), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n847), .A2(KEYINPUT40), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n324), .A2(new_n331), .A3(new_n258), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n329), .A2(new_n327), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n258), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT99), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n306), .A2(new_n682), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n283), .A2(new_n682), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT37), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n311), .A2(new_n857), .A3(new_n850), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n682), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n853), .A2(new_n861), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n335), .A2(KEYINPUT100), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT100), .B1(new_n335), .B2(new_n862), .ZN(new_n864));
  OAI211_X1 g0664(.A(KEYINPUT38), .B(new_n860), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n857), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n671), .A2(new_n672), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n319), .A2(new_n332), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n311), .A2(new_n857), .A3(new_n850), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n859), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT101), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT101), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n876), .B(KEYINPUT38), .C1(new_n869), .C2(new_n872), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n849), .B1(new_n865), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n847), .A2(new_n848), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n335), .A2(new_n862), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT100), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n335), .A2(KEYINPUT100), .A3(new_n862), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n886), .B2(new_n860), .ZN(new_n887));
  INV_X1    g0687(.A(new_n865), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n881), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  XOR2_X1   g0689(.A(KEYINPUT103), .B(KEYINPUT40), .Z(new_n890));
  AOI21_X1  g0690(.A(new_n879), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n891), .B(KEYINPUT104), .Z(new_n892));
  NAND2_X1  g0692(.A1(new_n632), .A2(new_n848), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(G330), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n865), .A2(new_n878), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT39), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n874), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(KEYINPUT39), .A3(new_n865), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n436), .A2(new_n684), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n807), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n810), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n845), .A2(new_n846), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT98), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n908), .A2(KEYINPUT98), .A3(new_n909), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n912), .B(new_n913), .C1(new_n888), .C2(new_n887), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n867), .A2(new_n861), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n906), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n674), .B1(new_n444), .B2(new_n712), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT102), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n917), .B(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n843), .B1(new_n896), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n920), .B2(new_n896), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n216), .A2(G116), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n506), .B2(KEYINPUT35), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(KEYINPUT35), .B2(new_n506), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT36), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n213), .A2(new_n271), .A3(new_n351), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n426), .A2(G50), .ZN(new_n928));
  OAI211_X1 g0728(.A(G1), .B(new_n782), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n922), .A2(new_n926), .A3(new_n929), .ZN(G367));
  OAI21_X1  g0730(.A(new_n714), .B1(new_n488), .B2(new_n695), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n657), .A2(new_n684), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(new_n693), .A3(new_n697), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT42), .Z(new_n935));
  INV_X1    g0735(.A(new_n933), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n936), .A2(new_n620), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n695), .B1(new_n937), .B2(new_n633), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n695), .A2(new_n553), .ZN(new_n939));
  MUX2_X1   g0739(.A(new_n655), .B(new_n646), .S(new_n939), .Z(new_n940));
  AOI22_X1  g0740(.A1(new_n935), .A2(new_n938), .B1(KEYINPUT43), .B2(new_n940), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n694), .A2(new_n936), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n943), .B(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n701), .B(KEYINPUT41), .Z(new_n946));
  NAND2_X1  g0746(.A1(new_n698), .A2(new_n933), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT45), .Z(new_n948));
  NOR2_X1   g0748(.A1(new_n698), .A2(new_n933), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT44), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(new_n694), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n697), .B(new_n693), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(new_n689), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n732), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n946), .B1(new_n957), .B2(new_n732), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n945), .B1(new_n958), .B2(new_n785), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT105), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT105), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n945), .B(new_n961), .C1(new_n785), .C2(new_n958), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n760), .A2(new_n426), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n348), .B1(new_n756), .B2(new_n202), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n964), .B(new_n965), .C1(G143), .C2(new_n749), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n742), .A2(new_n338), .B1(new_n754), .B2(new_n351), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n745), .A2(new_n201), .B1(new_n764), .B2(new_n817), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n966), .B(new_n969), .C1(new_n269), .C2(new_n837), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n754), .A2(new_n469), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n772), .A2(G317), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n971), .B(new_n972), .C1(G303), .C2(new_n743), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n756), .A2(new_n568), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n974), .A2(KEYINPUT46), .B1(new_n831), .B2(new_n750), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(KEYINPUT46), .B2(new_n974), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n261), .B1(new_n745), .B2(new_n834), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(G107), .B2(new_n770), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n973), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n837), .A2(new_n596), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n970), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT47), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n739), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n982), .B2(new_n981), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n237), .A2(new_n791), .ZN(new_n985));
  INV_X1    g0785(.A(new_n381), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n796), .B1(new_n700), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n800), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT106), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n984), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT107), .Z(new_n991));
  INV_X1    g0791(.A(new_n736), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n991), .B1(new_n940), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT108), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n963), .A2(new_n995), .ZN(G387));
  OAI21_X1  g0796(.A(new_n736), .B1(new_n691), .B2(new_n692), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n787), .A2(new_n703), .B1(G107), .B2(new_n210), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n232), .A2(G45), .ZN(new_n999));
  INV_X1    g0799(.A(new_n703), .ZN(new_n1000));
  AOI211_X1 g0800(.A(G45), .B(new_n1000), .C1(G68), .C2(G77), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n251), .A2(G50), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT50), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n792), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n998), .B1(new_n999), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n786), .B1(new_n1005), .B2(new_n796), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n251), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n261), .B(new_n971), .C1(new_n1007), .C2(new_n762), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G68), .A2(new_n746), .B1(new_n772), .B2(G150), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n756), .A2(new_n351), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G50), .B2(new_n743), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n770), .A2(new_n986), .B1(G159), .B2(new_n749), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n348), .B1(new_n774), .B2(G116), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n756), .A2(new_n596), .B1(new_n760), .B2(new_n834), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G317), .A2(new_n743), .B1(new_n746), .B2(G303), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n768), .B2(new_n750), .C1(new_n837), .C2(new_n831), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT48), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n1018), .B2(new_n1017), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT49), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1014), .B1(new_n764), .B2(new_n776), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1013), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1006), .B1(new_n1024), .B2(new_n738), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n954), .A2(new_n785), .B1(new_n997), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n955), .A2(new_n701), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n732), .A2(new_n954), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(G393));
  AOI21_X1  g0829(.A(new_n702), .B1(new_n952), .B2(new_n956), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n956), .B2(new_n952), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n936), .A2(new_n736), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n795), .B1(new_n469), .B2(new_n210), .C1(new_n792), .C2(new_n245), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n786), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n837), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(G50), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n750), .A2(new_n338), .B1(new_n742), .B2(new_n269), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT51), .ZN(new_n1038));
  INV_X1    g0838(.A(G143), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n745), .A2(new_n251), .B1(new_n764), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G68), .B2(new_n757), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n348), .B1(new_n754), .B2(new_n536), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(G77), .B2(new_n770), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1036), .A2(new_n1038), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n745), .A2(new_n596), .B1(new_n764), .B2(new_n768), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(G283), .B2(new_n757), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n348), .B(new_n755), .C1(G116), .C2(new_n770), .ZN(new_n1047));
  INV_X1    g0847(.A(G303), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1046), .B(new_n1047), .C1(new_n837), .C2(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n743), .A2(G311), .B1(G317), .B2(new_n749), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT52), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1044), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT109), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1034), .B1(new_n1053), .B2(new_n738), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n952), .A2(new_n785), .B1(new_n1032), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1031), .A2(new_n1055), .ZN(G390));
  INV_X1    g0856(.A(new_n908), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n630), .A2(new_n516), .A3(new_n684), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n727), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1059), .A2(new_n725), .ZN(new_n1060));
  OAI211_X1 g0860(.A(G330), .B(new_n808), .C1(new_n1058), .C2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n909), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1063), .A2(KEYINPUT113), .B1(new_n729), .B2(new_n847), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n909), .B1(new_n729), .B2(new_n808), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT113), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1057), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT114), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n907), .B(new_n1069), .C1(new_n805), .C2(new_n388), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1061), .B1(new_n909), .B2(new_n1071), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n845), .A2(new_n846), .A3(new_n1070), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1073), .A2(new_n729), .A3(new_n808), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n805), .A2(new_n388), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n695), .B(new_n1076), .C1(new_n709), .C2(new_n664), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT110), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n1077), .A2(new_n1078), .A3(new_n907), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1078), .B1(new_n1077), .B2(new_n907), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(KEYINPUT115), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1077), .A2(new_n907), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT110), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1077), .A2(new_n1078), .A3(new_n907), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT115), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1068), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT116), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n396), .A2(new_n442), .A3(new_n443), .A4(new_n729), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1092), .B(new_n674), .C1(new_n444), .C2(new_n712), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n1090), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n847), .A2(new_n729), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1063), .A2(KEYINPUT113), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n908), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1088), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1093), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT116), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(KEYINPUT117), .B1(new_n1094), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1091), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT117), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1101), .A2(KEYINPUT116), .A3(new_n1102), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT112), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n904), .B1(new_n865), .B2(new_n878), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1084), .A2(new_n909), .A3(new_n1085), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1110), .A2(new_n1111), .A3(KEYINPUT111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT111), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n910), .A2(new_n905), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n899), .B2(new_n902), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1109), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT111), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1110), .A2(new_n1111), .A3(KEYINPUT111), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n903), .A2(new_n1115), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(KEYINPUT112), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1095), .B1(new_n1118), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1095), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n899), .A2(new_n902), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n1128), .A2(new_n1116), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1127), .B1(new_n1129), .B2(new_n1109), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1104), .B(new_n1108), .C1(new_n1126), .C2(new_n1130), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n1114), .A2(new_n1109), .A3(new_n1117), .ZN(new_n1132));
  AOI21_X1  g0932(.A(KEYINPUT112), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1127), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1130), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1131), .A2(new_n701), .A3(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT54), .B(G143), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n261), .B1(new_n746), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(G128), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1141), .B1(new_n269), .B2(new_n760), .C1(new_n750), .C2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n756), .A2(new_n338), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT53), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G132), .A2(new_n743), .B1(new_n772), .B2(G125), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1145), .B(new_n1146), .C1(new_n201), .C2(new_n754), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1143), .B(new_n1147), .C1(G137), .C2(new_n1035), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n348), .B1(new_n757), .B2(G87), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1149), .B1(new_n351), .B2(new_n760), .C1(new_n750), .C2(new_n834), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n837), .A2(new_n372), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n742), .A2(new_n568), .B1(new_n754), .B2(new_n426), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n745), .A2(new_n469), .B1(new_n764), .B2(new_n596), .ZN(new_n1153));
  NOR4_X1   g0953(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n738), .B1(new_n1148), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n814), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1155), .B(new_n786), .C1(new_n1007), .C2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n903), .B2(new_n734), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1118), .A2(new_n1125), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1130), .B1(new_n1159), .B2(new_n1127), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1158), .B1(new_n1160), .B2(new_n785), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1138), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT118), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1138), .A2(KEYINPUT118), .A3(new_n1161), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(G378));
  INV_X1    g0966(.A(KEYINPUT57), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1093), .B1(new_n1160), .B2(new_n1136), .ZN(new_n1168));
  OAI21_X1  g0968(.A(KEYINPUT120), .B1(new_n906), .B2(new_n916), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n367), .A2(new_n370), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n345), .A2(new_n682), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1170), .B(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1172), .B(new_n1173), .Z(new_n1174));
  INV_X1    g0974(.A(KEYINPUT119), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n891), .B2(G330), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n849), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n897), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n880), .B1(new_n901), .B2(new_n865), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n890), .ZN(new_n1180));
  OAI211_X1 g0980(.A(G330), .B(new_n1178), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1181), .A2(KEYINPUT119), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1174), .B1(new_n1176), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1174), .B1(new_n1181), .B2(KEYINPUT119), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1169), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1174), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1181), .A2(KEYINPUT119), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n889), .A2(new_n890), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1189), .A2(new_n1175), .A3(G330), .A4(new_n1178), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1187), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT120), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n914), .A2(new_n915), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1128), .A2(new_n904), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1191), .A2(new_n1195), .A3(new_n1184), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1186), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1167), .B1(new_n1168), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1137), .A2(new_n1102), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT121), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n917), .A2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(KEYINPUT121), .B1(new_n906), .B2(new_n916), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1183), .A2(new_n1201), .A3(new_n1185), .A4(new_n1202), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1200), .B(new_n917), .C1(new_n1191), .C2(new_n1184), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1199), .A2(new_n1205), .A3(KEYINPUT57), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1198), .A2(new_n701), .A3(new_n1206), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n818), .A2(new_n824), .B1(new_n338), .B2(new_n760), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G128), .A2(new_n743), .B1(new_n757), .B2(new_n1140), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n817), .B2(new_n745), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1208), .B(new_n1210), .C1(G125), .C2(new_n749), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n471), .B(new_n291), .C1(new_n754), .C2(new_n269), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G124), .B2(new_n772), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n348), .A2(G41), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1219), .A2(new_n1010), .A3(new_n964), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n469), .B2(new_n818), .C1(new_n568), .C2(new_n750), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n381), .A2(new_n745), .B1(new_n754), .B2(new_n202), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n742), .A2(new_n372), .B1(new_n764), .B2(new_n834), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(KEYINPUT58), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1219), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1224), .A2(KEYINPUT58), .ZN(new_n1227));
  AND4_X1   g1027(.A1(new_n1217), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n786), .B1(G50), .B2(new_n1156), .C1(new_n1228), .C2(new_n739), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1174), .B2(new_n734), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1197), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1230), .B1(new_n1231), .B2(new_n785), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1207), .A2(new_n1232), .ZN(G375));
  INV_X1    g1033(.A(new_n946), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1104), .A2(new_n1234), .A3(new_n1108), .A4(new_n1235), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT122), .Z(new_n1237));
  NAND2_X1  g1037(.A1(new_n1062), .A2(new_n734), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n786), .B1(G68), .B2(new_n1156), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n742), .A2(new_n817), .B1(new_n745), .B2(new_n338), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n348), .B1(new_n754), .B2(new_n202), .C1(new_n750), .C2(new_n824), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n756), .A2(new_n269), .B1(new_n764), .B2(new_n1142), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n760), .A2(new_n201), .ZN(new_n1243));
  OR4_X1    g1043(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n837), .A2(new_n1139), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n261), .B1(new_n754), .B2(new_n351), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT123), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G107), .A2(new_n746), .B1(new_n772), .B2(G303), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G97), .A2(new_n757), .B1(new_n743), .B2(G283), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n770), .A2(new_n986), .B1(G294), .B2(new_n749), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n837), .A2(new_n568), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n1244), .A2(new_n1245), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1253), .A2(KEYINPUT124), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n739), .B1(new_n1253), .B2(KEYINPUT124), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1239), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1101), .A2(new_n785), .B1(new_n1238), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1237), .A2(new_n1257), .ZN(G381));
  OR4_X1    g1058(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1259));
  NOR4_X1   g1059(.A1(G381), .A2(G387), .A3(new_n1162), .A4(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(G375), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(G407));
  INV_X1    g1062(.A(new_n1162), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n680), .A2(G343), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G407), .B(G213), .C1(G375), .C2(new_n1265), .ZN(G409));
  INV_X1    g1066(.A(KEYINPUT127), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(G393), .B(new_n803), .ZN(new_n1268));
  AOI21_X1  g1068(.A(G390), .B1(new_n963), .B2(new_n995), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n963), .A2(new_n995), .A3(G390), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1268), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1271), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1268), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1273), .A2(new_n1269), .A3(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(KEYINPUT126), .B1(new_n1272), .B2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1274), .B1(new_n1273), .B2(new_n1269), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1270), .A2(new_n1268), .A3(new_n1271), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT126), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1276), .A2(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1207), .A2(new_n1164), .A3(new_n1165), .A4(new_n1232), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1231), .A2(new_n1199), .A3(new_n1234), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1230), .B1(new_n1205), .B2(new_n785), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1263), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1282), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1264), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1105), .A2(KEYINPUT60), .A3(new_n1107), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1235), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT60), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1290), .B(new_n701), .C1(new_n1291), .C2(new_n1235), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1257), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n841), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1292), .A2(G384), .A3(new_n1257), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1287), .A2(new_n1288), .A3(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1264), .B1(new_n1282), .B2(new_n1286), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1299), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(new_n1297), .A3(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1300), .A2(new_n1301), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1296), .A2(G2897), .A3(new_n1264), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1296), .B1(G2897), .B2(new_n1264), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT61), .B1(new_n1306), .B2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1281), .B1(new_n1305), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT63), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1298), .A2(new_n1312), .ZN(new_n1313));
  AOI211_X1 g1113(.A(new_n1264), .B(new_n1296), .C1(new_n1282), .C2(new_n1286), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(KEYINPUT63), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1316));
  AND4_X1   g1116(.A1(new_n1313), .A2(new_n1310), .A3(new_n1315), .A4(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1267), .B1(new_n1311), .B2(new_n1317), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1310), .A2(new_n1315), .A3(new_n1313), .A4(new_n1316), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT61), .ZN(new_n1320));
  OR2_X1    g1120(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1320), .B1(new_n1321), .B2(new_n1302), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1301), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1323), .B1(new_n1314), .B2(new_n1303), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1322), .B1(new_n1324), .B2(new_n1300), .ZN(new_n1325));
  OAI211_X1 g1125(.A(KEYINPUT127), .B(new_n1319), .C1(new_n1325), .C2(new_n1281), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1318), .A2(new_n1326), .ZN(G405));
  OAI21_X1  g1127(.A(new_n1282), .B1(new_n1261), .B2(new_n1162), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1328), .B(new_n1296), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(new_n1329), .B(new_n1316), .ZN(G402));
endmodule


