//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT2), .B(G113), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G116), .B(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G116), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n188), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT0), .A2(G128), .ZN(new_n198));
  XNOR2_X1  g012(.A(G143), .B(G146), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(KEYINPUT64), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n198), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n200), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  INV_X1    g025(.A(G134), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(G137), .ZN(new_n213));
  INV_X1    g027(.A(G137), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT11), .A3(G134), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(G137), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G131), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n213), .A2(new_n215), .A3(new_n219), .A4(new_n216), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(KEYINPUT66), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n217), .A2(new_n222), .A3(G131), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n221), .A2(KEYINPUT67), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT67), .B1(new_n221), .B2(new_n223), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n210), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n205), .A2(new_n227), .A3(G128), .ZN(new_n228));
  INV_X1    g042(.A(new_n216), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n212), .A2(G137), .ZN(new_n230));
  OAI21_X1  g044(.A(G131), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n202), .B(new_n204), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n228), .A2(new_n231), .A3(new_n220), .A4(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n226), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n197), .B1(new_n235), .B2(KEYINPUT69), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n226), .A2(new_n237), .A3(new_n234), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT28), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT28), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n235), .A2(new_n197), .ZN(new_n241));
  INV_X1    g055(.A(new_n197), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n226), .A2(new_n242), .A3(new_n234), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n240), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G237), .ZN(new_n245));
  INV_X1    g059(.A(G953), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(G210), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(KEYINPUT27), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G101), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n248), .B(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT29), .ZN(new_n251));
  NOR3_X1   g065(.A1(new_n239), .A2(new_n244), .A3(new_n251), .ZN(new_n252));
  XOR2_X1   g066(.A(KEYINPUT72), .B(G902), .Z(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n187), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n210), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n221), .A2(new_n223), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n221), .A2(KEYINPUT67), .A3(new_n223), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n234), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT69), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(new_n242), .A3(new_n238), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n240), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n241), .A2(new_n243), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n265), .B1(new_n267), .B2(new_n240), .ZN(new_n268));
  OAI211_X1 g082(.A(KEYINPUT73), .B(new_n253), .C1(new_n268), .C2(new_n251), .ZN(new_n269));
  INV_X1    g083(.A(new_n250), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n200), .A2(new_n209), .A3(KEYINPUT65), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT65), .B1(new_n200), .B2(new_n209), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n221), .A2(new_n223), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n234), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n197), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n240), .B1(new_n277), .B2(new_n243), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n270), .B1(new_n265), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT30), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n242), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT68), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n262), .A2(new_n281), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n226), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n283), .B1(new_n226), .B2(new_n284), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n287), .A2(new_n243), .A3(new_n270), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n280), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n255), .B(new_n269), .C1(new_n289), .C2(KEYINPUT29), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G472), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT32), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n262), .B1(new_n273), .B2(new_n274), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n197), .B1(new_n294), .B2(KEYINPUT30), .ZN(new_n295));
  INV_X1    g109(.A(new_n284), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT68), .B1(new_n261), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n226), .A2(new_n283), .A3(new_n284), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n295), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n243), .A2(new_n250), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT31), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT31), .ZN(new_n302));
  INV_X1    g116(.A(new_n300), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n287), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n250), .B1(new_n265), .B2(new_n279), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n293), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n270), .B1(new_n239), .B2(new_n278), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n308), .A2(KEYINPUT70), .A3(new_n301), .A4(new_n304), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(G472), .A2(G902), .ZN(new_n311));
  XOR2_X1   g125(.A(new_n311), .B(KEYINPUT71), .Z(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n292), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  AOI211_X1 g128(.A(KEYINPUT32), .B(new_n312), .C1(new_n307), .C2(new_n309), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n291), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G217), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n317), .B1(new_n253), .B2(G234), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT74), .B1(new_n232), .B2(G119), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n194), .A3(G128), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n232), .A2(G119), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT75), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n320), .A2(new_n322), .A3(new_n326), .A4(new_n323), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT24), .B(G110), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n325), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT23), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n323), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n232), .A2(KEYINPUT23), .A3(G119), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n332), .B(new_n333), .C1(G119), .C2(new_n232), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G110), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT16), .ZN(new_n337));
  INV_X1    g151(.A(G140), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(G125), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(G125), .ZN(new_n340));
  INV_X1    g154(.A(G125), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G140), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n336), .B(new_n339), .C1(new_n343), .C2(new_n337), .ZN(new_n344));
  XNOR2_X1  g158(.A(G125), .B(G140), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(KEYINPUT76), .A3(KEYINPUT16), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n201), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n201), .A3(new_n346), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n330), .B(new_n335), .C1(new_n347), .C2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n347), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT77), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n343), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n345), .A2(KEYINPUT77), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n201), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n329), .B1(new_n325), .B2(new_n327), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n334), .A2(G110), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n351), .B(new_n355), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(KEYINPUT78), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n353), .A2(new_n354), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n347), .B1(new_n201), .B2(new_n361), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n356), .A2(new_n357), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n350), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT22), .B(G137), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n246), .A2(G221), .A3(G234), .ZN(new_n367));
  XOR2_X1   g181(.A(new_n366), .B(new_n367), .Z(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n358), .A2(KEYINPUT78), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n362), .A2(new_n363), .A3(new_n360), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n350), .A3(new_n368), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n370), .A2(new_n253), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT25), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n370), .A2(KEYINPUT25), .A3(new_n253), .A4(new_n374), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n319), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n370), .A2(new_n374), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G902), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n319), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(KEYINPUT79), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n379), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT9), .B(G234), .ZN(new_n388));
  OAI21_X1  g202(.A(G221), .B1(new_n388), .B2(G902), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G469), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(new_n382), .ZN(new_n392));
  INV_X1    g206(.A(G104), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT3), .B1(new_n393), .B2(G107), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT3), .ZN(new_n395));
  INV_X1    g209(.A(G107), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n396), .A3(G104), .ZN(new_n397));
  INV_X1    g211(.A(G101), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n393), .A2(G107), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n394), .A2(new_n397), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n393), .A2(G107), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n396), .A2(G104), .ZN(new_n402));
  OAI21_X1  g216(.A(G101), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n228), .A2(new_n233), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n228), .A2(new_n233), .A3(new_n400), .A4(new_n403), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT12), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n257), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n259), .A2(new_n260), .B1(new_n408), .B2(new_n407), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(KEYINPUT12), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n408), .B(KEYINPUT10), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n394), .A2(new_n397), .A3(new_n399), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G101), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(KEYINPUT4), .A3(new_n400), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT4), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n419), .A3(G101), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n210), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n415), .A2(new_n260), .A3(new_n259), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n414), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G140), .ZN(new_n424));
  INV_X1    g238(.A(G227), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(G953), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n424), .B(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n415), .A2(new_n421), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n259), .A2(new_n260), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n423), .A2(new_n427), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n392), .B1(new_n434), .B2(G469), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n430), .A2(new_n414), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n428), .B1(new_n433), .B2(new_n422), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n391), .B(new_n253), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n390), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G952), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n440), .A2(KEYINPUT93), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n440), .A2(KEYINPUT93), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n246), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(G234), .B2(G237), .ZN(new_n444));
  AOI211_X1 g258(.A(new_n246), .B(new_n253), .C1(G234), .C2(G237), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(G898), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(KEYINPUT94), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n444), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G214), .B1(G237), .B2(G902), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n451), .B(KEYINPUT80), .Z(new_n452));
  OAI21_X1  g266(.A(G210), .B1(G237), .B2(G902), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n190), .A2(KEYINPUT5), .ZN(new_n455));
  INV_X1    g269(.A(G113), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT5), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n456), .B1(new_n193), .B2(new_n457), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n455), .A2(new_n458), .B1(new_n189), .B2(new_n190), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n404), .ZN(new_n460));
  INV_X1    g274(.A(new_n418), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n197), .A2(new_n420), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G110), .B(G122), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT81), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n464), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n466), .A2(new_n467), .A3(KEYINPUT6), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n406), .A2(new_n341), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n470), .B1(new_n210), .B2(new_n341), .ZN(new_n471));
  INV_X1    g285(.A(G224), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(G953), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n471), .B(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n467), .A2(KEYINPUT6), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n463), .A2(new_n465), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n469), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n405), .A2(new_n459), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n464), .B(KEYINPUT8), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n455), .A2(KEYINPUT82), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n194), .A2(G116), .ZN(new_n483));
  OAI21_X1  g297(.A(G113), .B1(new_n483), .B2(KEYINPUT5), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT83), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n458), .A2(KEYINPUT83), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT82), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n190), .A2(new_n488), .A3(KEYINPUT5), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n482), .A2(new_n486), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n191), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT84), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n490), .A2(KEYINPUT84), .A3(new_n191), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n481), .B1(new_n495), .B2(new_n404), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT7), .B1(new_n472), .B2(G953), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n471), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n471), .A2(new_n497), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n468), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n382), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n454), .B1(new_n478), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n501), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n453), .A3(new_n477), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n452), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n439), .A2(new_n450), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT89), .B1(new_n349), .B2(new_n347), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT89), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n351), .A2(new_n508), .A3(new_n348), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n245), .A2(new_n246), .A3(G214), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT85), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(G143), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n203), .A2(KEYINPUT85), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n510), .B1(new_n514), .B2(new_n512), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G131), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n513), .A2(new_n515), .A3(new_n219), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n517), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT17), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n507), .A2(new_n509), .A3(new_n520), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(KEYINPUT18), .A2(G131), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n513), .A2(new_n515), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(KEYINPUT87), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n521), .A2(KEYINPUT18), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT86), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n343), .A2(G146), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n355), .B2(new_n529), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n355), .A2(new_n528), .A3(new_n529), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n526), .B(new_n527), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(G113), .B(G122), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(new_n393), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n523), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n534), .B1(new_n523), .B2(new_n532), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n382), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(G475), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT20), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n347), .B1(new_n519), .B2(new_n517), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT19), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n361), .A2(new_n541), .ZN(new_n542));
  OR3_X1    g356(.A1(new_n345), .A2(KEYINPUT88), .A3(new_n541), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT88), .B1(new_n345), .B2(new_n541), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n540), .B1(new_n545), .B2(G146), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n532), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n534), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n523), .A2(new_n532), .A3(new_n534), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(G475), .A2(G902), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n539), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n552), .ZN(new_n554));
  AOI211_X1 g368(.A(KEYINPUT20), .B(new_n554), .C1(new_n549), .C2(new_n550), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n538), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n388), .A2(new_n317), .A3(G953), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n232), .A2(G143), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n203), .A2(G128), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT13), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT13), .B1(new_n203), .B2(G128), .ZN(new_n562));
  OAI21_X1  g376(.A(G134), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT90), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n559), .A2(new_n558), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n212), .ZN(new_n566));
  INV_X1    g380(.A(G122), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G116), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n192), .A2(G122), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(new_n396), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n396), .B1(new_n568), .B2(new_n569), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n566), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n569), .A2(KEYINPUT14), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n192), .A2(G122), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n569), .B1(new_n575), .B2(KEYINPUT14), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n574), .B1(new_n576), .B2(KEYINPUT91), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(KEYINPUT91), .B2(new_n576), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n578), .A2(G107), .ZN(new_n579));
  INV_X1    g393(.A(new_n566), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n565), .A2(new_n212), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n570), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI221_X1 g396(.A(new_n557), .B1(new_n564), .B2(new_n573), .C1(new_n579), .C2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n557), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n564), .A2(new_n573), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n582), .B1(new_n578), .B2(G107), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n583), .A2(new_n587), .A3(KEYINPUT92), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT92), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n589), .B(new_n584), .C1(new_n585), .C2(new_n586), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n588), .A2(new_n253), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G478), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(KEYINPUT15), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n591), .B(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n556), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n506), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n316), .A2(new_n387), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT95), .B(G101), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G3));
  INV_X1    g414(.A(G472), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(new_n310), .B2(new_n253), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n312), .B1(new_n307), .B2(new_n309), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n505), .A2(new_n450), .ZN(new_n605));
  INV_X1    g419(.A(new_n556), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n588), .A2(new_n607), .A3(new_n590), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n583), .A2(new_n587), .A3(KEYINPUT33), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n608), .A2(G478), .A3(new_n253), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n591), .A2(new_n592), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n605), .A2(new_n606), .A3(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n604), .A2(new_n387), .A3(new_n439), .A4(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT34), .B(G104), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  NAND2_X1  g431(.A1(new_n606), .A2(new_n594), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n605), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n604), .A2(new_n387), .A3(new_n439), .A4(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT35), .B(G107), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  NOR2_X1   g438(.A1(new_n369), .A2(KEYINPUT36), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n365), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n373), .A2(new_n350), .A3(new_n625), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n384), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT98), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n379), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n506), .A2(new_n596), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n604), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT37), .B(G110), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G12));
  XOR2_X1   g449(.A(KEYINPUT99), .B(G900), .Z(new_n636));
  NAND2_X1  g450(.A1(new_n445), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n444), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n618), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n435), .A2(new_n438), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n389), .ZN(new_n643));
  INV_X1    g457(.A(new_n505), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n631), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n316), .A2(new_n641), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G128), .ZN(G30));
  XNOR2_X1  g461(.A(new_n639), .B(KEYINPUT39), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n439), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT40), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n502), .A2(new_n504), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n652), .B(KEYINPUT38), .Z(new_n653));
  NOR2_X1   g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n649), .A2(new_n650), .ZN(new_n655));
  INV_X1    g469(.A(new_n452), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n631), .A2(new_n594), .A3(new_n556), .A4(new_n656), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n657), .A2(KEYINPUT101), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(KEYINPUT101), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n654), .B(new_n655), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(G902), .B1(new_n267), .B2(new_n270), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n270), .B1(new_n287), .B2(new_n243), .ZN(new_n663));
  OAI21_X1  g477(.A(G472), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n664), .B1(new_n314), .B2(new_n315), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT100), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n665), .A2(KEYINPUT100), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n660), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(new_n203), .ZN(G45));
  NAND3_X1  g483(.A1(new_n556), .A2(new_n612), .A3(new_n639), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n316), .A2(new_n645), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  AOI21_X1  g487(.A(new_n437), .B1(new_n414), .B2(new_n430), .ZN(new_n674));
  OAI21_X1  g488(.A(G469), .B1(new_n674), .B2(new_n254), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(new_n438), .A3(new_n389), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT102), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT102), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n675), .A2(new_n438), .A3(new_n678), .A4(new_n389), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n316), .A2(new_n387), .A3(new_n614), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  NAND4_X1  g497(.A1(new_n316), .A2(new_n387), .A3(new_n619), .A4(new_n680), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT103), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT104), .B(G116), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G18));
  NOR2_X1   g502(.A1(new_n644), .A2(new_n676), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n629), .B(KEYINPUT98), .Z(new_n690));
  NAND2_X1  g504(.A1(new_n377), .A2(new_n378), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n318), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  AND4_X1   g507(.A1(new_n595), .A2(new_n689), .A3(new_n693), .A4(new_n450), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n316), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT105), .B(G119), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G21));
  INV_X1    g511(.A(new_n305), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n268), .A2(new_n270), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n312), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n310), .A2(new_n253), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n700), .B1(new_n701), .B2(G472), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n387), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g518(.A(KEYINPUT106), .B1(new_n379), .B2(new_n386), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n505), .A2(new_n594), .A3(new_n556), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT107), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n505), .A2(new_n709), .A3(new_n556), .A4(new_n594), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n677), .A2(new_n450), .A3(new_n679), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n702), .A2(new_n706), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G122), .ZN(G24));
  INV_X1    g528(.A(new_n700), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n254), .B1(new_n307), .B2(new_n309), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n693), .B(new_n715), .C1(new_n716), .C2(new_n601), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n671), .A3(new_n689), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  NAND3_X1  g534(.A1(new_n502), .A2(new_n504), .A3(new_n656), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n643), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n671), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n316), .A2(new_n706), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT42), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n670), .A2(KEYINPUT42), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n316), .A2(new_n727), .A3(new_n387), .A4(new_n722), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n219), .ZN(G33));
  NAND4_X1  g544(.A1(new_n316), .A2(new_n387), .A3(new_n641), .A4(new_n722), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G134), .ZN(G36));
  INV_X1    g546(.A(new_n434), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n391), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n434), .A2(KEYINPUT45), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n392), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n737), .A2(KEYINPUT46), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n438), .B1(new_n737), .B2(KEYINPUT46), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n389), .B(new_n648), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  XOR2_X1   g554(.A(new_n740), .B(KEYINPUT108), .Z(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n556), .A2(KEYINPUT109), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n538), .B(new_n745), .C1(new_n553), .C2(new_n555), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n744), .A2(KEYINPUT43), .A3(new_n612), .A4(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT110), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n749), .B1(new_n613), .B2(new_n556), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n747), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n693), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n748), .B1(new_n747), .B2(new_n750), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n755));
  INV_X1    g569(.A(new_n604), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n754), .A2(new_n755), .A3(KEYINPUT44), .A4(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n747), .A2(new_n750), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT110), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n693), .A3(new_n751), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n758), .B1(new_n761), .B2(new_n604), .ZN(new_n762));
  INV_X1    g576(.A(new_n721), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n757), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n761), .A2(new_n604), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n755), .B1(new_n765), .B2(KEYINPUT44), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n743), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n754), .A2(new_n756), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT111), .B1(new_n768), .B2(new_n758), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n721), .B1(new_n768), .B2(new_n758), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n769), .A2(new_n770), .A3(KEYINPUT112), .A4(new_n757), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n742), .B1(new_n767), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT113), .B(G137), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(G39));
  OR2_X1    g588(.A1(new_n738), .A2(new_n739), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n389), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT47), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(KEYINPUT47), .A3(new_n389), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n316), .ZN(new_n781));
  INV_X1    g595(.A(new_n387), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n781), .A2(new_n782), .A3(new_n671), .A4(new_n763), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  NAND2_X1  g600(.A1(new_n667), .A2(new_n666), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n676), .A2(new_n638), .A3(new_n721), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n787), .A2(new_n782), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(new_n556), .A3(new_n612), .ZN(new_n791));
  INV_X1    g605(.A(new_n706), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n781), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n789), .B1(new_n750), .B2(new_n747), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(KEYINPUT120), .B(KEYINPUT48), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  AND4_X1   g612(.A1(new_n444), .A2(new_n702), .A3(new_n706), .A4(new_n759), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n443), .B1(new_n799), .B2(new_n689), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n791), .A2(new_n797), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n790), .A2(new_n606), .A3(new_n613), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n794), .A2(new_n718), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n653), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n805), .A2(new_n656), .A3(new_n676), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n799), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT50), .Z(new_n808));
  NAND3_X1  g622(.A1(new_n675), .A2(new_n438), .A3(new_n390), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n778), .A2(new_n779), .A3(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n799), .A2(new_n763), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n808), .A2(KEYINPUT51), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n809), .B(KEYINPUT119), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n811), .B1(new_n780), .B2(new_n814), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n803), .A2(new_n808), .A3(new_n802), .A4(new_n815), .ZN(new_n816));
  OAI221_X1 g630(.A(new_n801), .B1(new_n804), .B2(new_n813), .C1(new_n816), .C2(KEYINPUT51), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n690), .A2(new_n692), .A3(new_n439), .A4(new_n639), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n710), .B2(new_n708), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n665), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n820), .B1(new_n665), .B2(new_n822), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n646), .A2(new_n672), .A3(new_n719), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n819), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n646), .A2(new_n672), .A3(new_n719), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n665), .A2(new_n822), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT118), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n665), .A2(new_n820), .A3(new_n822), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n828), .A2(new_n832), .A3(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n827), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT53), .B1(new_n834), .B2(KEYINPUT117), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n827), .A2(new_n833), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n631), .A2(new_n643), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n595), .A2(new_n639), .A3(new_n763), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n316), .A2(new_n837), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n718), .B2(new_n724), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n717), .A2(new_n723), .A3(KEYINPUT116), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n731), .B(new_n842), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n729), .A2(new_n846), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n606), .A2(new_n613), .A3(KEYINPUT114), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT114), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(new_n556), .B2(new_n612), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n848), .A2(new_n506), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n604), .A2(new_n851), .A3(new_n387), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n695), .A2(new_n852), .A3(new_n713), .A4(new_n633), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n598), .A2(new_n620), .ZN(new_n854));
  INV_X1    g668(.A(new_n681), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n684), .B(KEYINPUT103), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n847), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n835), .B1(new_n836), .B2(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n847), .A2(new_n856), .A3(new_n857), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n860), .B(new_n834), .C1(KEYINPUT117), .C2(KEYINPUT53), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n818), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT53), .B1(new_n836), .B2(new_n858), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n598), .A2(new_n620), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n852), .A2(new_n713), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n316), .A2(new_n694), .B1(new_n604), .B2(new_n632), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n864), .A2(new_n681), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n686), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n834), .A2(new_n868), .A3(new_n869), .A4(new_n847), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT54), .B1(new_n863), .B2(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n817), .A2(new_n862), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(G952), .A2(G953), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n675), .A2(new_n438), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n874), .A2(KEYINPUT49), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(KEYINPUT49), .ZN(new_n876));
  AND4_X1   g690(.A1(new_n744), .A2(new_n875), .A3(new_n746), .A4(new_n876), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n613), .A2(new_n452), .A3(new_n390), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n877), .A2(new_n653), .A3(new_n706), .A4(new_n878), .ZN(new_n879));
  OAI22_X1  g693(.A1(new_n872), .A2(new_n873), .B1(new_n787), .B2(new_n879), .ZN(G75));
  AOI21_X1  g694(.A(new_n869), .B1(new_n860), .B2(new_n834), .ZN(new_n881));
  AND4_X1   g695(.A1(new_n869), .A2(new_n834), .A3(new_n868), .A4(new_n847), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n881), .A2(new_n882), .A3(new_n253), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n454), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT56), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n469), .A2(new_n476), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n474), .ZN(new_n887));
  XOR2_X1   g701(.A(KEYINPUT121), .B(KEYINPUT55), .Z(new_n888));
  XNOR2_X1  g702(.A(new_n887), .B(new_n888), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n884), .A2(new_n885), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n889), .B1(new_n884), .B2(new_n885), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n246), .A2(G952), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(G51));
  OAI21_X1  g707(.A(new_n818), .B1(new_n881), .B2(new_n882), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n863), .A2(KEYINPUT54), .A3(new_n870), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(KEYINPUT122), .B(new_n818), .C1(new_n881), .C2(new_n882), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n392), .B(KEYINPUT57), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n674), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n883), .A2(new_n736), .A3(new_n735), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n892), .B1(new_n902), .B2(new_n903), .ZN(G54));
  NAND3_X1  g718(.A1(new_n883), .A2(KEYINPUT58), .A3(G475), .ZN(new_n905));
  INV_X1    g719(.A(new_n551), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n907), .A2(new_n908), .A3(new_n892), .ZN(G60));
  NAND2_X1  g723(.A1(new_n608), .A2(new_n609), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n862), .A2(new_n871), .ZN(new_n911));
  NAND2_X1  g725(.A1(G478), .A2(G902), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT59), .Z(new_n913));
  OAI21_X1  g727(.A(new_n910), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n892), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n910), .A2(new_n913), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n897), .A2(new_n898), .A3(new_n916), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(G63));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n919));
  NAND2_X1  g733(.A1(G217), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT60), .Z(new_n921));
  NAND3_X1  g735(.A1(new_n863), .A2(new_n870), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n863), .A2(KEYINPUT123), .A3(new_n870), .A4(new_n921), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n380), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n915), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n627), .A2(new_n628), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n924), .B2(new_n925), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n919), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n924), .A2(new_n925), .ZN(new_n931));
  INV_X1    g745(.A(new_n928), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n933), .A2(KEYINPUT61), .A3(new_n915), .A4(new_n926), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n930), .A2(new_n934), .ZN(G66));
  OAI21_X1  g749(.A(G953), .B1(new_n448), .B2(new_n472), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n868), .B2(G953), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n886), .B1(G898), .B2(new_n246), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G69));
  INV_X1    g753(.A(G900), .ZN(new_n940));
  OAI21_X1  g754(.A(G953), .B1(new_n425), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT124), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n767), .A2(new_n771), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n741), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n948));
  INV_X1    g762(.A(new_n787), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n948), .B(new_n828), .C1(new_n949), .C2(new_n660), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT62), .B1(new_n668), .B2(new_n826), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n781), .A2(new_n782), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n649), .A2(new_n763), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n848), .A2(new_n850), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n953), .B1(new_n954), .B2(new_n618), .ZN(new_n955));
  AOI22_X1  g769(.A1(new_n780), .A2(new_n784), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n950), .A2(new_n951), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(G953), .B1(new_n947), .B2(new_n957), .ZN(new_n958));
  OAI22_X1  g772(.A1(new_n285), .A2(new_n286), .B1(KEYINPUT30), .B2(new_n294), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(new_n545), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n945), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n960), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n741), .A2(new_n711), .A3(new_n793), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n729), .A2(new_n826), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n963), .A2(new_n731), .A3(new_n964), .A4(new_n785), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n246), .B1(new_n772), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n940), .A2(G953), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n962), .B1(new_n968), .B2(KEYINPUT125), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT125), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n966), .A2(new_n970), .A3(new_n967), .ZN(new_n971));
  AOI211_X1 g785(.A(new_n944), .B(new_n961), .C1(new_n969), .C2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n944), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n968), .A2(KEYINPUT125), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(new_n971), .A3(new_n960), .ZN(new_n975));
  INV_X1    g789(.A(new_n961), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n972), .A2(new_n977), .ZN(G72));
  INV_X1    g792(.A(new_n663), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n947), .A2(new_n868), .A3(new_n957), .ZN(new_n980));
  NAND2_X1  g794(.A1(G472), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT63), .Z(new_n982));
  AOI21_X1  g796(.A(new_n979), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n982), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n772), .A2(new_n965), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(new_n868), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n288), .B(KEYINPUT127), .Z(new_n987));
  OAI21_X1  g801(.A(new_n915), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n859), .A2(new_n861), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n288), .A2(new_n663), .A3(new_n984), .ZN(new_n990));
  AOI211_X1 g804(.A(new_n983), .B(new_n988), .C1(new_n989), .C2(new_n990), .ZN(G57));
endmodule


