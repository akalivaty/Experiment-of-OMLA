

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577;

  XNOR2_X1 U320 ( .A(n324), .B(n323), .ZN(n545) );
  XNOR2_X1 U321 ( .A(n353), .B(n352), .ZN(n563) );
  AND2_X1 U322 ( .A1(G229GAT), .A2(G233GAT), .ZN(n288) );
  XOR2_X1 U323 ( .A(G92GAT), .B(G85GAT), .Z(n289) );
  NOR2_X1 U324 ( .A1(n570), .A2(n359), .ZN(n360) );
  XNOR2_X1 U325 ( .A(n315), .B(n375), .ZN(n320) );
  XNOR2_X1 U326 ( .A(n421), .B(n288), .ZN(n343) );
  XNOR2_X1 U327 ( .A(n320), .B(n319), .ZN(n322) );
  XNOR2_X1 U328 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n427) );
  XNOR2_X1 U329 ( .A(n428), .B(n427), .ZN(n446) );
  NOR2_X1 U330 ( .A1(n446), .A2(n455), .ZN(n553) );
  XNOR2_X1 U331 ( .A(n325), .B(n545), .ZN(n552) );
  XNOR2_X1 U332 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U333 ( .A(n450), .B(n449), .ZN(G1349GAT) );
  XOR2_X1 U334 ( .A(G15GAT), .B(G1GAT), .Z(n349) );
  XOR2_X1 U335 ( .A(G78GAT), .B(G155GAT), .Z(n291) );
  XNOR2_X1 U336 ( .A(G22GAT), .B(G211GAT), .ZN(n290) );
  XNOR2_X1 U337 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U338 ( .A(n349), .B(n292), .Z(n294) );
  NAND2_X1 U339 ( .A1(G231GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U341 ( .A(n295), .B(KEYINPUT78), .Z(n299) );
  XOR2_X1 U342 ( .A(KEYINPUT66), .B(KEYINPUT13), .Z(n297) );
  XNOR2_X1 U343 ( .A(G71GAT), .B(G57GAT), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n338) );
  XNOR2_X1 U345 ( .A(n338), .B(KEYINPUT77), .ZN(n298) );
  XNOR2_X1 U346 ( .A(n299), .B(n298), .ZN(n307) );
  XOR2_X1 U347 ( .A(G64GAT), .B(G183GAT), .Z(n301) );
  XNOR2_X1 U348 ( .A(G8GAT), .B(G127GAT), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U350 ( .A(KEYINPUT14), .B(KEYINPUT76), .Z(n303) );
  XNOR2_X1 U351 ( .A(KEYINPUT15), .B(KEYINPUT12), .ZN(n302) );
  XNOR2_X1 U352 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U353 ( .A(n305), .B(n304), .Z(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n570) );
  INV_X1 U355 ( .A(n570), .ZN(n479) );
  INV_X1 U356 ( .A(KEYINPUT75), .ZN(n325) );
  XOR2_X1 U357 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n309) );
  XNOR2_X1 U358 ( .A(KEYINPUT9), .B(KEYINPUT70), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n324) );
  XOR2_X1 U360 ( .A(KEYINPUT71), .B(KEYINPUT74), .Z(n311) );
  NAND2_X1 U361 ( .A1(G232GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n312), .B(KEYINPUT69), .ZN(n315) );
  XOR2_X1 U364 ( .A(KEYINPUT73), .B(G218GAT), .Z(n314) );
  XNOR2_X1 U365 ( .A(G36GAT), .B(G190GAT), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n375) );
  XOR2_X1 U367 ( .A(G29GAT), .B(G43GAT), .Z(n317) );
  XNOR2_X1 U368 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n317), .B(n316), .ZN(n344) );
  XNOR2_X1 U370 ( .A(G99GAT), .B(G106GAT), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n289), .B(n318), .ZN(n334) );
  XNOR2_X1 U372 ( .A(n344), .B(n334), .ZN(n319) );
  XOR2_X1 U373 ( .A(G50GAT), .B(G162GAT), .Z(n420) );
  XOR2_X1 U374 ( .A(G134GAT), .B(KEYINPUT72), .Z(n401) );
  XNOR2_X1 U375 ( .A(n420), .B(n401), .ZN(n321) );
  XNOR2_X1 U376 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U377 ( .A(n552), .B(KEYINPUT102), .Z(n326) );
  XNOR2_X1 U378 ( .A(n326), .B(KEYINPUT36), .ZN(n575) );
  NOR2_X1 U379 ( .A1(n479), .A2(n575), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n327), .B(KEYINPUT45), .ZN(n355) );
  XOR2_X1 U381 ( .A(G176GAT), .B(G64GAT), .Z(n371) );
  XOR2_X1 U382 ( .A(KEYINPUT67), .B(KEYINPUT33), .Z(n329) );
  XNOR2_X1 U383 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n371), .B(n330), .ZN(n332) );
  AND2_X1 U386 ( .A1(G230GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n333), .B(KEYINPUT32), .ZN(n336) );
  XOR2_X1 U389 ( .A(n334), .B(KEYINPUT68), .Z(n335) );
  XNOR2_X1 U390 ( .A(n336), .B(n335), .ZN(n340) );
  XNOR2_X1 U391 ( .A(G78GAT), .B(G204GAT), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n337), .B(G148GAT), .ZN(n418) );
  XNOR2_X1 U393 ( .A(n418), .B(n338), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n340), .B(n339), .ZN(n566) );
  XOR2_X1 U395 ( .A(G113GAT), .B(G197GAT), .Z(n342) );
  XNOR2_X1 U396 ( .A(G50GAT), .B(G36GAT), .ZN(n341) );
  XNOR2_X1 U397 ( .A(n342), .B(n341), .ZN(n353) );
  XOR2_X1 U398 ( .A(G141GAT), .B(G22GAT), .Z(n421) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U400 ( .A(KEYINPUT65), .B(KEYINPUT30), .Z(n346) );
  XNOR2_X1 U401 ( .A(KEYINPUT64), .B(KEYINPUT29), .ZN(n345) );
  XNOR2_X1 U402 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U403 ( .A(n348), .B(n347), .Z(n351) );
  XOR2_X1 U404 ( .A(G169GAT), .B(G8GAT), .Z(n379) );
  XNOR2_X1 U405 ( .A(n379), .B(n349), .ZN(n350) );
  XNOR2_X1 U406 ( .A(n351), .B(n350), .ZN(n352) );
  INV_X1 U407 ( .A(n563), .ZN(n493) );
  AND2_X1 U408 ( .A1(n566), .A2(n493), .ZN(n354) );
  AND2_X1 U409 ( .A1(n355), .A2(n354), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n356), .B(KEYINPUT116), .ZN(n364) );
  XNOR2_X1 U411 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n358) );
  XNOR2_X1 U412 ( .A(KEYINPUT41), .B(n566), .ZN(n492) );
  NAND2_X1 U413 ( .A1(n563), .A2(n492), .ZN(n357) );
  XOR2_X1 U414 ( .A(n358), .B(n357), .Z(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(KEYINPUT115), .ZN(n361) );
  NOR2_X1 U416 ( .A1(n545), .A2(n361), .ZN(n362) );
  XOR2_X1 U417 ( .A(KEYINPUT47), .B(n362), .Z(n363) );
  NOR2_X1 U418 ( .A1(n364), .A2(n363), .ZN(n365) );
  XNOR2_X1 U419 ( .A(n365), .B(KEYINPUT48), .ZN(n536) );
  XOR2_X1 U420 ( .A(KEYINPUT83), .B(KEYINPUT17), .Z(n367) );
  XNOR2_X1 U421 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U423 ( .A(KEYINPUT19), .B(n368), .Z(n441) );
  XOR2_X1 U424 ( .A(G211GAT), .B(KEYINPUT21), .Z(n370) );
  XNOR2_X1 U425 ( .A(G197GAT), .B(KEYINPUT87), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n415) );
  XOR2_X1 U427 ( .A(n371), .B(n415), .Z(n373) );
  NAND2_X1 U428 ( .A1(G226GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U429 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U430 ( .A(n374), .B(KEYINPUT94), .Z(n377) );
  XNOR2_X1 U431 ( .A(n375), .B(KEYINPUT95), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U433 ( .A(n378), .B(G92GAT), .Z(n381) );
  XNOR2_X1 U434 ( .A(n379), .B(G204GAT), .ZN(n380) );
  XNOR2_X1 U435 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U436 ( .A(n441), .B(n382), .ZN(n469) );
  NOR2_X1 U437 ( .A1(n536), .A2(n469), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n383), .B(KEYINPUT54), .ZN(n559) );
  XOR2_X1 U439 ( .A(KEYINPUT89), .B(KEYINPUT93), .Z(n385) );
  XNOR2_X1 U440 ( .A(G148GAT), .B(KEYINPUT5), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U442 ( .A(G85GAT), .B(G162GAT), .Z(n387) );
  XNOR2_X1 U443 ( .A(G29GAT), .B(G141GAT), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n389), .B(n388), .ZN(n408) );
  XOR2_X1 U446 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n391) );
  XNOR2_X1 U447 ( .A(KEYINPUT4), .B(KEYINPUT92), .ZN(n390) );
  XNOR2_X1 U448 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U449 ( .A(G57GAT), .B(KEYINPUT1), .Z(n393) );
  XNOR2_X1 U450 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U452 ( .A(n395), .B(n394), .Z(n406) );
  XOR2_X1 U453 ( .A(KEYINPUT79), .B(G127GAT), .Z(n397) );
  XNOR2_X1 U454 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U456 ( .A(G113GAT), .B(n398), .Z(n445) );
  XOR2_X1 U457 ( .A(G155GAT), .B(KEYINPUT88), .Z(n400) );
  XNOR2_X1 U458 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n400), .B(n399), .ZN(n414) );
  XOR2_X1 U460 ( .A(n401), .B(n414), .Z(n403) );
  NAND2_X1 U461 ( .A1(G225GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n445), .B(n404), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n509) );
  INV_X1 U466 ( .A(n509), .ZN(n560) );
  XOR2_X1 U467 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n410) );
  XNOR2_X1 U468 ( .A(G218GAT), .B(G106GAT), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n410), .B(n409), .ZN(n425) );
  XOR2_X1 U470 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n412) );
  NAND2_X1 U471 ( .A1(G228GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U472 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U473 ( .A(n413), .B(KEYINPUT22), .Z(n417) );
  XNOR2_X1 U474 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n417), .B(n416), .ZN(n419) );
  XOR2_X1 U476 ( .A(n419), .B(n418), .Z(n423) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U479 ( .A(n425), .B(n424), .Z(n457) );
  AND2_X1 U480 ( .A1(n560), .A2(n457), .ZN(n426) );
  NAND2_X1 U481 ( .A1(n559), .A2(n426), .ZN(n428) );
  XOR2_X1 U482 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n430) );
  XNOR2_X1 U483 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U485 ( .A(KEYINPUT82), .B(KEYINPUT84), .Z(n432) );
  XNOR2_X1 U486 ( .A(G71GAT), .B(G176GAT), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U488 ( .A(n434), .B(n433), .Z(n443) );
  XOR2_X1 U489 ( .A(G190GAT), .B(G134GAT), .Z(n436) );
  XNOR2_X1 U490 ( .A(G43GAT), .B(G99GAT), .ZN(n435) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U492 ( .A(G15GAT), .B(n437), .Z(n439) );
  NAND2_X1 U493 ( .A1(G227GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n455) );
  NAND2_X1 U498 ( .A1(n553), .A2(n492), .ZN(n450) );
  XOR2_X1 U499 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n448) );
  XNOR2_X1 U500 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n447) );
  XOR2_X1 U501 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n467) );
  NAND2_X1 U502 ( .A1(n563), .A2(n566), .ZN(n482) );
  NOR2_X1 U503 ( .A1(n479), .A2(n552), .ZN(n451) );
  XNOR2_X1 U504 ( .A(n451), .B(KEYINPUT16), .ZN(n465) );
  XOR2_X1 U505 ( .A(n457), .B(KEYINPUT28), .Z(n518) );
  XOR2_X1 U506 ( .A(KEYINPUT27), .B(n469), .Z(n454) );
  NAND2_X1 U507 ( .A1(n509), .A2(n454), .ZN(n535) );
  NOR2_X1 U508 ( .A1(n518), .A2(n535), .ZN(n523) );
  NAND2_X1 U509 ( .A1(n523), .A2(n455), .ZN(n464) );
  XNOR2_X1 U510 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n453) );
  INV_X1 U511 ( .A(n455), .ZN(n524) );
  NOR2_X1 U512 ( .A1(n524), .A2(n457), .ZN(n452) );
  XNOR2_X1 U513 ( .A(n453), .B(n452), .ZN(n561) );
  NAND2_X1 U514 ( .A1(n454), .A2(n561), .ZN(n461) );
  NOR2_X1 U515 ( .A1(n455), .A2(n469), .ZN(n456) );
  XNOR2_X1 U516 ( .A(KEYINPUT97), .B(n456), .ZN(n458) );
  NAND2_X1 U517 ( .A1(n458), .A2(n457), .ZN(n459) );
  XOR2_X1 U518 ( .A(KEYINPUT25), .B(n459), .Z(n460) );
  NAND2_X1 U519 ( .A1(n461), .A2(n460), .ZN(n462) );
  NAND2_X1 U520 ( .A1(n462), .A2(n560), .ZN(n463) );
  NAND2_X1 U521 ( .A1(n464), .A2(n463), .ZN(n478) );
  NAND2_X1 U522 ( .A1(n465), .A2(n478), .ZN(n494) );
  NOR2_X1 U523 ( .A1(n482), .A2(n494), .ZN(n475) );
  NAND2_X1 U524 ( .A1(n475), .A2(n509), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U526 ( .A(G1GAT), .B(n468), .Z(G1324GAT) );
  INV_X1 U527 ( .A(n469), .ZN(n512) );
  NAND2_X1 U528 ( .A1(n475), .A2(n512), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n470), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U530 ( .A(KEYINPUT35), .B(KEYINPUT100), .Z(n472) );
  NAND2_X1 U531 ( .A1(n475), .A2(n524), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n472), .B(n471), .ZN(n474) );
  XOR2_X1 U533 ( .A(G15GAT), .B(KEYINPUT99), .Z(n473) );
  XNOR2_X1 U534 ( .A(n474), .B(n473), .ZN(G1326GAT) );
  XOR2_X1 U535 ( .A(G22GAT), .B(KEYINPUT101), .Z(n477) );
  NAND2_X1 U536 ( .A1(n475), .A2(n518), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n477), .B(n476), .ZN(G1327GAT) );
  XOR2_X1 U538 ( .A(G29GAT), .B(KEYINPUT39), .Z(n485) );
  NAND2_X1 U539 ( .A1(n479), .A2(n478), .ZN(n480) );
  NOR2_X1 U540 ( .A1(n575), .A2(n480), .ZN(n481) );
  XNOR2_X1 U541 ( .A(KEYINPUT37), .B(n481), .ZN(n506) );
  NOR2_X1 U542 ( .A1(n482), .A2(n506), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n483), .B(KEYINPUT38), .ZN(n489) );
  NAND2_X1 U544 ( .A1(n509), .A2(n489), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n485), .B(n484), .ZN(G1328GAT) );
  NAND2_X1 U546 ( .A1(n512), .A2(n489), .ZN(n486) );
  XNOR2_X1 U547 ( .A(G36GAT), .B(n486), .ZN(G1329GAT) );
  NAND2_X1 U548 ( .A1(n489), .A2(n524), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n487), .B(KEYINPUT40), .ZN(n488) );
  XNOR2_X1 U550 ( .A(G43GAT), .B(n488), .ZN(G1330GAT) );
  XOR2_X1 U551 ( .A(G50GAT), .B(KEYINPUT103), .Z(n491) );
  NAND2_X1 U552 ( .A1(n518), .A2(n489), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(G1331GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n497) );
  NAND2_X1 U555 ( .A1(n493), .A2(n492), .ZN(n507) );
  NOR2_X1 U556 ( .A1(n507), .A2(n494), .ZN(n495) );
  XOR2_X1 U557 ( .A(KEYINPUT105), .B(n495), .Z(n501) );
  NAND2_X1 U558 ( .A1(n501), .A2(n509), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U560 ( .A(G57GAT), .B(n498), .Z(G1332GAT) );
  NAND2_X1 U561 ( .A1(n501), .A2(n512), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n499), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U563 ( .A1(n501), .A2(n524), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n500), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n503) );
  NAND2_X1 U566 ( .A1(n501), .A2(n518), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(n505) );
  XOR2_X1 U568 ( .A(G78GAT), .B(KEYINPUT106), .Z(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(G1335GAT) );
  XOR2_X1 U570 ( .A(G85GAT), .B(KEYINPUT109), .Z(n511) );
  NOR2_X1 U571 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n508), .B(KEYINPUT108), .ZN(n517) );
  NAND2_X1 U573 ( .A1(n509), .A2(n517), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(G1336GAT) );
  NAND2_X1 U575 ( .A1(n517), .A2(n512), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n513), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n515) );
  NAND2_X1 U578 ( .A1(n524), .A2(n517), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U580 ( .A(G99GAT), .B(n516), .ZN(G1338GAT) );
  XNOR2_X1 U581 ( .A(G106GAT), .B(KEYINPUT112), .ZN(n522) );
  XOR2_X1 U582 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n520) );
  NAND2_X1 U583 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n522), .B(n521), .ZN(G1339GAT) );
  NAND2_X1 U586 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U587 ( .A1(n536), .A2(n525), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n563), .A2(n532), .ZN(n526) );
  XNOR2_X1 U589 ( .A(n526), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n528) );
  NAND2_X1 U591 ( .A1(n532), .A2(n492), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U593 ( .A(G120GAT), .B(n529), .Z(G1341GAT) );
  NAND2_X1 U594 ( .A1(n570), .A2(n532), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n530), .B(KEYINPUT50), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G127GAT), .B(n531), .ZN(G1342GAT) );
  XOR2_X1 U597 ( .A(G134GAT), .B(KEYINPUT51), .Z(n534) );
  NAND2_X1 U598 ( .A1(n532), .A2(n552), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(G1343GAT) );
  NOR2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U601 ( .A1(n537), .A2(n561), .ZN(n538) );
  XOR2_X1 U602 ( .A(KEYINPUT118), .B(n538), .Z(n546) );
  NAND2_X1 U603 ( .A1(n546), .A2(n563), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n539), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n541) );
  NAND2_X1 U606 ( .A1(n546), .A2(n492), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(n542), .ZN(G1345GAT) );
  XOR2_X1 U609 ( .A(G155GAT), .B(KEYINPUT119), .Z(n544) );
  NAND2_X1 U610 ( .A1(n546), .A2(n570), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(G1346GAT) );
  NAND2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n547), .B(KEYINPUT120), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G162GAT), .B(n548), .ZN(G1347GAT) );
  NAND2_X1 U615 ( .A1(n563), .A2(n553), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n549), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U617 ( .A(G183GAT), .B(KEYINPUT123), .Z(n551) );
  NAND2_X1 U618 ( .A1(n553), .A2(n570), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(G1350GAT) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT58), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n557) );
  XNOR2_X1 U624 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U626 ( .A(KEYINPUT124), .B(n558), .Z(n565) );
  AND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n574) );
  INV_X1 U629 ( .A(n574), .ZN(n569) );
  NAND2_X1 U630 ( .A1(n569), .A2(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1352GAT) );
  XOR2_X1 U632 ( .A(G204GAT), .B(KEYINPUT61), .Z(n568) );
  OR2_X1 U633 ( .A1(n574), .A2(n566), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1353GAT) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n573) );
  XNOR2_X1 U638 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n577) );
  NOR2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(n577), .B(n576), .Z(G1355GAT) );
endmodule

