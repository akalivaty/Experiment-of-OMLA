

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U552 ( .A1(n719), .A2(n601), .ZN(n662) );
  AND2_X1 U553 ( .A1(n616), .A2(n615), .ZN(n520) );
  AND2_X1 U554 ( .A1(n750), .A2(n741), .ZN(n521) );
  OR2_X1 U555 ( .A1(KEYINPUT33), .A2(n686), .ZN(n522) );
  INV_X1 U556 ( .A(KEYINPUT95), .ZN(n602) );
  XNOR2_X1 U557 ( .A(n603), .B(n602), .ZN(n605) );
  AND2_X1 U558 ( .A1(n520), .A2(n969), .ZN(n629) );
  INV_X1 U559 ( .A(KEYINPUT29), .ZN(n643) );
  XNOR2_X1 U560 ( .A(n644), .B(n643), .ZN(n649) );
  INV_X1 U561 ( .A(KEYINPUT97), .ZN(n678) );
  XNOR2_X1 U562 ( .A(n679), .B(n678), .ZN(n698) );
  INV_X1 U563 ( .A(KEYINPUT64), .ZN(n523) );
  NOR2_X1 U564 ( .A1(G164), .A2(G1384), .ZN(n719) );
  XNOR2_X1 U565 ( .A(n523), .B(KEYINPUT17), .ZN(n524) );
  NAND2_X1 U566 ( .A1(n521), .A2(n742), .ZN(n743) );
  NOR2_X1 U567 ( .A1(G651), .A2(G543), .ZN(n783) );
  XNOR2_X1 U568 ( .A(n525), .B(n524), .ZN(n889) );
  NOR2_X1 U569 ( .A1(G651), .A2(n580), .ZN(n787) );
  NOR2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  NAND2_X1 U571 ( .A1(G138), .A2(n889), .ZN(n528) );
  INV_X1 U572 ( .A(G2105), .ZN(n529) );
  AND2_X1 U573 ( .A1(n529), .A2(G2104), .ZN(n888) );
  NAND2_X1 U574 ( .A1(G102), .A2(n888), .ZN(n526) );
  XOR2_X1 U575 ( .A(KEYINPUT85), .B(n526), .Z(n527) );
  NAND2_X1 U576 ( .A1(n528), .A2(n527), .ZN(n533) );
  NOR2_X1 U577 ( .A1(G2104), .A2(n529), .ZN(n892) );
  NAND2_X1 U578 ( .A1(G126), .A2(n892), .ZN(n531) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n894) );
  NAND2_X1 U580 ( .A1(G114), .A2(n894), .ZN(n530) );
  NAND2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U582 ( .A1(n533), .A2(n532), .ZN(G164) );
  NAND2_X1 U583 ( .A1(n894), .A2(G113), .ZN(n536) );
  NAND2_X1 U584 ( .A1(G101), .A2(n888), .ZN(n534) );
  XOR2_X1 U585 ( .A(KEYINPUT23), .B(n534), .Z(n535) );
  NAND2_X1 U586 ( .A1(n536), .A2(n535), .ZN(n540) );
  NAND2_X1 U587 ( .A1(n892), .A2(G125), .ZN(n538) );
  NAND2_X1 U588 ( .A1(G137), .A2(n889), .ZN(n537) );
  NAND2_X1 U589 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U590 ( .A1(n540), .A2(n539), .ZN(G160) );
  NAND2_X1 U591 ( .A1(G91), .A2(n783), .ZN(n543) );
  XNOR2_X1 U592 ( .A(G543), .B(KEYINPUT0), .ZN(n541) );
  XNOR2_X1 U593 ( .A(n541), .B(KEYINPUT65), .ZN(n580) );
  INV_X1 U594 ( .A(G651), .ZN(n544) );
  NOR2_X1 U595 ( .A1(n580), .A2(n544), .ZN(n784) );
  NAND2_X1 U596 ( .A1(G78), .A2(n784), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n543), .A2(n542), .ZN(n550) );
  NAND2_X1 U598 ( .A1(n787), .A2(G53), .ZN(n548) );
  NOR2_X1 U599 ( .A1(G543), .A2(n544), .ZN(n545) );
  XOR2_X1 U600 ( .A(KEYINPUT1), .B(n545), .Z(n546) );
  XNOR2_X1 U601 ( .A(KEYINPUT66), .B(n546), .ZN(n788) );
  NAND2_X1 U602 ( .A1(G65), .A2(n788), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U604 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U605 ( .A(n551), .B(KEYINPUT71), .ZN(G299) );
  XNOR2_X1 U606 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n557) );
  NAND2_X1 U607 ( .A1(n784), .A2(G77), .ZN(n552) );
  XNOR2_X1 U608 ( .A(n552), .B(KEYINPUT68), .ZN(n554) );
  NAND2_X1 U609 ( .A1(G90), .A2(n783), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U611 ( .A(n555), .B(KEYINPUT9), .ZN(n556) );
  XNOR2_X1 U612 ( .A(n557), .B(n556), .ZN(n561) );
  NAND2_X1 U613 ( .A1(n787), .A2(G52), .ZN(n559) );
  NAND2_X1 U614 ( .A1(G64), .A2(n788), .ZN(n558) );
  NAND2_X1 U615 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U616 ( .A1(n561), .A2(n560), .ZN(G171) );
  INV_X1 U617 ( .A(G171), .ZN(G301) );
  NAND2_X1 U618 ( .A1(n783), .A2(G89), .ZN(n562) );
  XNOR2_X1 U619 ( .A(n562), .B(KEYINPUT4), .ZN(n564) );
  NAND2_X1 U620 ( .A1(G76), .A2(n784), .ZN(n563) );
  NAND2_X1 U621 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U622 ( .A(n565), .B(KEYINPUT5), .ZN(n570) );
  NAND2_X1 U623 ( .A1(n787), .A2(G51), .ZN(n567) );
  NAND2_X1 U624 ( .A1(G63), .A2(n788), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U626 ( .A(KEYINPUT6), .B(n568), .Z(n569) );
  NAND2_X1 U627 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U628 ( .A(n571), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U629 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U630 ( .A1(G88), .A2(n783), .ZN(n573) );
  NAND2_X1 U631 ( .A1(G75), .A2(n784), .ZN(n572) );
  NAND2_X1 U632 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U633 ( .A(KEYINPUT82), .B(n574), .Z(n576) );
  NAND2_X1 U634 ( .A1(G62), .A2(n788), .ZN(n575) );
  NAND2_X1 U635 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U636 ( .A1(G50), .A2(n787), .ZN(n577) );
  XNOR2_X1 U637 ( .A(KEYINPUT81), .B(n577), .ZN(n578) );
  NOR2_X1 U638 ( .A1(n579), .A2(n578), .ZN(G166) );
  XOR2_X1 U639 ( .A(KEYINPUT86), .B(G166), .Z(G303) );
  NAND2_X1 U640 ( .A1(G87), .A2(n580), .ZN(n582) );
  NAND2_X1 U641 ( .A1(G74), .A2(G651), .ZN(n581) );
  NAND2_X1 U642 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U643 ( .A1(n788), .A2(n583), .ZN(n585) );
  NAND2_X1 U644 ( .A1(n787), .A2(G49), .ZN(n584) );
  NAND2_X1 U645 ( .A1(n585), .A2(n584), .ZN(G288) );
  NAND2_X1 U646 ( .A1(G86), .A2(n783), .ZN(n592) );
  NAND2_X1 U647 ( .A1(n787), .A2(G48), .ZN(n587) );
  NAND2_X1 U648 ( .A1(G61), .A2(n788), .ZN(n586) );
  NAND2_X1 U649 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U650 ( .A1(n784), .A2(G73), .ZN(n588) );
  XOR2_X1 U651 ( .A(KEYINPUT2), .B(n588), .Z(n589) );
  NOR2_X1 U652 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U653 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U654 ( .A(n593), .B(KEYINPUT80), .ZN(G305) );
  NAND2_X1 U655 ( .A1(n787), .A2(G47), .ZN(n595) );
  NAND2_X1 U656 ( .A1(G60), .A2(n788), .ZN(n594) );
  NAND2_X1 U657 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U658 ( .A(KEYINPUT67), .B(n596), .ZN(n600) );
  NAND2_X1 U659 ( .A1(G85), .A2(n783), .ZN(n598) );
  NAND2_X1 U660 ( .A1(G72), .A2(n784), .ZN(n597) );
  AND2_X1 U661 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U662 ( .A1(n600), .A2(n599), .ZN(G290) );
  NAND2_X1 U663 ( .A1(G160), .A2(G40), .ZN(n718) );
  INV_X1 U664 ( .A(n718), .ZN(n601) );
  INV_X1 U665 ( .A(n662), .ZN(n645) );
  NAND2_X1 U666 ( .A1(n645), .A2(G2067), .ZN(n603) );
  NAND2_X1 U667 ( .A1(G1348), .A2(n662), .ZN(n604) );
  NAND2_X1 U668 ( .A1(n605), .A2(n604), .ZN(n631) );
  NAND2_X1 U669 ( .A1(G92), .A2(n783), .ZN(n607) );
  NAND2_X1 U670 ( .A1(G79), .A2(n784), .ZN(n606) );
  NAND2_X1 U671 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U672 ( .A1(n787), .A2(G54), .ZN(n609) );
  NAND2_X1 U673 ( .A1(G66), .A2(n788), .ZN(n608) );
  NAND2_X1 U674 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U675 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U676 ( .A(n612), .B(KEYINPUT15), .ZN(n975) );
  NAND2_X1 U677 ( .A1(n631), .A2(n975), .ZN(n630) );
  XNOR2_X1 U678 ( .A(G1996), .B(KEYINPUT93), .ZN(n946) );
  NOR2_X1 U679 ( .A1(n662), .A2(n946), .ZN(n614) );
  XOR2_X1 U680 ( .A(KEYINPUT26), .B(KEYINPUT94), .Z(n613) );
  XNOR2_X1 U681 ( .A(n614), .B(n613), .ZN(n616) );
  NAND2_X1 U682 ( .A1(n662), .A2(G1341), .ZN(n615) );
  NAND2_X1 U683 ( .A1(G56), .A2(n788), .ZN(n617) );
  XNOR2_X1 U684 ( .A(n617), .B(KEYINPUT14), .ZN(n619) );
  NAND2_X1 U685 ( .A1(G43), .A2(n787), .ZN(n618) );
  NAND2_X1 U686 ( .A1(n619), .A2(n618), .ZN(n627) );
  NAND2_X1 U687 ( .A1(G81), .A2(n783), .ZN(n620) );
  XNOR2_X1 U688 ( .A(n620), .B(KEYINPUT72), .ZN(n621) );
  XNOR2_X1 U689 ( .A(n621), .B(KEYINPUT12), .ZN(n623) );
  NAND2_X1 U690 ( .A1(G68), .A2(n784), .ZN(n622) );
  NAND2_X1 U691 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U692 ( .A(KEYINPUT13), .B(n624), .ZN(n625) );
  XNOR2_X1 U693 ( .A(KEYINPUT73), .B(n625), .ZN(n626) );
  NOR2_X1 U694 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X2 U695 ( .A(KEYINPUT74), .B(n628), .ZN(n969) );
  AND2_X1 U696 ( .A1(n630), .A2(n629), .ZN(n633) );
  NOR2_X1 U697 ( .A1(n631), .A2(n975), .ZN(n632) );
  NOR2_X1 U698 ( .A1(n633), .A2(n632), .ZN(n638) );
  NAND2_X1 U699 ( .A1(n645), .A2(G2072), .ZN(n634) );
  XNOR2_X1 U700 ( .A(n634), .B(KEYINPUT27), .ZN(n636) );
  AND2_X1 U701 ( .A1(G1956), .A2(n662), .ZN(n635) );
  NOR2_X1 U702 ( .A1(n636), .A2(n635), .ZN(n639) );
  INV_X1 U703 ( .A(G299), .ZN(n800) );
  NAND2_X1 U704 ( .A1(n639), .A2(n800), .ZN(n637) );
  NAND2_X1 U705 ( .A1(n638), .A2(n637), .ZN(n642) );
  NOR2_X1 U706 ( .A1(n639), .A2(n800), .ZN(n640) );
  XOR2_X1 U707 ( .A(n640), .B(KEYINPUT28), .Z(n641) );
  NAND2_X1 U708 ( .A1(n642), .A2(n641), .ZN(n644) );
  XOR2_X1 U709 ( .A(G2078), .B(KEYINPUT25), .Z(n955) );
  NOR2_X1 U710 ( .A1(n955), .A2(n662), .ZN(n647) );
  NOR2_X1 U711 ( .A1(n645), .A2(G1961), .ZN(n646) );
  NOR2_X1 U712 ( .A1(n647), .A2(n646), .ZN(n656) );
  OR2_X1 U713 ( .A1(n656), .A2(G301), .ZN(n648) );
  NAND2_X1 U714 ( .A1(n649), .A2(n648), .ZN(n661) );
  INV_X1 U715 ( .A(G8), .ZN(n650) );
  NOR2_X1 U716 ( .A1(n650), .A2(G1966), .ZN(n651) );
  AND2_X1 U717 ( .A1(n662), .A2(n651), .ZN(n673) );
  NOR2_X1 U718 ( .A1(G2084), .A2(n662), .ZN(n670) );
  NOR2_X1 U719 ( .A1(n673), .A2(n670), .ZN(n652) );
  NAND2_X1 U720 ( .A1(G8), .A2(n652), .ZN(n653) );
  XNOR2_X1 U721 ( .A(KEYINPUT30), .B(n653), .ZN(n654) );
  NOR2_X1 U722 ( .A1(G168), .A2(n654), .ZN(n655) );
  XOR2_X1 U723 ( .A(KEYINPUT96), .B(n655), .Z(n658) );
  NAND2_X1 U724 ( .A1(n656), .A2(G301), .ZN(n657) );
  NAND2_X1 U725 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U726 ( .A(KEYINPUT31), .B(n659), .ZN(n660) );
  NAND2_X1 U727 ( .A1(n661), .A2(n660), .ZN(n671) );
  NAND2_X1 U728 ( .A1(n671), .A2(G286), .ZN(n668) );
  NAND2_X1 U729 ( .A1(G8), .A2(n662), .ZN(n700) );
  NOR2_X1 U730 ( .A1(G1971), .A2(n700), .ZN(n664) );
  NOR2_X1 U731 ( .A1(G2090), .A2(n662), .ZN(n663) );
  NOR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U733 ( .A1(n665), .A2(G303), .ZN(n666) );
  OR2_X1 U734 ( .A1(n650), .A2(n666), .ZN(n667) );
  AND2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U736 ( .A(n669), .B(KEYINPUT32), .ZN(n677) );
  NAND2_X1 U737 ( .A1(G8), .A2(n670), .ZN(n675) );
  INV_X1 U738 ( .A(n671), .ZN(n672) );
  NOR2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n679) );
  NOR2_X1 U742 ( .A1(G1976), .A2(G288), .ZN(n688) );
  NOR2_X1 U743 ( .A1(G303), .A2(G1971), .ZN(n680) );
  NOR2_X1 U744 ( .A1(n688), .A2(n680), .ZN(n681) );
  NAND2_X1 U745 ( .A1(n698), .A2(n681), .ZN(n682) );
  XNOR2_X1 U746 ( .A(n682), .B(KEYINPUT98), .ZN(n685) );
  NAND2_X1 U747 ( .A1(G1976), .A2(G288), .ZN(n980) );
  INV_X1 U748 ( .A(n980), .ZN(n683) );
  NOR2_X1 U749 ( .A1(n700), .A2(n683), .ZN(n684) );
  AND2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U751 ( .A(G1981), .B(G305), .ZN(n687) );
  XNOR2_X1 U752 ( .A(n687), .B(KEYINPUT100), .ZN(n971) );
  INV_X1 U753 ( .A(n971), .ZN(n693) );
  INV_X1 U754 ( .A(KEYINPUT99), .ZN(n691) );
  INV_X1 U755 ( .A(n688), .ZN(n979) );
  NOR2_X1 U756 ( .A1(n700), .A2(n979), .ZN(n689) );
  NAND2_X1 U757 ( .A1(KEYINPUT33), .A2(n689), .ZN(n690) );
  XNOR2_X1 U758 ( .A(n691), .B(n690), .ZN(n692) );
  AND2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n694) );
  AND2_X1 U760 ( .A1(n522), .A2(n694), .ZN(n707) );
  NOR2_X1 U761 ( .A1(G303), .A2(G2090), .ZN(n695) );
  NAND2_X1 U762 ( .A1(G8), .A2(n695), .ZN(n696) );
  XOR2_X1 U763 ( .A(KEYINPUT101), .B(n696), .Z(n697) );
  NAND2_X1 U764 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U765 ( .A1(n700), .A2(n699), .ZN(n705) );
  INV_X1 U766 ( .A(n700), .ZN(n703) );
  NOR2_X1 U767 ( .A1(G1981), .A2(G305), .ZN(n701) );
  XNOR2_X1 U768 ( .A(n701), .B(KEYINPUT24), .ZN(n702) );
  NAND2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U770 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U771 ( .A1(n707), .A2(n706), .ZN(n744) );
  NAND2_X1 U772 ( .A1(n888), .A2(G104), .ZN(n708) );
  XOR2_X1 U773 ( .A(KEYINPUT87), .B(n708), .Z(n710) );
  NAND2_X1 U774 ( .A1(G140), .A2(n889), .ZN(n709) );
  NAND2_X1 U775 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U776 ( .A(KEYINPUT34), .B(n711), .ZN(n716) );
  NAND2_X1 U777 ( .A1(G128), .A2(n892), .ZN(n713) );
  NAND2_X1 U778 ( .A1(G116), .A2(n894), .ZN(n712) );
  NAND2_X1 U779 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U780 ( .A(KEYINPUT35), .B(n714), .Z(n715) );
  NOR2_X1 U781 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U782 ( .A(KEYINPUT36), .B(n717), .ZN(n901) );
  XNOR2_X1 U783 ( .A(KEYINPUT37), .B(G2067), .ZN(n753) );
  NOR2_X1 U784 ( .A1(n901), .A2(n753), .ZN(n918) );
  NOR2_X1 U785 ( .A1(n719), .A2(n718), .ZN(n755) );
  NAND2_X1 U786 ( .A1(n918), .A2(n755), .ZN(n720) );
  XNOR2_X1 U787 ( .A(n720), .B(KEYINPUT88), .ZN(n750) );
  NAND2_X1 U788 ( .A1(G105), .A2(n888), .ZN(n721) );
  XNOR2_X1 U789 ( .A(n721), .B(KEYINPUT38), .ZN(n729) );
  NAND2_X1 U790 ( .A1(G117), .A2(n894), .ZN(n722) );
  XNOR2_X1 U791 ( .A(n722), .B(KEYINPUT90), .ZN(n724) );
  NAND2_X1 U792 ( .A1(n892), .A2(G129), .ZN(n723) );
  NAND2_X1 U793 ( .A1(n724), .A2(n723), .ZN(n727) );
  NAND2_X1 U794 ( .A1(G141), .A2(n889), .ZN(n725) );
  XNOR2_X1 U795 ( .A(KEYINPUT91), .B(n725), .ZN(n726) );
  NOR2_X1 U796 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U797 ( .A1(n729), .A2(n728), .ZN(n880) );
  NAND2_X1 U798 ( .A1(G1996), .A2(n880), .ZN(n730) );
  XOR2_X1 U799 ( .A(KEYINPUT92), .B(n730), .Z(n739) );
  NAND2_X1 U800 ( .A1(n894), .A2(G107), .ZN(n732) );
  NAND2_X1 U801 ( .A1(G131), .A2(n889), .ZN(n731) );
  NAND2_X1 U802 ( .A1(n732), .A2(n731), .ZN(n735) );
  NAND2_X1 U803 ( .A1(G119), .A2(n892), .ZN(n733) );
  XNOR2_X1 U804 ( .A(KEYINPUT89), .B(n733), .ZN(n734) );
  NOR2_X1 U805 ( .A1(n735), .A2(n734), .ZN(n737) );
  NAND2_X1 U806 ( .A1(n888), .A2(G95), .ZN(n736) );
  NAND2_X1 U807 ( .A1(n737), .A2(n736), .ZN(n879) );
  AND2_X1 U808 ( .A1(n879), .A2(G1991), .ZN(n738) );
  NOR2_X1 U809 ( .A1(n739), .A2(n738), .ZN(n926) );
  INV_X1 U810 ( .A(n755), .ZN(n740) );
  NOR2_X1 U811 ( .A1(n926), .A2(n740), .ZN(n747) );
  INV_X1 U812 ( .A(n747), .ZN(n741) );
  XNOR2_X1 U813 ( .A(G1986), .B(G290), .ZN(n983) );
  NAND2_X1 U814 ( .A1(n983), .A2(n755), .ZN(n742) );
  OR2_X1 U815 ( .A1(n744), .A2(n743), .ZN(n758) );
  NOR2_X1 U816 ( .A1(G1996), .A2(n880), .ZN(n934) );
  NOR2_X1 U817 ( .A1(G1986), .A2(G290), .ZN(n745) );
  NOR2_X1 U818 ( .A1(G1991), .A2(n879), .ZN(n924) );
  NOR2_X1 U819 ( .A1(n745), .A2(n924), .ZN(n746) );
  NOR2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U821 ( .A1(n934), .A2(n748), .ZN(n749) );
  XNOR2_X1 U822 ( .A(KEYINPUT39), .B(n749), .ZN(n751) );
  NAND2_X1 U823 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U824 ( .A(n752), .B(KEYINPUT102), .ZN(n754) );
  NAND2_X1 U825 ( .A1(n901), .A2(n753), .ZN(n920) );
  NAND2_X1 U826 ( .A1(n754), .A2(n920), .ZN(n756) );
  NAND2_X1 U827 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U828 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U829 ( .A(n759), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U830 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U831 ( .A1(n894), .A2(G111), .ZN(n761) );
  NAND2_X1 U832 ( .A1(G135), .A2(n889), .ZN(n760) );
  NAND2_X1 U833 ( .A1(n761), .A2(n760), .ZN(n764) );
  NAND2_X1 U834 ( .A1(n892), .A2(G123), .ZN(n762) );
  XOR2_X1 U835 ( .A(KEYINPUT18), .B(n762), .Z(n763) );
  NOR2_X1 U836 ( .A1(n764), .A2(n763), .ZN(n766) );
  NAND2_X1 U837 ( .A1(n888), .A2(G99), .ZN(n765) );
  NAND2_X1 U838 ( .A1(n766), .A2(n765), .ZN(n921) );
  XNOR2_X1 U839 ( .A(G2096), .B(n921), .ZN(n767) );
  OR2_X1 U840 ( .A1(G2100), .A2(n767), .ZN(G156) );
  INV_X1 U841 ( .A(G57), .ZN(G237) );
  INV_X1 U842 ( .A(G132), .ZN(G219) );
  INV_X1 U843 ( .A(G82), .ZN(G220) );
  NAND2_X1 U844 ( .A1(G7), .A2(G661), .ZN(n768) );
  XNOR2_X1 U845 ( .A(n768), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U846 ( .A(G223), .ZN(n824) );
  NAND2_X1 U847 ( .A1(n824), .A2(G567), .ZN(n769) );
  XOR2_X1 U848 ( .A(KEYINPUT11), .B(n769), .Z(G234) );
  NAND2_X1 U849 ( .A1(G860), .A2(n969), .ZN(G153) );
  NAND2_X1 U850 ( .A1(G868), .A2(G301), .ZN(n771) );
  INV_X1 U851 ( .A(G868), .ZN(n808) );
  NAND2_X1 U852 ( .A1(n975), .A2(n808), .ZN(n770) );
  NAND2_X1 U853 ( .A1(n771), .A2(n770), .ZN(G284) );
  XNOR2_X1 U854 ( .A(KEYINPUT75), .B(G868), .ZN(n772) );
  NOR2_X1 U855 ( .A1(G286), .A2(n772), .ZN(n773) );
  XNOR2_X1 U856 ( .A(n773), .B(KEYINPUT76), .ZN(n775) );
  NOR2_X1 U857 ( .A1(G299), .A2(G868), .ZN(n774) );
  NOR2_X1 U858 ( .A1(n775), .A2(n774), .ZN(G297) );
  INV_X1 U859 ( .A(G559), .ZN(n776) );
  NOR2_X1 U860 ( .A1(G860), .A2(n776), .ZN(n777) );
  XNOR2_X1 U861 ( .A(KEYINPUT77), .B(n777), .ZN(n778) );
  INV_X1 U862 ( .A(n975), .ZN(n794) );
  NAND2_X1 U863 ( .A1(n778), .A2(n794), .ZN(n779) );
  XNOR2_X1 U864 ( .A(n779), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U865 ( .A1(n794), .A2(G868), .ZN(n780) );
  NOR2_X1 U866 ( .A1(G559), .A2(n780), .ZN(n782) );
  AND2_X1 U867 ( .A1(n969), .A2(n808), .ZN(n781) );
  NOR2_X1 U868 ( .A1(n782), .A2(n781), .ZN(G282) );
  NAND2_X1 U869 ( .A1(G93), .A2(n783), .ZN(n786) );
  NAND2_X1 U870 ( .A1(G80), .A2(n784), .ZN(n785) );
  NAND2_X1 U871 ( .A1(n786), .A2(n785), .ZN(n793) );
  NAND2_X1 U872 ( .A1(n787), .A2(G55), .ZN(n790) );
  NAND2_X1 U873 ( .A1(G67), .A2(n788), .ZN(n789) );
  NAND2_X1 U874 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U875 ( .A(KEYINPUT79), .B(n791), .Z(n792) );
  OR2_X1 U876 ( .A1(n793), .A2(n792), .ZN(n807) );
  NAND2_X1 U877 ( .A1(G559), .A2(n794), .ZN(n795) );
  XOR2_X1 U878 ( .A(n969), .B(n795), .Z(n805) );
  XNOR2_X1 U879 ( .A(KEYINPUT78), .B(n805), .ZN(n796) );
  NOR2_X1 U880 ( .A1(G860), .A2(n796), .ZN(n797) );
  XOR2_X1 U881 ( .A(n807), .B(n797), .Z(G145) );
  XOR2_X1 U882 ( .A(G305), .B(n807), .Z(n804) );
  XOR2_X1 U883 ( .A(KEYINPUT19), .B(KEYINPUT83), .Z(n798) );
  XNOR2_X1 U884 ( .A(G288), .B(n798), .ZN(n799) );
  XNOR2_X1 U885 ( .A(G166), .B(n799), .ZN(n802) );
  XNOR2_X1 U886 ( .A(G290), .B(n800), .ZN(n801) );
  XNOR2_X1 U887 ( .A(n802), .B(n801), .ZN(n803) );
  XNOR2_X1 U888 ( .A(n804), .B(n803), .ZN(n907) );
  XNOR2_X1 U889 ( .A(n805), .B(n907), .ZN(n806) );
  NAND2_X1 U890 ( .A1(n806), .A2(G868), .ZN(n810) );
  NAND2_X1 U891 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U892 ( .A1(n810), .A2(n809), .ZN(G295) );
  NAND2_X1 U893 ( .A1(G2078), .A2(G2084), .ZN(n811) );
  XOR2_X1 U894 ( .A(KEYINPUT20), .B(n811), .Z(n812) );
  NAND2_X1 U895 ( .A1(G2090), .A2(n812), .ZN(n814) );
  XNOR2_X1 U896 ( .A(KEYINPUT84), .B(KEYINPUT21), .ZN(n813) );
  XNOR2_X1 U897 ( .A(n814), .B(n813), .ZN(n815) );
  NAND2_X1 U898 ( .A1(G2072), .A2(n815), .ZN(G158) );
  XNOR2_X1 U899 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U900 ( .A1(G220), .A2(G219), .ZN(n816) );
  XOR2_X1 U901 ( .A(KEYINPUT22), .B(n816), .Z(n817) );
  NOR2_X1 U902 ( .A1(G218), .A2(n817), .ZN(n818) );
  NAND2_X1 U903 ( .A1(G96), .A2(n818), .ZN(n829) );
  NAND2_X1 U904 ( .A1(n829), .A2(G2106), .ZN(n822) );
  NAND2_X1 U905 ( .A1(G69), .A2(G120), .ZN(n819) );
  NOR2_X1 U906 ( .A1(G237), .A2(n819), .ZN(n820) );
  NAND2_X1 U907 ( .A1(G108), .A2(n820), .ZN(n830) );
  NAND2_X1 U908 ( .A1(n830), .A2(G567), .ZN(n821) );
  NAND2_X1 U909 ( .A1(n822), .A2(n821), .ZN(n841) );
  NAND2_X1 U910 ( .A1(G483), .A2(G661), .ZN(n823) );
  NOR2_X1 U911 ( .A1(n841), .A2(n823), .ZN(n828) );
  NAND2_X1 U912 ( .A1(n828), .A2(G36), .ZN(G176) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n824), .ZN(G217) );
  NAND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n825) );
  XNOR2_X1 U915 ( .A(KEYINPUT105), .B(n825), .ZN(n826) );
  NAND2_X1 U916 ( .A1(n826), .A2(G661), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U918 ( .A1(n828), .A2(n827), .ZN(G188) );
  INV_X1 U920 ( .A(G120), .ZN(G236) );
  INV_X1 U921 ( .A(G96), .ZN(G221) );
  INV_X1 U922 ( .A(G69), .ZN(G235) );
  NOR2_X1 U923 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U924 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U925 ( .A(G1341), .B(G2454), .ZN(n831) );
  XNOR2_X1 U926 ( .A(n831), .B(G2430), .ZN(n832) );
  XNOR2_X1 U927 ( .A(n832), .B(G1348), .ZN(n838) );
  XOR2_X1 U928 ( .A(G2443), .B(G2427), .Z(n834) );
  XNOR2_X1 U929 ( .A(G2438), .B(G2446), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n834), .B(n833), .ZN(n836) );
  XOR2_X1 U931 ( .A(G2451), .B(G2435), .Z(n835) );
  XNOR2_X1 U932 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U933 ( .A(n838), .B(n837), .ZN(n839) );
  NAND2_X1 U934 ( .A1(n839), .A2(G14), .ZN(n840) );
  XNOR2_X1 U935 ( .A(KEYINPUT103), .B(n840), .ZN(n915) );
  XNOR2_X1 U936 ( .A(n915), .B(KEYINPUT104), .ZN(G401) );
  INV_X1 U937 ( .A(n841), .ZN(G319) );
  XOR2_X1 U938 ( .A(KEYINPUT43), .B(G2678), .Z(n843) );
  XNOR2_X1 U939 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U941 ( .A(KEYINPUT42), .B(G2090), .Z(n845) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2072), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U944 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U945 ( .A(G2096), .B(G2100), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(n851) );
  XOR2_X1 U947 ( .A(G2078), .B(G2084), .Z(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(G227) );
  XOR2_X1 U949 ( .A(G1976), .B(G1971), .Z(n853) );
  XNOR2_X1 U950 ( .A(G1966), .B(G1961), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U952 ( .A(n854), .B(G2474), .Z(n856) );
  XNOR2_X1 U953 ( .A(G1986), .B(G1956), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U955 ( .A(KEYINPUT41), .B(G1981), .Z(n858) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(G229) );
  NAND2_X1 U959 ( .A1(n888), .A2(G100), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n861), .B(KEYINPUT108), .ZN(n863) );
  NAND2_X1 U961 ( .A1(G112), .A2(n894), .ZN(n862) );
  NAND2_X1 U962 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n864), .B(KEYINPUT109), .ZN(n866) );
  NAND2_X1 U964 ( .A1(G136), .A2(n889), .ZN(n865) );
  NAND2_X1 U965 ( .A1(n866), .A2(n865), .ZN(n869) );
  NAND2_X1 U966 ( .A1(n892), .A2(G124), .ZN(n867) );
  XOR2_X1 U967 ( .A(KEYINPUT44), .B(n867), .Z(n868) );
  NOR2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U969 ( .A(KEYINPUT110), .B(n870), .ZN(G162) );
  NAND2_X1 U970 ( .A1(G130), .A2(n892), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G118), .A2(n894), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n878) );
  NAND2_X1 U973 ( .A1(G106), .A2(n888), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G142), .A2(n889), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U976 ( .A(KEYINPUT111), .B(n875), .ZN(n876) );
  XNOR2_X1 U977 ( .A(KEYINPUT45), .B(n876), .ZN(n877) );
  NOR2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n887) );
  XNOR2_X1 U979 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n882) );
  XOR2_X1 U980 ( .A(n880), .B(n879), .Z(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n921), .B(n883), .ZN(n885) );
  XNOR2_X1 U983 ( .A(G164), .B(G160), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n903) );
  NAND2_X1 U986 ( .A1(G103), .A2(n888), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G139), .A2(n889), .ZN(n890) );
  NAND2_X1 U988 ( .A1(n891), .A2(n890), .ZN(n900) );
  NAND2_X1 U989 ( .A1(n892), .A2(G127), .ZN(n893) );
  XNOR2_X1 U990 ( .A(n893), .B(KEYINPUT112), .ZN(n896) );
  NAND2_X1 U991 ( .A1(G115), .A2(n894), .ZN(n895) );
  NAND2_X1 U992 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U993 ( .A(KEYINPUT47), .B(n897), .ZN(n898) );
  XNOR2_X1 U994 ( .A(KEYINPUT113), .B(n898), .ZN(n899) );
  NOR2_X1 U995 ( .A1(n900), .A2(n899), .ZN(n927) );
  XNOR2_X1 U996 ( .A(n901), .B(n927), .ZN(n902) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U998 ( .A(n904), .B(G162), .ZN(n905) );
  NOR2_X1 U999 ( .A1(G37), .A2(n905), .ZN(G395) );
  XNOR2_X1 U1000 ( .A(KEYINPUT114), .B(n969), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n906), .B(n975), .ZN(n908) );
  XOR2_X1 U1002 ( .A(n908), .B(n907), .Z(n910) );
  XNOR2_X1 U1003 ( .A(G171), .B(G286), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n910), .B(n909), .ZN(n911) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n911), .ZN(G397) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n912) );
  XOR2_X1 U1007 ( .A(KEYINPUT49), .B(n912), .Z(n913) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n913), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1011 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  INV_X1 U1014 ( .A(n918), .ZN(n919) );
  NAND2_X1 U1015 ( .A1(n920), .A2(n919), .ZN(n940) );
  XNOR2_X1 U1016 ( .A(G160), .B(G2084), .ZN(n922) );
  NAND2_X1 U1017 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1018 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1019 ( .A1(n926), .A2(n925), .ZN(n933) );
  XNOR2_X1 U1020 ( .A(G2072), .B(n927), .ZN(n929) );
  XNOR2_X1 U1021 ( .A(G164), .B(G2078), .ZN(n928) );
  NAND2_X1 U1022 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1023 ( .A(KEYINPUT115), .B(n930), .Z(n931) );
  XNOR2_X1 U1024 ( .A(KEYINPUT50), .B(n931), .ZN(n932) );
  NOR2_X1 U1025 ( .A1(n933), .A2(n932), .ZN(n938) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n935) );
  NOR2_X1 U1027 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1028 ( .A(KEYINPUT51), .B(n936), .Z(n937) );
  NAND2_X1 U1029 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1030 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1031 ( .A(KEYINPUT52), .B(n941), .ZN(n943) );
  INV_X1 U1032 ( .A(KEYINPUT55), .ZN(n942) );
  NAND2_X1 U1033 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1034 ( .A1(n944), .A2(G29), .ZN(n1027) );
  XNOR2_X1 U1035 ( .A(G29), .B(KEYINPUT119), .ZN(n967) );
  XNOR2_X1 U1036 ( .A(G2084), .B(G34), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(n945), .B(KEYINPUT54), .ZN(n964) );
  XNOR2_X1 U1038 ( .A(G32), .B(n946), .ZN(n954) );
  XNOR2_X1 U1039 ( .A(G1991), .B(G25), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(G2072), .B(G33), .ZN(n947) );
  NOR2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1042 ( .A1(G28), .A2(n949), .ZN(n952) );
  XNOR2_X1 U1043 ( .A(KEYINPUT116), .B(G2067), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(G26), .B(n950), .ZN(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1046 ( .A1(n954), .A2(n953), .ZN(n957) );
  XNOR2_X1 U1047 ( .A(G27), .B(n955), .ZN(n956) );
  NOR2_X1 U1048 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1049 ( .A(n958), .B(KEYINPUT117), .Z(n959) );
  XNOR2_X1 U1050 ( .A(KEYINPUT53), .B(n959), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(G35), .B(G2090), .ZN(n960) );
  NOR2_X1 U1052 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1053 ( .A(KEYINPUT118), .B(n962), .Z(n963) );
  NOR2_X1 U1054 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1055 ( .A(KEYINPUT55), .B(n965), .ZN(n966) );
  NAND2_X1 U1056 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n968), .ZN(n1025) );
  XNOR2_X1 U1058 ( .A(G16), .B(KEYINPUT56), .ZN(n995) );
  XOR2_X1 U1059 ( .A(n969), .B(G1341), .Z(n974) );
  XOR2_X1 U1060 ( .A(G168), .B(G1966), .Z(n970) );
  NOR2_X1 U1061 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1062 ( .A(KEYINPUT57), .B(n972), .ZN(n973) );
  NOR2_X1 U1063 ( .A1(n974), .A2(n973), .ZN(n993) );
  XNOR2_X1 U1064 ( .A(G301), .B(G1961), .ZN(n977) );
  XNOR2_X1 U1065 ( .A(n975), .B(G1348), .ZN(n976) );
  NOR2_X1 U1066 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1067 ( .A(KEYINPUT120), .B(n978), .Z(n991) );
  NAND2_X1 U1068 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1069 ( .A(n981), .B(KEYINPUT121), .ZN(n985) );
  XNOR2_X1 U1070 ( .A(G1956), .B(G299), .ZN(n982) );
  NOR2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1072 ( .A1(n985), .A2(n984), .ZN(n988) );
  XNOR2_X1 U1073 ( .A(G1971), .B(G303), .ZN(n986) );
  XNOR2_X1 U1074 ( .A(KEYINPUT122), .B(n986), .ZN(n987) );
  NOR2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(KEYINPUT123), .B(n989), .ZN(n990) );
  NOR2_X1 U1077 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1078 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1079 ( .A1(n995), .A2(n994), .ZN(n1023) );
  INV_X1 U1080 ( .A(G16), .ZN(n1021) );
  XNOR2_X1 U1081 ( .A(KEYINPUT125), .B(G1981), .ZN(n996) );
  XNOR2_X1 U1082 ( .A(n996), .B(G6), .ZN(n1001) );
  XOR2_X1 U1083 ( .A(G1348), .B(KEYINPUT59), .Z(n997) );
  XNOR2_X1 U1084 ( .A(G4), .B(n997), .ZN(n999) );
  XNOR2_X1 U1085 ( .A(G20), .B(G1956), .ZN(n998) );
  NOR2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1004) );
  XNOR2_X1 U1088 ( .A(G19), .B(G1341), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(KEYINPUT124), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(KEYINPUT60), .B(n1005), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(n1006), .B(KEYINPUT126), .ZN(n1010) );
  XNOR2_X1 U1093 ( .A(G1966), .B(G21), .ZN(n1008) );
  XNOR2_X1 U1094 ( .A(G5), .B(G1961), .ZN(n1007) );
  NOR2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1018) );
  XOR2_X1 U1097 ( .A(G1986), .B(G24), .Z(n1014) );
  XNOR2_X1 U1098 ( .A(G1971), .B(G22), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(G23), .B(G1976), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(KEYINPUT127), .B(n1015), .Z(n1016) );
  XNOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(KEYINPUT61), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1109 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

