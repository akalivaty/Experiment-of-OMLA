//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n451, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n536, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1156, new_n1157;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g024(.A(G2106), .ZN(new_n450));
  NOR2_X1   g025(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT67), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n454), .A2(new_n450), .B1(new_n458), .B2(new_n455), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT68), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT69), .ZN(new_n464));
  OAI21_X1  g039(.A(G2105), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G101), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n465), .A2(new_n475), .ZN(G160));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n477), .B1(new_n471), .B2(new_n474), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n461), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT71), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n461), .A2(new_n474), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G112), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n467), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n484), .A2(G136), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND4_X1  g065(.A1(new_n468), .A2(new_n470), .A3(KEYINPUT4), .A4(G138), .ZN(new_n491));
  NAND2_X1  g066(.A1(G102), .A2(G2104), .ZN(new_n492));
  AOI21_X1  g067(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(G114), .A2(G2104), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n461), .B2(G126), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n496), .B2(new_n474), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n484), .A2(G138), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n493), .B1(new_n497), .B2(new_n498), .ZN(G164));
  XNOR2_X1  g074(.A(KEYINPUT5), .B(G543), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT6), .B(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G88), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n502), .A2(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n506), .A2(new_n509), .ZN(G303));
  INV_X1    g085(.A(G303), .ZN(G166));
  NAND3_X1  g086(.A1(new_n500), .A2(G63), .A3(G651), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n512), .B(KEYINPUT72), .ZN(new_n513));
  INV_X1    g088(.A(new_n504), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G51), .ZN(new_n515));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  INV_X1    g092(.A(new_n502), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G89), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n513), .A2(new_n515), .A3(new_n517), .A4(new_n519), .ZN(G286));
  INV_X1    g095(.A(G286), .ZN(G168));
  INV_X1    g096(.A(G90), .ZN(new_n522));
  INV_X1    g097(.A(G52), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n502), .A2(new_n522), .B1(new_n504), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n508), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n524), .A2(new_n526), .ZN(G301));
  INV_X1    g102(.A(G301), .ZN(G171));
  INV_X1    g103(.A(G81), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT73), .B(G43), .Z(new_n530));
  OAI22_X1  g105(.A1(new_n502), .A2(new_n529), .B1(new_n504), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n508), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G860), .ZN(G153));
  AND3_X1   g110(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G36), .ZN(G176));
  NAND2_X1  g112(.A1(G1), .A2(G3), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT8), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g115(.A(new_n540), .B(KEYINPUT74), .Z(G188));
  NAND3_X1  g116(.A1(new_n501), .A2(G53), .A3(G543), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT9), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n542), .B(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n500), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G91), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n545), .A2(new_n508), .B1(new_n502), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(G299));
  NAND2_X1  g124(.A1(new_n518), .A2(G87), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n514), .A2(G49), .ZN(new_n551));
  OAI21_X1  g126(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(G288));
  INV_X1    g128(.A(G86), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT77), .B1(new_n502), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n500), .A2(new_n501), .A3(new_n556), .A4(G86), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n558));
  INV_X1    g133(.A(G48), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n504), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n501), .A2(KEYINPUT78), .A3(G48), .A4(G543), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n555), .A2(new_n557), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT5), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT5), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G543), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n566), .A3(G61), .ZN(new_n567));
  NAND2_X1  g142(.A1(G73), .A2(G543), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(KEYINPUT75), .B1(new_n569), .B2(G651), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  AOI211_X1 g146(.A(new_n571), .B(new_n508), .C1(new_n567), .C2(new_n568), .ZN(new_n572));
  NOR3_X1   g147(.A1(new_n570), .A2(new_n572), .A3(KEYINPUT76), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  INV_X1    g149(.A(new_n568), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n500), .B2(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n571), .B1(new_n576), .B2(new_n508), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n569), .A2(KEYINPUT75), .A3(G651), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n574), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n562), .B1(new_n573), .B2(new_n579), .ZN(G305));
  INV_X1    g155(.A(G85), .ZN(new_n581));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n502), .A2(new_n581), .B1(new_n504), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT79), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n584), .A2(KEYINPUT79), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n586), .A2(new_n587), .B1(new_n508), .B2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT80), .Z(new_n591));
  INV_X1    g166(.A(G92), .ZN(new_n592));
  OR3_X1    g167(.A1(new_n502), .A2(KEYINPUT81), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(KEYINPUT81), .B1(new_n502), .B2(new_n592), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n500), .A2(G66), .ZN(new_n598));
  INV_X1    g173(.A(G79), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(new_n563), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n600), .A2(G651), .B1(G54), .B2(new_n514), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n593), .A2(KEYINPUT10), .A3(new_n594), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n591), .B1(G868), .B2(new_n603), .ZN(G321));
  XNOR2_X1  g179(.A(G321), .B(KEYINPUT82), .ZN(G284));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G868), .B2(new_n548), .ZN(G280));
  XNOR2_X1  g182(.A(G280), .B(KEYINPUT83), .ZN(G297));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n603), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n603), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n534), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n484), .A2(G2104), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT12), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  INV_X1    g192(.A(G2100), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n480), .A2(G123), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n484), .A2(G135), .ZN(new_n621));
  NOR2_X1   g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(new_n474), .B2(G111), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n619), .A2(new_n625), .ZN(G156));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2435), .ZN(new_n628));
  XOR2_X1   g203(.A(G2427), .B(G2438), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT14), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2451), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n631), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n637), .B(new_n638), .Z(new_n639));
  AND2_X1   g214(.A1(new_n639), .A2(G14), .ZN(G401));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT85), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  NOR3_X1   g221(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT18), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n643), .A2(new_n644), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n644), .B(KEYINPUT17), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n649), .B(new_n646), .C1(new_n643), .C2(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n643), .A2(new_n650), .A3(new_n645), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n648), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2096), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(new_n618), .ZN(G227));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT20), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n657), .A2(new_n660), .A3(new_n662), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n665), .B(new_n666), .C1(new_n664), .C2(new_n663), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT86), .B(KEYINPUT87), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  INV_X1    g245(.A(G1981), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(G229));
  XNOR2_X1  g251(.A(KEYINPUT31), .B(G11), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n603), .A2(G16), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(G4), .B2(G16), .ZN(new_n679));
  INV_X1    g254(.A(G1348), .ZN(new_n680));
  INV_X1    g255(.A(G29), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT30), .B(G28), .ZN(new_n682));
  AOI22_X1  g257(.A1(new_n679), .A2(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AND2_X1   g258(.A1(KEYINPUT88), .A2(G29), .ZN(new_n684));
  NOR2_X1   g259(.A1(KEYINPUT88), .A2(G29), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n624), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G5), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G171), .B2(new_n689), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT98), .B(G1961), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  AND4_X1   g268(.A1(new_n677), .A2(new_n683), .A3(new_n688), .A4(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n687), .A2(KEYINPUT28), .A3(G26), .ZN(new_n695));
  AOI22_X1  g270(.A1(new_n480), .A2(G128), .B1(G140), .B2(new_n484), .ZN(new_n696));
  OR2_X1    g271(.A1(G104), .A2(G2105), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n697), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n695), .B1(new_n699), .B2(new_n681), .ZN(new_n700));
  AOI21_X1  g275(.A(KEYINPUT28), .B1(new_n687), .B2(G26), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G2067), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(G29), .A2(G32), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT96), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT26), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n480), .A2(G129), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n461), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(G2105), .ZN(new_n712));
  AND3_X1   g287(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n706), .B1(new_n713), .B2(G29), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT27), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1996), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n689), .A2(KEYINPUT23), .A3(G20), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT23), .ZN(new_n718));
  INV_X1    g293(.A(G20), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(G16), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n717), .B(new_n720), .C1(new_n548), .C2(new_n689), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1956), .ZN(new_n722));
  INV_X1    g297(.A(G27), .ZN(new_n723));
  OAI21_X1  g298(.A(KEYINPUT100), .B1(new_n686), .B2(new_n723), .ZN(new_n724));
  OR3_X1    g299(.A1(new_n686), .A2(KEYINPUT100), .A3(new_n723), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n724), .B(new_n725), .C1(G164), .C2(new_n687), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G2078), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n694), .A2(new_n705), .A3(new_n716), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT24), .B(G34), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n687), .A2(KEYINPUT95), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G160), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(new_n681), .ZN(new_n733));
  AOI21_X1  g308(.A(KEYINPUT95), .B1(new_n687), .B2(new_n730), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G2084), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT99), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n679), .A2(new_n680), .ZN(new_n739));
  OR2_X1    g314(.A1(G29), .A2(G33), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n484), .A2(G139), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT25), .Z(new_n743));
  AOI22_X1  g318(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n741), .B(new_n743), .C1(new_n474), .C2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n740), .B1(new_n745), .B2(new_n681), .ZN(new_n746));
  INV_X1    g321(.A(G2072), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(G16), .A2(G21), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G168), .B2(G16), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT97), .B(G1966), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n739), .A2(new_n748), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n689), .A2(G19), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n534), .B2(new_n689), .ZN(new_n755));
  MUX2_X1   g330(.A(new_n754), .B(new_n755), .S(KEYINPUT94), .Z(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(G1341), .Z(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  NOR4_X1   g333(.A1(new_n729), .A2(new_n738), .A3(new_n753), .A4(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n735), .A2(new_n736), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT36), .ZN(new_n761));
  NAND2_X1  g336(.A1(G305), .A2(G16), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n689), .A2(G6), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT32), .B(G1981), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT90), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n766), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n762), .A2(new_n763), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n689), .A2(G23), .ZN(new_n771));
  INV_X1    g346(.A(G288), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(new_n689), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT33), .B(G1976), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT91), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n773), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G16), .A2(G22), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G166), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT92), .B(G1971), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n770), .A2(new_n776), .A3(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT93), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n770), .A2(KEYINPUT93), .A3(new_n776), .A4(new_n780), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(KEYINPUT34), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT34), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n783), .A2(new_n787), .A3(new_n784), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G24), .ZN(new_n790));
  OAI21_X1  g365(.A(KEYINPUT89), .B1(new_n790), .B2(G16), .ZN(new_n791));
  OR3_X1    g366(.A1(new_n790), .A2(KEYINPUT89), .A3(G16), .ZN(new_n792));
  INV_X1    g367(.A(G290), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n791), .B(new_n792), .C1(new_n793), .C2(new_n689), .ZN(new_n794));
  INV_X1    g369(.A(G1986), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n687), .A2(G25), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n480), .A2(G119), .B1(G131), .B2(new_n484), .ZN(new_n798));
  OR2_X1    g373(.A1(G95), .A2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G107), .C2(new_n474), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n797), .B1(new_n801), .B2(new_n687), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT35), .B(G1991), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n802), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n796), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n761), .B1(new_n789), .B2(new_n807), .ZN(new_n808));
  AOI211_X1 g383(.A(KEYINPUT36), .B(new_n806), .C1(new_n786), .C2(new_n788), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n759), .B(new_n760), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n746), .A2(new_n747), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(G162), .A2(new_n687), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G35), .B2(new_n687), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT29), .B(G2090), .Z(new_n815));
  XOR2_X1   g390(.A(new_n814), .B(new_n815), .Z(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n810), .A2(new_n812), .A3(new_n817), .ZN(G311));
  OR3_X1    g393(.A1(new_n810), .A2(new_n812), .A3(new_n817), .ZN(G150));
  INV_X1    g394(.A(G93), .ZN(new_n820));
  INV_X1    g395(.A(G55), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n502), .A2(new_n820), .B1(new_n504), .B2(new_n821), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n823), .A2(new_n508), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G860), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  INV_X1    g403(.A(new_n534), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n825), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n826), .A2(new_n534), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n835), .A2(new_n609), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n834), .B(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n828), .B1(new_n837), .B2(G860), .ZN(G145));
  INV_X1    g413(.A(KEYINPUT40), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n468), .A2(new_n470), .A3(G126), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n474), .B1(new_n840), .B2(new_n494), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT4), .ZN(new_n842));
  INV_X1    g417(.A(G138), .ZN(new_n843));
  OAI22_X1  g418(.A1(new_n841), .A2(new_n842), .B1(new_n843), .B2(new_n483), .ZN(new_n844));
  INV_X1    g419(.A(new_n493), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n699), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n713), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n696), .A2(new_n698), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G164), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n848), .B1(new_n847), .B2(new_n850), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n745), .B(KEYINPUT101), .ZN(new_n853));
  OR3_X1    g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT101), .ZN(new_n855));
  OAI22_X1  g430(.A1(new_n851), .A2(new_n852), .B1(new_n855), .B2(new_n745), .ZN(new_n856));
  INV_X1    g431(.A(G142), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n483), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(new_n480), .B2(G130), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n474), .A2(G118), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(G2104), .ZN(new_n861));
  NOR2_X1   g436(.A1(G106), .A2(G2105), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n801), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n798), .A2(new_n800), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n866), .A2(new_n859), .A3(new_n863), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n868), .B1(new_n865), .B2(new_n867), .ZN(new_n871));
  INV_X1    g446(.A(new_n616), .ZN(new_n872));
  NOR3_X1   g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n865), .A2(new_n867), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT102), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n616), .B1(new_n875), .B2(new_n869), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n854), .B(new_n856), .C1(new_n873), .C2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n616), .A3(new_n869), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n872), .B1(new_n870), .B2(new_n871), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n745), .A2(new_n855), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n847), .A2(new_n850), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n713), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n878), .B(new_n879), .C1(new_n880), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n877), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n624), .B(G160), .ZN(new_n888));
  XNOR2_X1  g463(.A(G162), .B(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(G37), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n877), .A2(new_n886), .A3(new_n889), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT103), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n891), .A2(new_n897), .A3(new_n892), .A4(new_n893), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n896), .B1(new_n895), .B2(new_n898), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n839), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n877), .A2(new_n889), .A3(new_n886), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n889), .B1(new_n877), .B2(new_n886), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n897), .B1(new_n904), .B2(new_n892), .ZN(new_n905));
  INV_X1    g480(.A(new_n898), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT104), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(KEYINPUT40), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n901), .A2(new_n909), .ZN(G395));
  XNOR2_X1  g485(.A(G303), .B(G288), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(G290), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(G305), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n914));
  OAI21_X1  g489(.A(KEYINPUT106), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT42), .ZN(new_n916));
  INV_X1    g491(.A(G305), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n912), .B(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g496(.A(KEYINPUT106), .B(new_n916), .C1(new_n913), .C2(new_n914), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n611), .B(new_n832), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n603), .A2(new_n548), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n835), .A2(G299), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT41), .B1(new_n925), .B2(new_n926), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g508(.A(KEYINPUT105), .B(KEYINPUT41), .C1(new_n925), .C2(new_n926), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n928), .B1(new_n935), .B2(new_n924), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n923), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n923), .A2(new_n936), .ZN(new_n938));
  OAI21_X1  g513(.A(G868), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(G868), .B2(new_n825), .ZN(G295));
  OAI21_X1  g515(.A(new_n939), .B1(G868), .B2(new_n825), .ZN(G331));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n832), .A2(G171), .ZN(new_n943));
  AOI21_X1  g518(.A(G301), .B1(new_n831), .B2(new_n830), .ZN(new_n944));
  OR3_X1    g519(.A1(new_n943), .A2(G286), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(G286), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n933), .A2(new_n934), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n945), .A2(new_n927), .A3(new_n946), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n913), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n892), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n913), .B1(new_n948), .B2(new_n949), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n942), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n930), .A2(KEYINPUT108), .A3(new_n932), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n927), .A2(new_n957), .A3(new_n929), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n947), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n913), .B1(new_n959), .B2(new_n949), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT43), .B1(new_n951), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT109), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n963), .B(KEYINPUT43), .C1(new_n951), .C2(new_n960), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n955), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n960), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n966), .A2(new_n954), .A3(new_n892), .A4(new_n950), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(new_n953), .B2(new_n954), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n942), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n965), .A2(new_n969), .ZN(G397));
  INV_X1    g545(.A(G1384), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n846), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n465), .A2(G40), .A3(new_n475), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n793), .A2(new_n977), .A3(new_n795), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(G1986), .A3(G290), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g555(.A(new_n980), .B(KEYINPUT110), .Z(new_n981));
  XNOR2_X1  g556(.A(new_n849), .B(new_n703), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n848), .A2(G1996), .ZN(new_n983));
  INV_X1    g558(.A(G1996), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n713), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n866), .B(new_n804), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n977), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n981), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n671), .B(new_n562), .C1(new_n573), .C2(new_n579), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n560), .A2(new_n561), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT114), .B(G86), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n518), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n993), .A2(new_n578), .A3(new_n577), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(G1981), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT49), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n976), .A2(new_n972), .ZN(new_n1001));
  INV_X1    g576(.A(G8), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n992), .A2(KEYINPUT49), .A3(new_n997), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1000), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT115), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1000), .A2(new_n1007), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(G288), .A2(G1976), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n1009), .A2(new_n1010), .B1(new_n671), .B2(new_n917), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1003), .ZN(new_n1012));
  INV_X1    g587(.A(new_n972), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n975), .ZN(new_n1014));
  INV_X1    g589(.A(G1976), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT113), .B1(G288), .B2(new_n1015), .ZN(new_n1016));
  OR3_X1    g591(.A1(G288), .A2(KEYINPUT113), .A3(new_n1015), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1014), .A2(G8), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT52), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n772), .A2(G1976), .ZN(new_n1022));
  OR3_X1    g597(.A1(new_n1018), .A2(KEYINPUT52), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n846), .A2(KEYINPUT45), .A3(new_n971), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n974), .A2(new_n975), .A3(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT111), .B(G1971), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n1029));
  NOR3_X1   g604(.A1(G164), .A2(new_n1029), .A3(G1384), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT50), .B1(new_n846), .B2(new_n971), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n975), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1028), .B1(G2090), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(KEYINPUT112), .A2(KEYINPUT55), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(G166), .B2(new_n1002), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n1036));
  NAND3_X1  g611(.A1(G303), .A2(G8), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1033), .A2(G8), .A3(new_n1038), .ZN(new_n1039));
  OAI22_X1  g614(.A1(new_n1011), .A2(new_n1012), .B1(new_n1024), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1038), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1029), .B1(G164), .B2(G1384), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n846), .A2(KEYINPUT50), .A3(new_n971), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n976), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n1045));
  AOI21_X1  g620(.A(G2090), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1032), .A2(KEYINPUT116), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1046), .A2(new_n1047), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1041), .B1(new_n1048), .B2(new_n1002), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1021), .A2(new_n1049), .A3(new_n1039), .A4(new_n1023), .ZN(new_n1050));
  INV_X1    g625(.A(G1966), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1026), .A2(new_n1051), .B1(new_n1044), .B2(new_n736), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT51), .B1(new_n1052), .B2(G168), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1002), .B1(new_n1052), .B2(G168), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1055), .B1(new_n1056), .B2(new_n1054), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT62), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1050), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1044), .A2(G1961), .ZN(new_n1061));
  INV_X1    g636(.A(G2078), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n974), .A2(new_n1062), .A3(new_n975), .A4(new_n1025), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT125), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1063), .A2(new_n1064), .A3(KEYINPUT53), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT53), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1061), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(G171), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(new_n1057), .B2(KEYINPUT62), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1040), .B1(new_n1060), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(KEYINPUT118), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(KEYINPUT118), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n548), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1076), .B(KEYINPUT57), .C1(new_n544), .C2(new_n547), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT56), .B(G2072), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n974), .A2(new_n975), .A3(new_n1025), .A4(new_n1080), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1079), .B(new_n1081), .C1(G1956), .C2(new_n1044), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1081), .B1(G1956), .B2(new_n1044), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1078), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT120), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1087), .A3(new_n1078), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1013), .A2(new_n703), .A3(new_n975), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n1044), .B2(G1348), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n603), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1086), .A2(new_n1088), .B1(KEYINPUT119), .B2(new_n1091), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1091), .A2(KEYINPUT119), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1083), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(KEYINPUT60), .B(new_n1089), .C1(new_n1044), .C2(G1348), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1095), .A2(new_n1096), .A3(new_n835), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n835), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1090), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1101), .A2(KEYINPUT60), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1100), .A2(KEYINPUT124), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT124), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT61), .B1(new_n1085), .B2(new_n1082), .ZN(new_n1106));
  XOR2_X1   g681(.A(KEYINPUT58), .B(G1341), .Z(new_n1107));
  NAND2_X1  g682(.A1(new_n1014), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n974), .A2(new_n984), .A3(new_n975), .A4(new_n1025), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n829), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1111));
  XNOR2_X1  g686(.A(new_n1110), .B(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT61), .B1(new_n1082), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1082), .A2(new_n1113), .ZN(new_n1116));
  AOI211_X1 g691(.A(new_n1106), .B(new_n1112), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1094), .B1(new_n1105), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1058), .A2(new_n1050), .ZN(new_n1119));
  OAI211_X1 g694(.A(G301), .B(new_n1061), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1068), .A2(new_n1120), .ZN(new_n1121));
  OR2_X1    g696(.A1(G171), .A2(KEYINPUT126), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1121), .A2(KEYINPUT54), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1121), .B1(KEYINPUT126), .B2(KEYINPUT54), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1119), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1070), .B1(new_n1118), .B2(new_n1125), .ZN(new_n1126));
  AND4_X1   g701(.A1(new_n1039), .A2(new_n1009), .A3(new_n1019), .A4(new_n1023), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT117), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1052), .A2(new_n1002), .A3(G286), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1127), .A2(new_n1128), .A3(new_n1049), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1129), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT117), .B1(new_n1050), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1130), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1033), .A2(G8), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1133), .B1(new_n1135), .B2(new_n1041), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1127), .A2(new_n1129), .A3(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n991), .B1(new_n1126), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n977), .A2(new_n984), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT46), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT127), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1140), .B(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n982), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n977), .B1(new_n1144), .B2(new_n848), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1143), .B(new_n1145), .C1(KEYINPUT127), .C2(new_n1141), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT47), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n801), .A2(new_n804), .ZN(new_n1148));
  OAI22_X1  g723(.A1(new_n986), .A2(new_n1148), .B1(G2067), .B2(new_n849), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n977), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n978), .B(KEYINPUT48), .Z(new_n1151));
  OAI211_X1 g726(.A(new_n1147), .B(new_n1150), .C1(new_n990), .C2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1139), .A2(new_n1153), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g729(.A1(G401), .A2(G227), .A3(G229), .ZN(new_n1156));
  NAND2_X1  g730(.A1(new_n895), .A2(new_n898), .ZN(new_n1157));
  NAND4_X1  g731(.A1(new_n968), .A2(new_n1156), .A3(new_n1157), .A4(G319), .ZN(G225));
  INV_X1    g732(.A(G225), .ZN(G308));
endmodule


