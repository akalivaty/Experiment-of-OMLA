

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  XNOR2_X1 U324 ( .A(n465), .B(n464), .ZN(n573) );
  XNOR2_X1 U325 ( .A(KEYINPUT100), .B(KEYINPUT26), .ZN(n464) );
  INV_X1 U326 ( .A(n533), .ZN(n535) );
  XOR2_X1 U327 ( .A(n458), .B(n457), .Z(n475) );
  XOR2_X1 U328 ( .A(n445), .B(KEYINPUT64), .Z(n292) );
  XOR2_X1 U329 ( .A(G120GAT), .B(KEYINPUT0), .Z(n293) );
  INV_X1 U330 ( .A(KEYINPUT14), .ZN(n387) );
  XNOR2_X1 U331 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U332 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U333 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U334 ( .A(n415), .B(KEYINPUT48), .ZN(n533) );
  XNOR2_X1 U335 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U336 ( .A(n440), .B(KEYINPUT120), .ZN(n441) );
  AND2_X1 U337 ( .A1(n491), .A2(n481), .ZN(n482) );
  XNOR2_X1 U338 ( .A(n442), .B(n441), .ZN(n459) );
  XOR2_X1 U339 ( .A(KEYINPUT37), .B(n482), .Z(n522) );
  XOR2_X1 U340 ( .A(KEYINPUT112), .B(n586), .Z(n571) );
  XOR2_X1 U341 ( .A(n404), .B(n403), .Z(n586) );
  XOR2_X1 U342 ( .A(n474), .B(KEYINPUT28), .Z(n529) );
  XNOR2_X1 U343 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U344 ( .A(n463), .B(n462), .ZN(G1351GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT11), .B(KEYINPUT65), .Z(n295) );
  XNOR2_X1 U346 ( .A(G106GAT), .B(KEYINPUT66), .ZN(n294) );
  XNOR2_X1 U347 ( .A(n295), .B(n294), .ZN(n311) );
  XNOR2_X1 U348 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n296), .B(KEYINPUT8), .ZN(n368) );
  XOR2_X1 U350 ( .A(G92GAT), .B(KEYINPUT76), .Z(n298) );
  XNOR2_X1 U351 ( .A(G99GAT), .B(G85GAT), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n348) );
  XNOR2_X1 U353 ( .A(n368), .B(n348), .ZN(n309) );
  XOR2_X1 U354 ( .A(KEYINPUT10), .B(KEYINPUT80), .Z(n300) );
  XNOR2_X1 U355 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n299) );
  XOR2_X1 U356 ( .A(n300), .B(n299), .Z(n305) );
  XNOR2_X1 U357 ( .A(G36GAT), .B(G190GAT), .ZN(n301) );
  XNOR2_X1 U358 ( .A(n301), .B(KEYINPUT81), .ZN(n332) );
  XNOR2_X1 U359 ( .A(KEYINPUT79), .B(n332), .ZN(n303) );
  AND2_X1 U360 ( .A1(G232GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U361 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n307) );
  XOR2_X1 U363 ( .A(G43GAT), .B(G134GAT), .Z(n451) );
  XOR2_X1 U364 ( .A(G50GAT), .B(G162GAT), .Z(n313) );
  XNOR2_X1 U365 ( .A(n451), .B(n313), .ZN(n306) );
  XNOR2_X1 U366 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U367 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U368 ( .A(n311), .B(n310), .ZN(n559) );
  INV_X1 U369 ( .A(n559), .ZN(n488) );
  XNOR2_X1 U370 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n312) );
  XNOR2_X1 U371 ( .A(n312), .B(KEYINPUT2), .ZN(n432) );
  XNOR2_X1 U372 ( .A(n313), .B(n432), .ZN(n314) );
  XOR2_X1 U373 ( .A(G22GAT), .B(G155GAT), .Z(n384) );
  XNOR2_X1 U374 ( .A(n314), .B(n384), .ZN(n319) );
  XNOR2_X1 U375 ( .A(G106GAT), .B(G78GAT), .ZN(n315) );
  XNOR2_X1 U376 ( .A(n315), .B(G148GAT), .ZN(n344) );
  XOR2_X1 U377 ( .A(n344), .B(G204GAT), .Z(n317) );
  NAND2_X1 U378 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U380 ( .A(n319), .B(n318), .Z(n327) );
  XOR2_X1 U381 ( .A(KEYINPUT92), .B(G218GAT), .Z(n321) );
  XNOR2_X1 U382 ( .A(KEYINPUT21), .B(KEYINPUT93), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U384 ( .A(G197GAT), .B(n322), .Z(n340) );
  XOR2_X1 U385 ( .A(G211GAT), .B(KEYINPUT24), .Z(n324) );
  XNOR2_X1 U386 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n323) );
  XNOR2_X1 U387 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U388 ( .A(n340), .B(n325), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n327), .B(n326), .ZN(n474) );
  XOR2_X1 U390 ( .A(G204GAT), .B(KEYINPUT77), .Z(n345) );
  XOR2_X1 U391 ( .A(KEYINPUT82), .B(G211GAT), .Z(n329) );
  XNOR2_X1 U392 ( .A(G8GAT), .B(G183GAT), .ZN(n328) );
  XNOR2_X1 U393 ( .A(n329), .B(n328), .ZN(n390) );
  XOR2_X1 U394 ( .A(n345), .B(n390), .Z(n331) );
  XNOR2_X1 U395 ( .A(G92GAT), .B(G64GAT), .ZN(n330) );
  XNOR2_X1 U396 ( .A(n331), .B(n330), .ZN(n336) );
  XOR2_X1 U397 ( .A(KEYINPUT99), .B(n332), .Z(n334) );
  NAND2_X1 U398 ( .A1(G226GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U399 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U400 ( .A(n336), .B(n335), .Z(n343) );
  XOR2_X1 U401 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n338) );
  XNOR2_X1 U402 ( .A(KEYINPUT19), .B(G176GAT), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U404 ( .A(G169GAT), .B(n339), .Z(n458) );
  INV_X1 U405 ( .A(n458), .ZN(n341) );
  XOR2_X1 U406 ( .A(n341), .B(n340), .Z(n342) );
  XNOR2_X1 U407 ( .A(n343), .B(n342), .ZN(n525) );
  XOR2_X1 U408 ( .A(n345), .B(n344), .Z(n347) );
  XNOR2_X1 U409 ( .A(G176GAT), .B(G120GAT), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n347), .B(n346), .ZN(n352) );
  XOR2_X1 U411 ( .A(n348), .B(KEYINPUT33), .Z(n350) );
  NAND2_X1 U412 ( .A1(G230GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U413 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U414 ( .A(n352), .B(n351), .Z(n360) );
  XOR2_X1 U415 ( .A(KEYINPUT74), .B(G64GAT), .Z(n354) );
  XNOR2_X1 U416 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U418 ( .A(G57GAT), .B(n355), .Z(n404) );
  XOR2_X1 U419 ( .A(KEYINPUT75), .B(KEYINPUT31), .Z(n357) );
  XNOR2_X1 U420 ( .A(KEYINPUT32), .B(KEYINPUT78), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n404), .B(n358), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n582) );
  XNOR2_X1 U424 ( .A(KEYINPUT41), .B(n582), .ZN(n565) );
  INV_X1 U425 ( .A(n565), .ZN(n553) );
  XOR2_X1 U426 ( .A(KEYINPUT72), .B(G1GAT), .Z(n396) );
  XOR2_X1 U427 ( .A(G36GAT), .B(G43GAT), .Z(n362) );
  XNOR2_X1 U428 ( .A(G169GAT), .B(G50GAT), .ZN(n361) );
  XNOR2_X1 U429 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U430 ( .A(n396), .B(n363), .Z(n365) );
  NAND2_X1 U431 ( .A1(G229GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U432 ( .A(n365), .B(n364), .ZN(n367) );
  INV_X1 U433 ( .A(G8GAT), .ZN(n366) );
  XNOR2_X1 U434 ( .A(n367), .B(n366), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n368), .B(KEYINPUT30), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U437 ( .A(G141GAT), .B(G197GAT), .Z(n372) );
  XNOR2_X1 U438 ( .A(G15GAT), .B(G113GAT), .ZN(n371) );
  XOR2_X1 U439 ( .A(n372), .B(n371), .Z(n373) );
  XOR2_X1 U440 ( .A(n374), .B(n373), .Z(n382) );
  XOR2_X1 U441 ( .A(KEYINPUT73), .B(KEYINPUT68), .Z(n376) );
  XNOR2_X1 U442 ( .A(KEYINPUT67), .B(KEYINPUT29), .ZN(n375) );
  XNOR2_X1 U443 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U444 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n378) );
  XNOR2_X1 U445 ( .A(G22GAT), .B(KEYINPUT71), .ZN(n377) );
  XNOR2_X1 U446 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U447 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U448 ( .A(n382), .B(n381), .ZN(n576) );
  NAND2_X1 U449 ( .A1(n553), .A2(n576), .ZN(n383) );
  XNOR2_X1 U450 ( .A(KEYINPUT46), .B(n383), .ZN(n405) );
  XOR2_X1 U451 ( .A(KEYINPUT84), .B(n384), .Z(n386) );
  XOR2_X1 U452 ( .A(G15GAT), .B(G127GAT), .Z(n449) );
  XNOR2_X1 U453 ( .A(n449), .B(G78GAT), .ZN(n385) );
  XNOR2_X1 U454 ( .A(n386), .B(n385), .ZN(n392) );
  NAND2_X1 U455 ( .A1(G231GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U456 ( .A(n392), .B(n391), .ZN(n397) );
  XOR2_X1 U457 ( .A(KEYINPUT83), .B(KEYINPUT85), .Z(n394) );
  XNOR2_X1 U458 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n393) );
  XNOR2_X1 U459 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U460 ( .A(n396), .B(n395), .Z(n398) );
  NAND2_X1 U461 ( .A1(n397), .A2(n398), .ZN(n402) );
  INV_X1 U462 ( .A(n397), .ZN(n400) );
  INV_X1 U463 ( .A(n398), .ZN(n399) );
  NAND2_X1 U464 ( .A1(n400), .A2(n399), .ZN(n401) );
  NAND2_X1 U465 ( .A1(n402), .A2(n401), .ZN(n403) );
  NAND2_X1 U466 ( .A1(n405), .A2(n571), .ZN(n406) );
  NOR2_X1 U467 ( .A1(n559), .A2(n406), .ZN(n408) );
  XNOR2_X1 U468 ( .A(KEYINPUT47), .B(KEYINPUT113), .ZN(n407) );
  XNOR2_X1 U469 ( .A(n408), .B(n407), .ZN(n414) );
  INV_X1 U470 ( .A(n576), .ZN(n563) );
  XOR2_X1 U471 ( .A(KEYINPUT45), .B(KEYINPUT114), .Z(n410) );
  XNOR2_X1 U472 ( .A(n559), .B(KEYINPUT36), .ZN(n588) );
  NAND2_X1 U473 ( .A1(n588), .A2(n586), .ZN(n409) );
  XNOR2_X1 U474 ( .A(n410), .B(n409), .ZN(n411) );
  NAND2_X1 U475 ( .A1(n563), .A2(n411), .ZN(n412) );
  NOR2_X1 U476 ( .A1(n582), .A2(n412), .ZN(n413) );
  NOR2_X1 U477 ( .A1(n414), .A2(n413), .ZN(n415) );
  NOR2_X1 U478 ( .A1(n525), .A2(n533), .ZN(n416) );
  XNOR2_X1 U479 ( .A(n416), .B(KEYINPUT54), .ZN(n439) );
  NAND2_X1 U480 ( .A1(G225GAT), .A2(G233GAT), .ZN(n422) );
  XOR2_X1 U481 ( .A(G85GAT), .B(G148GAT), .Z(n418) );
  XNOR2_X1 U482 ( .A(G29GAT), .B(G127GAT), .ZN(n417) );
  XNOR2_X1 U483 ( .A(n418), .B(n417), .ZN(n420) );
  XOR2_X1 U484 ( .A(G134GAT), .B(G162GAT), .Z(n419) );
  XNOR2_X1 U485 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n438) );
  XOR2_X1 U487 ( .A(KEYINPUT95), .B(KEYINPUT1), .Z(n424) );
  XNOR2_X1 U488 ( .A(KEYINPUT4), .B(KEYINPUT98), .ZN(n423) );
  XNOR2_X1 U489 ( .A(n424), .B(n423), .ZN(n436) );
  XOR2_X1 U490 ( .A(KEYINPUT96), .B(G57GAT), .Z(n426) );
  XNOR2_X1 U491 ( .A(G1GAT), .B(G155GAT), .ZN(n425) );
  XNOR2_X1 U492 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U493 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n428) );
  XNOR2_X1 U494 ( .A(KEYINPUT97), .B(KEYINPUT94), .ZN(n427) );
  XNOR2_X1 U495 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U496 ( .A(n430), .B(n429), .Z(n434) );
  XNOR2_X1 U497 ( .A(G113GAT), .B(KEYINPUT87), .ZN(n431) );
  XNOR2_X1 U498 ( .A(n293), .B(n431), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n445), .B(n432), .ZN(n433) );
  XNOR2_X1 U500 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U501 ( .A(n436), .B(n435), .Z(n437) );
  XNOR2_X1 U502 ( .A(n438), .B(n437), .ZN(n523) );
  NAND2_X1 U503 ( .A1(n439), .A2(n523), .ZN(n574) );
  NOR2_X1 U504 ( .A1(n474), .A2(n574), .ZN(n442) );
  INV_X1 U505 ( .A(KEYINPUT55), .ZN(n440) );
  XOR2_X1 U506 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n444) );
  XNOR2_X1 U507 ( .A(G183GAT), .B(KEYINPUT20), .ZN(n443) );
  XNOR2_X1 U508 ( .A(n444), .B(n443), .ZN(n456) );
  NAND2_X1 U509 ( .A1(G227GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U510 ( .A(n292), .B(n446), .ZN(n454) );
  XOR2_X1 U511 ( .A(G71GAT), .B(KEYINPUT88), .Z(n448) );
  XNOR2_X1 U512 ( .A(G190GAT), .B(G99GAT), .ZN(n447) );
  XNOR2_X1 U513 ( .A(n448), .B(n447), .ZN(n450) );
  XOR2_X1 U514 ( .A(n450), .B(n449), .Z(n452) );
  XOR2_X1 U515 ( .A(n456), .B(n455), .Z(n457) );
  NAND2_X1 U516 ( .A1(n459), .A2(n475), .ZN(n570) );
  NOR2_X1 U517 ( .A1(n488), .A2(n570), .ZN(n463) );
  XNOR2_X1 U518 ( .A(KEYINPUT122), .B(KEYINPUT58), .ZN(n461) );
  INV_X1 U519 ( .A(G190GAT), .ZN(n460) );
  INV_X1 U520 ( .A(G43GAT), .ZN(n487) );
  INV_X1 U521 ( .A(n475), .ZN(n536) );
  NAND2_X1 U522 ( .A1(n536), .A2(n474), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n525), .B(KEYINPUT27), .ZN(n473) );
  NOR2_X1 U524 ( .A1(n573), .A2(n473), .ZN(n466) );
  XNOR2_X1 U525 ( .A(KEYINPUT101), .B(n466), .ZN(n470) );
  NOR2_X1 U526 ( .A1(n525), .A2(n536), .ZN(n467) );
  NOR2_X1 U527 ( .A1(n474), .A2(n467), .ZN(n468) );
  XNOR2_X1 U528 ( .A(KEYINPUT25), .B(n468), .ZN(n469) );
  NAND2_X1 U529 ( .A1(n470), .A2(n469), .ZN(n471) );
  NAND2_X1 U530 ( .A1(n471), .A2(n523), .ZN(n472) );
  XNOR2_X1 U531 ( .A(n472), .B(KEYINPUT102), .ZN(n479) );
  NOR2_X1 U532 ( .A1(n523), .A2(n473), .ZN(n534) );
  INV_X1 U533 ( .A(n529), .ZN(n539) );
  XOR2_X1 U534 ( .A(KEYINPUT91), .B(n475), .Z(n476) );
  NOR2_X1 U535 ( .A1(n539), .A2(n476), .ZN(n477) );
  NAND2_X1 U536 ( .A1(n534), .A2(n477), .ZN(n478) );
  NAND2_X1 U537 ( .A1(n479), .A2(n478), .ZN(n491) );
  INV_X1 U538 ( .A(n586), .ZN(n480) );
  AND2_X1 U539 ( .A1(n480), .A2(n588), .ZN(n481) );
  NOR2_X1 U540 ( .A1(n563), .A2(n582), .ZN(n493) );
  NAND2_X1 U541 ( .A1(n522), .A2(n493), .ZN(n484) );
  XNOR2_X1 U542 ( .A(KEYINPUT106), .B(KEYINPUT38), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(n507) );
  NOR2_X1 U544 ( .A1(n536), .A2(n507), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n485), .B(KEYINPUT40), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(G1330GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT16), .B(KEYINPUT86), .Z(n490) );
  NAND2_X1 U548 ( .A1(n586), .A2(n488), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(n492) );
  AND2_X1 U550 ( .A1(n492), .A2(n491), .ZN(n510) );
  NAND2_X1 U551 ( .A1(n493), .A2(n510), .ZN(n494) );
  XOR2_X1 U552 ( .A(KEYINPUT103), .B(n494), .Z(n502) );
  NOR2_X1 U553 ( .A1(n523), .A2(n502), .ZN(n496) );
  XNOR2_X1 U554 ( .A(KEYINPUT34), .B(KEYINPUT104), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U556 ( .A(G1GAT), .B(n497), .Z(G1324GAT) );
  NOR2_X1 U557 ( .A1(n525), .A2(n502), .ZN(n498) );
  XOR2_X1 U558 ( .A(G8GAT), .B(n498), .Z(G1325GAT) );
  NOR2_X1 U559 ( .A1(n536), .A2(n502), .ZN(n500) );
  XNOR2_X1 U560 ( .A(KEYINPUT35), .B(KEYINPUT105), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U562 ( .A(G15GAT), .B(n501), .Z(G1326GAT) );
  NOR2_X1 U563 ( .A1(n529), .A2(n502), .ZN(n503) );
  XOR2_X1 U564 ( .A(G22GAT), .B(n503), .Z(G1327GAT) );
  NOR2_X1 U565 ( .A1(n523), .A2(n507), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n504), .B(KEYINPUT39), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(n505), .ZN(G1328GAT) );
  NOR2_X1 U568 ( .A1(n525), .A2(n507), .ZN(n506) );
  XOR2_X1 U569 ( .A(G36GAT), .B(n506), .Z(G1329GAT) );
  NOR2_X1 U570 ( .A1(n529), .A2(n507), .ZN(n508) );
  XOR2_X1 U571 ( .A(G50GAT), .B(n508), .Z(G1331GAT) );
  NAND2_X1 U572 ( .A1(n553), .A2(n563), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n509), .B(KEYINPUT107), .ZN(n521) );
  NAND2_X1 U574 ( .A1(n510), .A2(n521), .ZN(n517) );
  NOR2_X1 U575 ( .A1(n523), .A2(n517), .ZN(n512) );
  XNOR2_X1 U576 ( .A(KEYINPUT42), .B(KEYINPUT108), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U578 ( .A(G57GAT), .B(n513), .Z(G1332GAT) );
  NOR2_X1 U579 ( .A1(n525), .A2(n517), .ZN(n515) );
  XNOR2_X1 U580 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(G1333GAT) );
  NOR2_X1 U582 ( .A1(n536), .A2(n517), .ZN(n516) );
  XOR2_X1 U583 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  NOR2_X1 U584 ( .A1(n529), .A2(n517), .ZN(n519) );
  XNOR2_X1 U585 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(G78GAT), .B(n520), .ZN(G1335GAT) );
  NAND2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n528) );
  NOR2_X1 U589 ( .A1(n523), .A2(n528), .ZN(n524) );
  XOR2_X1 U590 ( .A(G85GAT), .B(n524), .Z(G1336GAT) );
  NOR2_X1 U591 ( .A1(n525), .A2(n528), .ZN(n526) );
  XOR2_X1 U592 ( .A(G92GAT), .B(n526), .Z(G1337GAT) );
  NOR2_X1 U593 ( .A1(n536), .A2(n528), .ZN(n527) );
  XOR2_X1 U594 ( .A(G99GAT), .B(n527), .Z(G1338GAT) );
  NOR2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n531) );
  XNOR2_X1 U596 ( .A(KEYINPUT111), .B(KEYINPUT44), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NAND2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n550) );
  NOR2_X1 U600 ( .A1(n536), .A2(n550), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n537), .B(KEYINPUT115), .ZN(n538) );
  NOR2_X1 U602 ( .A1(n539), .A2(n538), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n576), .A2(n547), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n540), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U606 ( .A1(n547), .A2(n553), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G120GAT), .B(n543), .ZN(G1341GAT) );
  INV_X1 U609 ( .A(n547), .ZN(n544) );
  NOR2_X1 U610 ( .A1(n571), .A2(n544), .ZN(n545) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(n545), .Z(n546) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U614 ( .A1(n547), .A2(n559), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  XOR2_X1 U616 ( .A(G141GAT), .B(KEYINPUT117), .Z(n552) );
  NOR2_X1 U617 ( .A1(n573), .A2(n550), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n560), .A2(n576), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1344GAT) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n557) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n555) );
  NAND2_X1 U622 ( .A1(n560), .A2(n553), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n560), .A2(n586), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n558), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U627 ( .A(G162GAT), .B(KEYINPUT119), .Z(n562) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1347GAT) );
  NOR2_X1 U630 ( .A1(n563), .A2(n570), .ZN(n564) );
  XOR2_X1 U631 ( .A(G169GAT), .B(n564), .Z(G1348GAT) );
  NOR2_X1 U632 ( .A1(n570), .A2(n565), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n567) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n566) );
  XNOR2_X1 U635 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(G183GAT), .B(n572), .Z(G1350GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U640 ( .A(KEYINPUT123), .B(n575), .Z(n589) );
  AND2_X1 U641 ( .A1(n576), .A2(n589), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(KEYINPUT59), .B(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n584) );
  NAND2_X1 U648 ( .A1(n589), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(G204GAT), .B(n585), .ZN(G1353GAT) );
  NAND2_X1 U651 ( .A1(n589), .A2(n586), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U653 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n591) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

