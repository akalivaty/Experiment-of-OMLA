//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n549, new_n550, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n617, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1228, new_n1229;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT68), .Z(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  OAI22_X1  g035(.A1(new_n455), .A2(new_n460), .B1(new_n449), .B2(new_n457), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT69), .ZN(G319));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n466), .A2(G137), .B1(G101), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n470), .B1(new_n464), .B2(new_n465), .ZN(new_n471));
  AND2_X1   g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  AOI21_X1  g050(.A(new_n467), .B1(new_n464), .B2(new_n465), .ZN(new_n476));
  AOI22_X1  g051(.A1(G124), .A2(new_n476), .B1(new_n466), .B2(G136), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT70), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NOR3_X1   g054(.A1(KEYINPUT70), .A2(G100), .A3(G2105), .ZN(new_n480));
  OAI221_X1 g055(.A(G2104), .B1(G112), .B2(new_n467), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n477), .A2(new_n481), .ZN(G162));
  NAND2_X1  g057(.A1(G114), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G102), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2104), .ZN(new_n486));
  AND2_X1   g061(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n487));
  OAI211_X1 g062(.A(G126), .B(G2105), .C1(new_n487), .C2(new_n463), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT71), .ZN(new_n490));
  OAI211_X1 g065(.A(G138), .B(new_n467), .C1(new_n487), .C2(new_n463), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT3), .B(G2104), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n493), .A2(new_n494), .A3(G138), .A4(new_n467), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n486), .A2(new_n488), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n490), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT72), .B1(new_n501), .B2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(G543), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n502), .A2(new_n505), .B1(KEYINPUT5), .B2(new_n501), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT74), .A3(G62), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(KEYINPUT74), .B1(new_n506), .B2(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(G651), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n506), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT73), .B(G88), .ZN(new_n516));
  OAI21_X1  g091(.A(G543), .B1(new_n512), .B2(new_n513), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(G50), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n511), .A2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  OAI211_X1 g098(.A(G51), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n506), .A2(G89), .A3(new_n514), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AND2_X1   g105(.A1(new_n506), .A2(G64), .ZN(new_n531));
  AND2_X1   g106(.A1(G77), .A2(G543), .ZN(new_n532));
  OAI21_X1  g107(.A(G651), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n506), .A2(G90), .A3(new_n514), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n518), .A2(G52), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n533), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AND2_X1   g113(.A1(G68), .A2(G543), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n539), .B1(new_n506), .B2(G56), .ZN(new_n540));
  INV_X1    g115(.A(G651), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n506), .A2(G81), .A3(new_n514), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n518), .A2(G43), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT75), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(new_n550));
  XOR2_X1   g125(.A(new_n550), .B(KEYINPUT76), .Z(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(new_n502), .A2(new_n505), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n555), .A2(G65), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G78), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(new_n501), .ZN(new_n559));
  OAI21_X1  g134(.A(G651), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n506), .A2(G91), .A3(new_n514), .ZN(new_n561));
  OAI211_X1 g136(.A(G53), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT78), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT77), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT77), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n514), .A2(new_n565), .A3(G53), .A4(G543), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n566), .A3(KEYINPUT9), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  OAI211_X1 g143(.A(KEYINPUT77), .B(new_n568), .C1(new_n562), .C2(new_n563), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n560), .A2(new_n561), .A3(new_n567), .A4(new_n569), .ZN(G299));
  OAI21_X1  g145(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n506), .A2(G87), .A3(new_n514), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n518), .A2(G49), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  NAND3_X1  g149(.A1(new_n506), .A2(G86), .A3(new_n514), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n518), .A2(G48), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n506), .A2(G61), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n578), .A2(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n518), .A2(G47), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n506), .A2(new_n514), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n506), .A2(G60), .ZN(new_n588));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n541), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n555), .A2(new_n556), .ZN(new_n594));
  XNOR2_X1  g169(.A(KEYINPUT81), .B(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G651), .ZN(new_n597));
  XOR2_X1   g172(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n515), .A2(G92), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT80), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n517), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G54), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n506), .A2(G92), .A3(new_n514), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(new_n598), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n597), .A2(new_n600), .A3(new_n603), .A4(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  MUX2_X1   g182(.A(G301), .B(new_n606), .S(new_n607), .Z(G284));
  MUX2_X1   g183(.A(G301), .B(new_n606), .S(new_n607), .Z(G321));
  NOR2_X1   g184(.A1(G286), .A2(new_n607), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n567), .A2(new_n569), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n559), .B1(new_n506), .B2(G65), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n561), .B1(new_n612), .B2(new_n541), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n610), .B1(new_n614), .B2(new_n607), .ZN(G297));
  XOR2_X1   g190(.A(G297), .B(KEYINPUT82), .Z(G280));
  INV_X1    g191(.A(new_n606), .ZN(new_n617));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G860), .ZN(G148));
  NOR3_X1   g194(.A1(new_n542), .A2(new_n545), .A3(G868), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n606), .A2(G559), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n466), .A2(G2104), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g201(.A(G2100), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n476), .A2(G123), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT83), .ZN(new_n631));
  MUX2_X1   g206(.A(G99), .B(G111), .S(G2105), .Z(new_n632));
  AOI22_X1  g207(.A1(new_n466), .A2(G135), .B1(new_n632), .B2(G2104), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G2096), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n628), .A2(new_n629), .A3(new_n636), .ZN(G156));
  INV_X1    g212(.A(KEYINPUT14), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT15), .B(G2435), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2427), .ZN(new_n641));
  INV_X1    g216(.A(G2430), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n638), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n644), .A2(new_n650), .ZN(new_n652));
  AND3_X1   g227(.A1(new_n651), .A2(G14), .A3(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(G2072), .A2(G2078), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n442), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g234(.A1(new_n655), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT18), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n659), .A2(KEYINPUT84), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(KEYINPUT84), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n657), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n659), .B(KEYINPUT17), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n664), .B(new_n655), .C1(new_n657), .C2(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(new_n657), .A3(new_n654), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n661), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(new_n635), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(new_n627), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  AND2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT20), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n673), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n673), .B2(new_n679), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n686), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G229));
  XNOR2_X1  g266(.A(KEYINPUT98), .B(G28), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n692), .A2(KEYINPUT30), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT99), .ZN(new_n694));
  AOI21_X1  g269(.A(G29), .B1(new_n692), .B2(KEYINPUT30), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT31), .B(G11), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  AND2_X1   g273(.A1(KEYINPUT24), .A2(G34), .ZN(new_n699));
  NOR2_X1   g274(.A1(KEYINPUT24), .A2(G34), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT93), .Z(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G160), .B2(G29), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n696), .B(new_n697), .C1(new_n703), .C2(G2084), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n476), .A2(G129), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT94), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n468), .A2(G105), .ZN(new_n707));
  NAND3_X1  g282(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT26), .ZN(new_n709));
  AOI211_X1 g284(.A(new_n707), .B(new_n709), .C1(G141), .C2(new_n466), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(new_n698), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n698), .B2(G32), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G1996), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G2078), .ZN(new_n717));
  NAND2_X1  g292(.A1(G164), .A2(G29), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G27), .B2(G29), .ZN(new_n719));
  AOI211_X1 g294(.A(new_n704), .B(new_n716), .C1(new_n717), .C2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(G16), .A2(G19), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n546), .B2(G16), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT92), .B(G1341), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G21), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G168), .B2(new_n725), .ZN(new_n727));
  INV_X1    g302(.A(G1966), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n634), .A2(new_n698), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT97), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n698), .A2(G26), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT28), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n466), .A2(G140), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n476), .A2(G128), .ZN(new_n735));
  MUX2_X1   g310(.A(G104), .B(G116), .S(G2105), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G2104), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n733), .B1(new_n739), .B2(new_n698), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G2067), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n731), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n720), .A2(new_n724), .A3(new_n729), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n698), .A2(G35), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT100), .Z(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G162), .B2(new_n698), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT29), .Z(new_n747));
  INV_X1    g322(.A(G2090), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n725), .A2(G5), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G171), .B2(new_n725), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n747), .A2(new_n748), .B1(G1961), .B2(new_n750), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n751), .B1(G1961), .B2(new_n750), .C1(new_n717), .C2(new_n719), .ZN(new_n752));
  NOR2_X1   g327(.A1(G4), .A2(G16), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n617), .B2(G16), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1348), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n743), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n714), .A2(new_n715), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT95), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n468), .A2(G103), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT25), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n468), .A2(KEYINPUT25), .A3(G103), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n762), .A2(new_n763), .B1(new_n466), .B2(G139), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n493), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n467), .B2(new_n765), .ZN(new_n766));
  MUX2_X1   g341(.A(G33), .B(new_n766), .S(G29), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G2072), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G2084), .B2(new_n703), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n759), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT96), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n725), .A2(G20), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT23), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n614), .B2(new_n725), .ZN(new_n775));
  INV_X1    g350(.A(G1956), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n748), .B2(new_n747), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT101), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n756), .A2(new_n772), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G25), .A2(G29), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n466), .A2(G131), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT86), .Z(new_n783));
  MUX2_X1   g358(.A(G95), .B(G107), .S(G2105), .Z(new_n784));
  AOI22_X1  g359(.A1(new_n476), .A2(G119), .B1(new_n784), .B2(G2104), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n781), .B1(new_n786), .B2(G29), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT35), .B(G1991), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT87), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n787), .B(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G16), .A2(G24), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n591), .B2(G16), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G1986), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n792), .A2(G1986), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n790), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G16), .A2(G22), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G303), .B2(new_n725), .ZN(new_n798));
  INV_X1    g373(.A(G1971), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(G288), .A2(KEYINPUT88), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT88), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n571), .A2(new_n572), .A3(new_n802), .A4(new_n573), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n801), .A2(G16), .A3(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(G16), .A2(G23), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT33), .B(G1976), .Z(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n804), .A2(new_n807), .A3(new_n805), .ZN(new_n810));
  AND3_X1   g385(.A1(new_n800), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n798), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT32), .B(G1981), .ZN(new_n813));
  NOR2_X1   g388(.A1(G305), .A2(new_n725), .ZN(new_n814));
  NOR2_X1   g389(.A1(G6), .A2(G16), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n541), .B1(new_n579), .B2(new_n580), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(new_n577), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n815), .B1(new_n818), .B2(G16), .ZN(new_n819));
  INV_X1    g394(.A(new_n813), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n812), .A2(G1971), .B1(new_n816), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n811), .A2(new_n822), .A3(KEYINPUT89), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT89), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n800), .A2(new_n809), .A3(new_n810), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n819), .A2(new_n820), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n819), .A2(new_n820), .ZN(new_n827));
  OAI22_X1  g402(.A1(new_n826), .A2(new_n827), .B1(new_n798), .B2(new_n799), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n824), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT34), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n795), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT90), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n823), .A2(new_n829), .A3(KEYINPUT34), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n833), .B1(new_n832), .B2(new_n834), .ZN(new_n837));
  OAI21_X1  g412(.A(KEYINPUT36), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT36), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n832), .A2(new_n839), .A3(new_n834), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT91), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n830), .A2(new_n831), .ZN(new_n844));
  INV_X1    g419(.A(new_n795), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n844), .A2(new_n834), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT90), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(new_n835), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n848), .A2(new_n841), .A3(KEYINPUT36), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n780), .B1(new_n843), .B2(new_n849), .ZN(G311));
  INV_X1    g425(.A(new_n780), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n848), .A2(KEYINPUT36), .B1(new_n841), .B2(new_n840), .ZN(new_n852));
  AOI211_X1 g427(.A(KEYINPUT91), .B(new_n839), .C1(new_n847), .C2(new_n835), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(G150));
  NAND2_X1  g429(.A1(new_n506), .A2(G67), .ZN(new_n855));
  NAND2_X1  g430(.A1(G80), .A2(G543), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G651), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n506), .A2(G93), .A3(new_n514), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n518), .A2(G55), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(G860), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT37), .Z(new_n864));
  NOR2_X1   g439(.A1(new_n606), .A2(new_n618), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n540), .A2(new_n541), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n543), .A2(new_n544), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n866), .A2(new_n858), .A3(new_n867), .A4(new_n861), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n541), .B1(new_n855), .B2(new_n856), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n859), .A2(new_n860), .ZN(new_n870));
  OAI22_X1  g445(.A1(new_n542), .A2(new_n545), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n865), .B(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n876), .A2(KEYINPUT39), .ZN(new_n877));
  INV_X1    g452(.A(G860), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n876), .B2(KEYINPUT39), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n864), .B1(new_n877), .B2(new_n879), .ZN(G145));
  XNOR2_X1  g455(.A(new_n634), .B(KEYINPUT103), .ZN(new_n881));
  XNOR2_X1  g456(.A(G162), .B(new_n474), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n711), .B(new_n738), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n489), .B1(new_n492), .B2(new_n495), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n766), .B(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n884), .B(new_n886), .ZN(new_n887));
  MUX2_X1   g462(.A(G106), .B(G118), .S(G2105), .Z(new_n888));
  AOI22_X1  g463(.A1(new_n476), .A2(G130), .B1(new_n888), .B2(G2104), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n466), .A2(G142), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n625), .B(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n786), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n887), .A2(new_n893), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n887), .A2(KEYINPUT104), .A3(new_n893), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n883), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n895), .A2(new_n883), .ZN(new_n900));
  AOI21_X1  g475(.A(G37), .B1(new_n900), .B2(new_n894), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g478(.A(new_n621), .B(new_n872), .ZN(new_n904));
  INV_X1    g479(.A(new_n611), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n604), .B(new_n599), .ZN(new_n906));
  AOI22_X1  g481(.A1(G651), .A2(new_n596), .B1(new_n602), .B2(G54), .ZN(new_n907));
  INV_X1    g482(.A(new_n613), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n905), .A2(new_n906), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n606), .A2(G299), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n904), .A2(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT41), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT41), .B1(new_n909), .B2(new_n910), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n904), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n801), .A2(new_n803), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(G290), .ZN(new_n919));
  NAND2_X1  g494(.A1(G303), .A2(G305), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n591), .A2(new_n801), .A3(new_n803), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n511), .A2(new_n818), .A3(new_n519), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n919), .A2(new_n920), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n921), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n591), .B1(new_n801), .B2(new_n803), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n511), .A2(new_n818), .A3(new_n519), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n818), .B1(new_n511), .B2(new_n519), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n931), .A3(KEYINPUT105), .ZN(new_n932));
  INV_X1    g507(.A(new_n928), .ZN(new_n933));
  INV_X1    g508(.A(new_n931), .ZN(new_n934));
  AOI22_X1  g509(.A1(new_n925), .A2(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n917), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n935), .A2(new_n912), .A3(new_n936), .A4(new_n916), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(KEYINPUT106), .B2(KEYINPUT42), .ZN(new_n941));
  NOR2_X1   g516(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n938), .A2(new_n942), .A3(new_n939), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(G868), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n941), .A2(new_n943), .A3(KEYINPUT107), .A4(G868), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n862), .A2(new_n607), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(G295));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(G331));
  AND4_X1   g525(.A1(G63), .A2(new_n555), .A3(G651), .A4(new_n556), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(new_n525), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n533), .A2(new_n536), .A3(new_n952), .A4(new_n527), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n532), .B1(new_n506), .B2(G64), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n954), .A2(new_n541), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n534), .A2(new_n535), .ZN(new_n956));
  OAI21_X1  g531(.A(G286), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n872), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n868), .A2(new_n953), .A3(new_n957), .A4(new_n871), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n915), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n963));
  INV_X1    g538(.A(new_n960), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n871), .A2(new_n868), .B1(new_n953), .B2(new_n957), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n911), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n961), .A2(KEYINPUT110), .A3(new_n911), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n962), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n935), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n933), .A2(new_n934), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n923), .A2(new_n924), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT105), .B1(new_n928), .B2(new_n931), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n966), .A2(new_n967), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT109), .B1(new_n915), .B2(new_n961), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT41), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n911), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT41), .ZN(new_n980));
  AND4_X1   g555(.A1(KEYINPUT109), .A2(new_n961), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n975), .B(new_n976), .C1(new_n977), .C2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G37), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n971), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n976), .B1(new_n977), .B2(new_n981), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n935), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n987), .A2(new_n988), .A3(new_n983), .A4(new_n982), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(KEYINPUT44), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n984), .A2(new_n988), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n987), .A2(KEYINPUT43), .A3(new_n983), .A4(new_n982), .ZN(new_n992));
  XOR2_X1   g567(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT111), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n990), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(G397));
  AND2_X1   g574(.A1(new_n486), .A2(new_n488), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1384), .B1(new_n496), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1001), .B(KEYINPUT112), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n469), .A2(new_n473), .A3(G40), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1996), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n1005), .A2(new_n1006), .A3(new_n712), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT113), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1005), .A2(G1996), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1005), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n738), .B(G2067), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n1009), .A2(new_n712), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n786), .B(new_n789), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n1010), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1005), .A2(G1986), .A3(G290), .ZN(new_n1017));
  XNOR2_X1  g592(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1014), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n1009), .A2(KEYINPUT46), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1009), .A2(KEYINPUT46), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1010), .B1(new_n711), .B2(new_n1011), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1024), .A2(KEYINPUT47), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(KEYINPUT47), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1020), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G2067), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n739), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n786), .A2(new_n789), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(new_n1013), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(KEYINPUT126), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(new_n1005), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(KEYINPUT126), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1027), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n496), .A2(new_n1000), .ZN(new_n1037));
  INV_X1    g612(.A(G1384), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(KEYINPUT45), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n469), .A2(new_n473), .A3(G40), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n1040), .A2(KEYINPUT124), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(G2078), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1040), .A2(KEYINPUT124), .ZN(new_n1044));
  AND4_X1   g619(.A1(new_n1039), .A2(new_n1041), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1040), .B1(new_n1001), .B2(KEYINPUT45), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n486), .A2(new_n488), .A3(new_n497), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n497), .B1(new_n486), .B2(new_n488), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1384), .B1(new_n1050), .B2(new_n496), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1047), .B(new_n717), .C1(new_n1051), .C2(KEYINPUT45), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1045), .A2(new_n1046), .B1(new_n1042), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n499), .A2(KEYINPUT50), .A3(new_n1038), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(new_n885), .B2(G1384), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n1004), .ZN(new_n1058));
  INV_X1    g633(.A(G1961), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT123), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1058), .A2(KEYINPUT123), .A3(new_n1059), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1053), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1064), .A2(G171), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n499), .A2(new_n1038), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT45), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1040), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1069), .A2(new_n1043), .B1(new_n1052), .B2(new_n1042), .ZN(new_n1070));
  AOI21_X1  g645(.A(G301), .B1(new_n1070), .B2(new_n1060), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1036), .B1(new_n1065), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1064), .A2(G171), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(G301), .A3(new_n1060), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1073), .A2(KEYINPUT54), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G2084), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1057), .A2(new_n1076), .A3(new_n1004), .ZN(new_n1077));
  OAI211_X1 g652(.A(G168), .B(new_n1077), .C1(new_n1069), .C2(G1966), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(G8), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT51), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT51), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1077), .B1(new_n1069), .B2(G1966), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1082), .B2(G286), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1080), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1039), .A2(new_n1004), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT45), .B1(new_n499), .B2(new_n1038), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n799), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT114), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1040), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n748), .ZN(new_n1091));
  OAI211_X1 g666(.A(KEYINPUT114), .B(new_n799), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(G303), .A2(G8), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT55), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1094), .B(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1093), .A2(new_n1096), .A3(G8), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT49), .ZN(new_n1098));
  INV_X1    g673(.A(G1981), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n578), .B2(new_n582), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n817), .A2(new_n577), .A3(G1981), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1098), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n818), .A2(new_n1099), .ZN(new_n1103));
  OAI21_X1  g678(.A(G1981), .B1(new_n817), .B2(new_n577), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1103), .A2(KEYINPUT49), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(G8), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n1004), .B2(new_n1001), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1102), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n801), .A2(G1976), .A3(new_n803), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n1107), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT52), .ZN(new_n1111));
  INV_X1    g686(.A(G1976), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT52), .B1(G288), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1109), .A2(new_n1107), .A3(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1108), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1094), .B(KEYINPUT55), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT50), .B1(new_n499), .B2(new_n1038), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n885), .A2(new_n1055), .A3(G1384), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n748), .B(new_n1004), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1087), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G8), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1116), .A2(new_n1121), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1097), .A2(new_n1115), .A3(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1072), .A2(new_n1075), .A3(new_n1084), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1047), .B(new_n1006), .C1(new_n1051), .C2(KEYINPUT45), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1086), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1129), .A2(KEYINPUT121), .A3(new_n1006), .A4(new_n1047), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1001), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1132), .A2(new_n1040), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT58), .B(G1341), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1125), .B1(new_n1131), .B2(new_n1136), .ZN(new_n1137));
  AOI211_X1 g712(.A(KEYINPUT122), .B(new_n1135), .C1(new_n1128), .C2(new_n1130), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n546), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT59), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1141), .B(new_n546), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT119), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1144), .B1(G299), .B2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n905), .A2(new_n908), .A3(KEYINPUT119), .A4(KEYINPUT57), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT118), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n614), .B2(KEYINPUT57), .ZN(new_n1150));
  OAI211_X1 g725(.A(KEYINPUT118), .B(new_n1145), .C1(new_n611), .C2(new_n613), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1001), .A2(KEYINPUT50), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(new_n1051), .B2(KEYINPUT50), .ZN(new_n1154));
  AOI21_X1  g729(.A(G1956), .B1(new_n1154), .B2(new_n1004), .ZN(new_n1155));
  XOR2_X1   g730(.A(KEYINPUT56), .B(G2072), .Z(new_n1156));
  NOR3_X1   g731(.A1(new_n1085), .A2(new_n1086), .A3(new_n1156), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1148), .B(new_n1152), .C1(new_n1155), .C2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1157), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1004), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n776), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1151), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT118), .B1(G299), .B2(new_n1145), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1159), .B(new_n1161), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1158), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1004), .A2(new_n1001), .A3(new_n1028), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT120), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1090), .A2(G1348), .ZN(new_n1172));
  OR4_X1    g747(.A1(KEYINPUT60), .A2(new_n1171), .A3(new_n1172), .A4(new_n606), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1158), .A2(new_n1166), .A3(KEYINPUT61), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1171), .A2(new_n1172), .A3(new_n617), .ZN(new_n1175));
  OR2_X1    g750(.A1(new_n1090), .A2(G1348), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT120), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1170), .B(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n606), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT60), .B1(new_n1175), .B2(new_n1179), .ZN(new_n1180));
  AND4_X1   g755(.A1(new_n1169), .A2(new_n1173), .A3(new_n1174), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1143), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1158), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1166), .B1(new_n1183), .B2(new_n1179), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1124), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1097), .A2(new_n1071), .A3(new_n1115), .A4(new_n1122), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1081), .B1(new_n1078), .B2(G8), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1079), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1068), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1003), .B1(new_n499), .B2(new_n1038), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1004), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AOI22_X1  g767(.A1(new_n1192), .A2(new_n728), .B1(new_n1090), .B2(new_n1076), .ZN(new_n1193));
  OAI21_X1  g768(.A(KEYINPUT51), .B1(new_n1193), .B2(G168), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1188), .B1(new_n1189), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1186), .B1(new_n1187), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1197), .B1(new_n1195), .B2(new_n1187), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1084), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1196), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1115), .A2(G8), .A3(new_n1096), .A4(new_n1093), .ZN(new_n1201));
  NOR2_X1   g776(.A1(G288), .A2(G1976), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1101), .B1(new_n1108), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT115), .ZN(new_n1204));
  AND2_X1   g779(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1107), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1201), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT116), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  OAI211_X1 g784(.A(new_n1201), .B(KEYINPUT116), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1200), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1097), .A2(new_n1115), .ZN(new_n1213));
  NOR3_X1   g788(.A1(new_n1193), .A2(new_n1106), .A3(G286), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1214), .A2(KEYINPUT63), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1096), .B1(new_n1093), .B2(G8), .ZN(new_n1216));
  NOR3_X1   g791(.A1(new_n1213), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1123), .A2(KEYINPUT117), .A3(new_n1214), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1097), .A2(new_n1214), .A3(new_n1122), .A4(new_n1115), .ZN(new_n1219));
  INV_X1    g794(.A(KEYINPUT117), .ZN(new_n1220));
  AOI21_X1  g795(.A(KEYINPUT63), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1217), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1222));
  NOR3_X1   g797(.A1(new_n1185), .A2(new_n1212), .A3(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g798(.A(new_n591), .B(G1986), .ZN(new_n1224));
  OAI211_X1 g799(.A(new_n1014), .B(new_n1016), .C1(new_n1005), .C2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g800(.A(new_n1035), .B1(new_n1223), .B2(new_n1225), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g801(.A1(G227), .A2(new_n461), .A3(G401), .ZN(new_n1228));
  AND3_X1   g802(.A1(new_n690), .A2(new_n902), .A3(new_n1228), .ZN(new_n1229));
  NAND3_X1  g803(.A1(new_n1229), .A2(new_n991), .A3(new_n992), .ZN(G225));
  INV_X1    g804(.A(G225), .ZN(G308));
endmodule


