//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G131), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n192), .B1(new_n188), .B2(G137), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n187), .A2(new_n189), .A3(new_n191), .A4(new_n193), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n193), .A2(new_n189), .A3(new_n191), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n194), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT68), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT67), .B(G128), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT1), .B1(new_n200), .B2(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT66), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n203), .B(KEYINPUT1), .C1(new_n200), .C2(G146), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n199), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n200), .A2(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n198), .B1(new_n205), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n199), .ZN(new_n212));
  INV_X1    g026(.A(new_n204), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n203), .B1(new_n207), .B2(KEYINPUT1), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT68), .A3(new_n209), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT79), .B(G101), .ZN(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT3), .B1(new_n219), .B2(G107), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(G107), .ZN(new_n221));
  OR2_X1    g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT77), .A2(G107), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT77), .A2(G107), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n219), .A2(KEYINPUT3), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT78), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT77), .ZN(new_n228));
  INV_X1    g042(.A(G107), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT77), .A2(G107), .ZN(new_n231));
  AND4_X1   g045(.A1(KEYINPUT78), .A2(new_n226), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n218), .B(new_n222), .C1(new_n227), .C2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n225), .A2(G104), .ZN(new_n234));
  OAI21_X1  g048(.A(G101), .B1(new_n234), .B2(new_n221), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G128), .ZN(new_n237));
  OR3_X1    g051(.A1(new_n209), .A2(KEYINPUT1), .A3(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n217), .A2(new_n236), .A3(KEYINPUT82), .A4(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n237), .B1(new_n207), .B2(KEYINPUT1), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n238), .B1(new_n240), .B2(new_n210), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(new_n233), .A3(new_n235), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n238), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(new_n211), .B2(new_n216), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT82), .B1(new_n245), .B2(new_n236), .ZN(new_n246));
  OAI211_X1 g060(.A(KEYINPUT12), .B(new_n197), .C1(new_n243), .C2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT83), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT82), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT68), .B1(new_n215), .B2(new_n209), .ZN(new_n250));
  NOR3_X1   g064(.A1(new_n205), .A2(new_n198), .A3(new_n210), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n238), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n236), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(new_n242), .A3(new_n239), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT83), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT12), .A4(new_n197), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n197), .B1(new_n243), .B2(new_n246), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT12), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n248), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n233), .A2(KEYINPUT10), .A3(new_n235), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n252), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  AND2_X1   g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n209), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n209), .B2(new_n265), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n222), .B1(new_n227), .B2(new_n232), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(G101), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n233), .A2(KEYINPUT4), .ZN(new_n271));
  INV_X1    g085(.A(G101), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n226), .A2(new_n230), .A3(new_n231), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT78), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n225), .A2(KEYINPUT78), .A3(new_n226), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n272), .B1(new_n277), .B2(new_n222), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n267), .B(new_n270), .C1(new_n271), .C2(new_n278), .ZN(new_n279));
  XOR2_X1   g093(.A(KEYINPUT81), .B(KEYINPUT10), .Z(new_n280));
  NAND2_X1  g094(.A1(new_n242), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n263), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  OR2_X1    g096(.A1(new_n282), .A2(new_n197), .ZN(new_n283));
  XNOR2_X1  g097(.A(G110), .B(G140), .ZN(new_n284));
  INV_X1    g098(.A(G953), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n285), .A2(G227), .ZN(new_n286));
  XOR2_X1   g100(.A(new_n284), .B(new_n286), .Z(new_n287));
  AND2_X1   g101(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n261), .A2(new_n288), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n282), .A2(KEYINPUT84), .A3(new_n197), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT84), .B1(new_n282), .B2(new_n197), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n283), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n287), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G469), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT85), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n289), .B2(new_n294), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT85), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n301), .A3(new_n296), .ZN(new_n302));
  OR2_X1    g116(.A1(new_n290), .A2(new_n291), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n303), .A2(new_n288), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n287), .B1(new_n261), .B2(new_n283), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n297), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n299), .A2(new_n302), .B1(G469), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT9), .B(G234), .ZN(new_n308));
  OAI21_X1  g122(.A(G221), .B1(new_n308), .B2(G902), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n309), .B(KEYINPUT76), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT86), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(G214), .B1(G237), .B2(G902), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT87), .ZN(new_n313));
  OAI21_X1  g127(.A(G210), .B1(G237), .B2(G902), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G119), .ZN(new_n316));
  OR2_X1    g130(.A1(new_n316), .A2(G116), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(G116), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT2), .B(G113), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g135(.A1(new_n318), .A2(KEYINPUT5), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n322), .A2(G113), .ZN(new_n323));
  INV_X1    g137(.A(new_n319), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT5), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT88), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n323), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(KEYINPUT88), .B1(new_n324), .B2(KEYINPUT5), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n321), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n253), .ZN(new_n330));
  XNOR2_X1  g144(.A(G110), .B(G122), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT8), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n325), .A2(new_n323), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n321), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n330), .B(new_n332), .C1(new_n253), .C2(new_n334), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n334), .A2(new_n236), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n319), .A2(new_n320), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n321), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n338), .B(new_n270), .C1(new_n271), .C2(new_n278), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n339), .A3(new_n331), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT73), .B(G125), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n267), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(new_n245), .B2(new_n341), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n285), .A2(G224), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n344), .A2(KEYINPUT7), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n335), .B(new_n340), .C1(new_n343), .C2(new_n345), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n343), .A2(KEYINPUT7), .A3(new_n344), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n297), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT89), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n336), .A2(new_n339), .ZN(new_n352));
  INV_X1    g166(.A(new_n331), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(KEYINPUT6), .A3(new_n340), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n343), .B(new_n344), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT6), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n352), .A2(new_n357), .A3(new_n353), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(new_n348), .B2(new_n349), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n315), .B1(new_n351), .B2(new_n360), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n348), .A2(new_n349), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n362), .A2(new_n314), .A3(new_n350), .A4(new_n359), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n313), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(G475), .A2(G902), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G113), .B(G122), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(new_n219), .ZN(new_n369));
  INV_X1    g183(.A(G237), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(new_n285), .A3(G214), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT90), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT91), .B1(new_n373), .B2(G143), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n372), .B(new_n374), .C1(KEYINPUT91), .C2(G143), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n371), .B(KEYINPUT91), .C1(new_n373), .C2(G143), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT18), .A2(G131), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(G125), .A2(G140), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(new_n341), .B2(G140), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G146), .ZN(new_n382));
  XNOR2_X1  g196(.A(G125), .B(G140), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n206), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT16), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n381), .A2(new_n388), .ZN(new_n389));
  XOR2_X1   g203(.A(KEYINPUT73), .B(G125), .Z(new_n390));
  NOR3_X1   g204(.A1(new_n390), .A2(KEYINPUT16), .A3(G140), .ZN(new_n391));
  OR3_X1    g205(.A1(new_n389), .A2(new_n206), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n187), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n375), .A2(new_n393), .A3(new_n376), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT17), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n206), .B1(new_n389), .B2(new_n391), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n392), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(KEYINPUT93), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n392), .A2(new_n396), .A3(KEYINPUT93), .A4(new_n397), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n377), .A2(new_n187), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n395), .A3(new_n394), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n369), .B(new_n387), .C1(new_n399), .C2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n369), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT92), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n383), .A2(KEYINPUT19), .ZN(new_n407));
  INV_X1    g221(.A(new_n380), .ZN(new_n408));
  INV_X1    g222(.A(G140), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n408), .B1(new_n390), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n407), .B1(new_n410), .B2(KEYINPUT19), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n406), .B1(new_n411), .B2(G146), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n401), .A2(new_n394), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n392), .A3(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n411), .A2(G146), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n414), .B1(KEYINPUT92), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n405), .B1(new_n416), .B2(new_n386), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n367), .B1(new_n404), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT20), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n404), .A2(new_n417), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n366), .B(KEYINPUT94), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n387), .B1(new_n399), .B2(new_n403), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n405), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT95), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(new_n404), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(KEYINPUT95), .A3(new_n405), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n297), .A3(new_n428), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n420), .A2(new_n423), .B1(new_n429), .B2(G475), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT97), .ZN(new_n431));
  XNOR2_X1  g245(.A(G116), .B(G122), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n225), .B(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT96), .ZN(new_n434));
  OR2_X1    g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n237), .A2(G143), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n199), .B2(G143), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT13), .ZN(new_n438));
  INV_X1    g252(.A(new_n436), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n438), .B(G134), .C1(KEYINPUT13), .C2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n437), .A2(new_n188), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n433), .A2(new_n434), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n435), .A2(new_n440), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n225), .A2(new_n432), .ZN(new_n444));
  INV_X1    g258(.A(G122), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT14), .B1(new_n445), .B2(G116), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n445), .A2(G116), .ZN(new_n447));
  MUX2_X1   g261(.A(new_n446), .B(KEYINPUT14), .S(new_n447), .Z(new_n448));
  INV_X1    g262(.A(new_n441), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n437), .A2(new_n188), .ZN(new_n450));
  OAI221_X1 g264(.A(new_n444), .B1(new_n448), .B2(new_n229), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G217), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n308), .A2(new_n452), .A3(G953), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n443), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n453), .B1(new_n443), .B2(new_n451), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n297), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n431), .B1(new_n456), .B2(KEYINPUT98), .ZN(new_n457));
  INV_X1    g271(.A(G478), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(KEYINPUT15), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n459), .B1(new_n456), .B2(new_n431), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n457), .B(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT99), .B(G952), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(G953), .ZN(new_n464));
  NAND2_X1  g278(.A1(G234), .A2(G237), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n465), .A2(G902), .A3(G953), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(G898), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n470), .B(KEYINPUT100), .Z(new_n471));
  NAND3_X1  g285(.A1(new_n430), .A2(new_n462), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n365), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n306), .A2(G469), .ZN(new_n474));
  AND4_X1   g288(.A1(new_n301), .A2(new_n295), .A3(new_n296), .A4(new_n297), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n301), .B1(new_n300), .B2(new_n296), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT86), .ZN(new_n478));
  INV_X1    g292(.A(new_n310), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n311), .A2(new_n473), .A3(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(G472), .A2(G902), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n197), .A2(new_n267), .ZN(new_n483));
  INV_X1    g297(.A(new_n189), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n188), .A2(G137), .ZN(new_n485));
  OAI21_X1  g299(.A(G131), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n194), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n483), .B1(new_n245), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT30), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT69), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n487), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n252), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT69), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT30), .A4(new_n483), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n487), .B(KEYINPUT65), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n483), .B1(new_n245), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n489), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n490), .A2(new_n494), .A3(new_n497), .A4(new_n338), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n370), .A2(new_n285), .A3(G210), .ZN(new_n499));
  XOR2_X1   g313(.A(new_n499), .B(KEYINPUT27), .Z(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT26), .B(G101), .ZN(new_n501));
  XOR2_X1   g315(.A(new_n500), .B(new_n501), .Z(new_n502));
  INV_X1    g316(.A(new_n338), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n503), .B(new_n483), .C1(new_n245), .C2(new_n487), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n498), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n483), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT65), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n487), .B(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n506), .B1(new_n252), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n504), .B1(new_n509), .B2(new_n503), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT28), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n488), .A2(KEYINPUT70), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT70), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n513), .B(new_n483), .C1(new_n245), .C2(new_n487), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n338), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n511), .B1(new_n515), .B2(KEYINPUT28), .ZN(new_n516));
  INV_X1    g330(.A(new_n502), .ZN(new_n517));
  AOI22_X1  g331(.A1(KEYINPUT31), .A2(new_n505), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT31), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n498), .A2(new_n519), .A3(new_n502), .A4(new_n504), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT71), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n505), .A2(KEYINPUT31), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n516), .A2(new_n517), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT71), .A4(new_n520), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n482), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT32), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g342(.A(KEYINPUT32), .B(new_n482), .C1(new_n521), .C2(new_n525), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n488), .B(new_n503), .ZN(new_n530));
  MUX2_X1   g344(.A(new_n515), .B(new_n530), .S(KEYINPUT28), .Z(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(KEYINPUT29), .A3(new_n502), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n498), .A2(new_n504), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(new_n502), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT29), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(new_n516), .B2(new_n517), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n532), .B(new_n297), .C1(new_n535), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G472), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n528), .A2(new_n529), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n392), .A2(new_n384), .ZN(new_n541));
  XOR2_X1   g355(.A(KEYINPUT72), .B(KEYINPUT23), .Z(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n316), .B2(G128), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n199), .A2(KEYINPUT23), .A3(G119), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n543), .B(new_n544), .C1(G119), .C2(new_n237), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(G110), .ZN(new_n546));
  OR2_X1    g360(.A1(new_n546), .A2(KEYINPUT74), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n237), .A2(G119), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n199), .B2(G119), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT24), .B(G110), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n546), .B2(KEYINPUT74), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n541), .B1(new_n547), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n392), .A2(new_n397), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n545), .A2(G110), .B1(new_n549), .B2(new_n551), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n285), .A2(G221), .A3(G234), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT75), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT22), .B(G137), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n555), .A2(new_n558), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n558), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n562), .B1(new_n554), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT25), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n568), .A3(new_n297), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n452), .B1(G234), .B2(new_n297), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n568), .B1(new_n567), .B2(new_n297), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n570), .A2(G902), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n573), .B1(new_n567), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n540), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n481), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT102), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n218), .B(KEYINPUT101), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(G3));
  INV_X1    g394(.A(G472), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n522), .A2(new_n523), .A3(new_n520), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT71), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(G902), .B1(new_n584), .B2(new_n524), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n575), .B(new_n526), .C1(new_n581), .C2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n587), .A2(new_n311), .A3(new_n480), .ZN(new_n588));
  INV_X1    g402(.A(new_n312), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(new_n361), .B2(new_n363), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n471), .ZN(new_n591));
  INV_X1    g405(.A(new_n430), .ZN(new_n592));
  OR3_X1    g406(.A1(new_n454), .A2(new_n455), .A3(KEYINPUT33), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT33), .B1(new_n454), .B2(new_n455), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(G478), .B1(new_n596), .B2(G902), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n456), .A2(G478), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n592), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n591), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n588), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT34), .B(G104), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G6));
  INV_X1    g419(.A(new_n418), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT103), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT20), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT103), .B1(new_n418), .B2(new_n419), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n421), .A2(new_n419), .A3(new_n366), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n429), .A2(G475), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n611), .A2(new_n612), .A3(new_n461), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(new_n590), .A3(new_n471), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT104), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT104), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n613), .A2(new_n590), .A3(new_n616), .A4(new_n471), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n588), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT35), .B(G107), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G9));
  NAND2_X1  g435(.A1(new_n555), .A2(new_n558), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n563), .A2(KEYINPUT36), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n574), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n625), .B1(new_n571), .B2(new_n572), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n526), .B(new_n626), .C1(new_n585), .C2(new_n581), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n311), .A2(new_n628), .A3(new_n473), .A4(new_n480), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT37), .B(G110), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G12));
  AND3_X1   g445(.A1(new_n311), .A2(new_n480), .A3(new_n590), .ZN(new_n632));
  INV_X1    g446(.A(G900), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n467), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n466), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n613), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n540), .A2(new_n637), .A3(new_n626), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n632), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n311), .A2(new_n480), .A3(new_n590), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT105), .B1(new_n642), .B2(new_n638), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G128), .ZN(G30));
  XOR2_X1   g459(.A(new_n635), .B(KEYINPUT39), .Z(new_n646));
  NAND3_X1  g460(.A1(new_n311), .A2(new_n480), .A3(new_n646), .ZN(new_n647));
  OR2_X1    g461(.A1(new_n647), .A2(KEYINPUT40), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(KEYINPUT40), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n505), .B1(new_n502), .B2(new_n530), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n650), .A2(new_n297), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n528), .B(new_n529), .C1(new_n581), .C2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n361), .A2(new_n363), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n653), .B(KEYINPUT38), .Z(new_n654));
  NOR2_X1   g468(.A1(new_n430), .A2(new_n462), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR4_X1   g470(.A1(new_n654), .A2(new_n589), .A3(new_n626), .A4(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n648), .A2(new_n649), .A3(new_n652), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT106), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G143), .ZN(G45));
  NAND3_X1  g474(.A1(new_n592), .A2(new_n600), .A3(new_n636), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n540), .A2(new_n626), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n642), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n206), .ZN(G48));
  OR2_X1    g479(.A1(new_n300), .A2(new_n296), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n479), .B(new_n666), .C1(new_n475), .C2(new_n476), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n299), .A2(new_n302), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n670), .A2(KEYINPUT107), .A3(new_n479), .A4(new_n666), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT108), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n540), .A2(new_n575), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n669), .A2(KEYINPUT108), .A3(new_n671), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n674), .A2(new_n602), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT41), .B(G113), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G15));
  NAND4_X1  g493(.A1(new_n674), .A2(new_n618), .A3(new_n675), .A4(new_n676), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G116), .ZN(G18));
  NAND2_X1  g495(.A1(new_n540), .A2(new_n626), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n472), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n669), .A2(new_n590), .A3(new_n671), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G119), .ZN(G21));
  OR2_X1    g500(.A1(new_n585), .A2(new_n581), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n522), .B(new_n520), .C1(new_n531), .C2(new_n502), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n482), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n687), .A2(new_n575), .A3(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n655), .A2(new_n590), .A3(new_n471), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n674), .A2(new_n676), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT109), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n674), .A2(new_n692), .A3(new_n695), .A4(new_n676), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G122), .ZN(G24));
  OAI211_X1 g512(.A(new_n626), .B(new_n689), .C1(new_n585), .C2(new_n581), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n661), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(new_n590), .A3(new_n669), .A4(new_n671), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G125), .ZN(G27));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n361), .A2(new_n363), .A3(new_n312), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n307), .A2(new_n310), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n675), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n703), .B1(new_n706), .B2(new_n661), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n526), .A2(new_n709), .A3(new_n527), .ZN(new_n710));
  INV_X1    g524(.A(new_n482), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n584), .B2(new_n524), .ZN(new_n712));
  AOI21_X1  g526(.A(KEYINPUT110), .B1(new_n712), .B2(KEYINPUT32), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(KEYINPUT32), .ZN(new_n714));
  OAI211_X1 g528(.A(KEYINPUT111), .B(new_n710), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n539), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n529), .A2(new_n709), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n528), .ZN(new_n718));
  AOI21_X1  g532(.A(KEYINPUT111), .B1(new_n718), .B2(new_n710), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n575), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(KEYINPUT112), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n722), .B(new_n575), .C1(new_n716), .C2(new_n719), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n704), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n477), .A2(new_n725), .A3(new_n479), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n726), .A2(new_n703), .A3(new_n661), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n708), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n196), .ZN(G33));
  NAND4_X1  g543(.A1(new_n705), .A2(new_n540), .A3(new_n575), .A4(new_n637), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G134), .ZN(G36));
  NAND2_X1  g545(.A1(new_n600), .A2(new_n430), .ZN(new_n732));
  XOR2_X1   g546(.A(new_n732), .B(KEYINPUT43), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT113), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n687), .A2(new_n526), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n734), .A2(new_n735), .A3(new_n626), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n704), .B1(new_n736), .B2(KEYINPUT44), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n737), .B1(KEYINPUT44), .B2(new_n736), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n304), .A2(new_n305), .ZN(new_n739));
  XOR2_X1   g553(.A(new_n739), .B(KEYINPUT45), .Z(new_n740));
  OAI21_X1  g554(.A(G469), .B1(new_n740), .B2(G902), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n741), .A2(KEYINPUT46), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(KEYINPUT46), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n670), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n479), .A3(new_n646), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n738), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n190), .ZN(G39));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n479), .ZN(new_n748));
  XOR2_X1   g562(.A(new_n748), .B(KEYINPUT47), .Z(new_n749));
  NOR4_X1   g563(.A1(new_n540), .A2(new_n704), .A3(new_n575), .A4(new_n661), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n409), .ZN(G42));
  INV_X1    g566(.A(new_n313), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n575), .A2(new_n479), .A3(new_n753), .ZN(new_n754));
  OR3_X1    g568(.A1(new_n754), .A2(KEYINPUT114), .A3(new_n732), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT114), .B1(new_n754), .B2(new_n732), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n654), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n670), .A2(new_n666), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n758), .A2(KEYINPUT49), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(KEYINPUT49), .ZN(new_n760));
  OR4_X1    g574(.A1(new_n652), .A2(new_n757), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n466), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n733), .A2(new_n762), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n763), .A2(new_n690), .ZN(new_n764));
  INV_X1    g578(.A(new_n684), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n464), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n601), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n669), .A2(new_n671), .A3(new_n725), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n575), .A2(new_n762), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n768), .A2(new_n652), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n766), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n654), .A2(new_n589), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n764), .A2(new_n672), .A3(new_n772), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT50), .Z(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n763), .A2(new_n768), .ZN(new_n776));
  INV_X1    g590(.A(new_n699), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n592), .A2(new_n600), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n776), .A2(new_n777), .B1(new_n770), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n775), .A2(KEYINPUT51), .A3(new_n779), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n764), .A2(new_n704), .ZN(new_n781));
  INV_X1    g595(.A(new_n749), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n758), .A2(new_n479), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n781), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n771), .B1(new_n780), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT48), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n724), .A2(new_n776), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n782), .A2(KEYINPUT119), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT119), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n783), .B1(new_n749), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n781), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n774), .A2(KEYINPUT120), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n779), .ZN(new_n795));
  AOI211_X1 g609(.A(new_n793), .B(new_n795), .C1(KEYINPUT120), .C2(new_n774), .ZN(new_n796));
  OAI221_X1 g610(.A(new_n789), .B1(new_n787), .B2(new_n788), .C1(new_n796), .C2(KEYINPUT51), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n680), .A2(new_n677), .A3(new_n685), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n626), .A2(new_n361), .A3(new_n363), .A4(new_n312), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n461), .A2(new_n635), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n612), .A3(new_n611), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n800), .A2(new_n611), .A3(KEYINPUT115), .A4(new_n612), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n799), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(new_n311), .A3(new_n540), .A4(new_n480), .ZN(new_n806));
  NOR4_X1   g620(.A1(new_n726), .A2(new_n699), .A3(KEYINPUT116), .A4(new_n661), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n705), .B2(new_n700), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n730), .B(new_n806), .C1(new_n807), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n420), .A2(new_n423), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n612), .A3(new_n461), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n812), .B1(new_n430), .B2(new_n599), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n813), .A2(new_n364), .A3(new_n471), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n587), .A2(new_n814), .A3(new_n311), .A4(new_n480), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n815), .B(new_n629), .C1(new_n576), .C2(new_n481), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n810), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n798), .A2(new_n817), .A3(new_n697), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n728), .ZN(new_n819));
  INV_X1    g633(.A(new_n663), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n632), .A2(new_n820), .B1(new_n684), .B2(new_n700), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n655), .A2(new_n590), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n822), .A2(new_n626), .A3(new_n635), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n823), .A2(new_n479), .A3(new_n477), .A4(new_n652), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n640), .B1(new_n632), .B2(new_n639), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n642), .A2(new_n638), .A3(KEYINPUT105), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n821), .B(new_n824), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n701), .B1(new_n642), .B2(new_n663), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n641), .B2(new_n643), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(KEYINPUT52), .A3(new_n824), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n819), .A2(KEYINPUT53), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT53), .B1(new_n819), .B2(new_n833), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n834), .B1(new_n835), .B2(KEYINPUT117), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n837));
  AOI211_X1 g651(.A(new_n837), .B(KEYINPUT53), .C1(new_n819), .C2(new_n833), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT54), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n798), .A2(new_n817), .A3(new_n697), .ZN(new_n841));
  INV_X1    g655(.A(new_n723), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n710), .B1(new_n713), .B2(new_n714), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT111), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n539), .A3(new_n715), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n722), .B1(new_n846), .B2(new_n575), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n727), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n707), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n841), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n829), .A2(new_n832), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n840), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(new_n853), .A3(new_n834), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT118), .B1(new_n839), .B2(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n839), .A2(KEYINPUT118), .A3(new_n854), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n797), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(G952), .A2(G953), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n761), .B1(new_n857), .B2(new_n858), .ZN(G75));
  NAND2_X1  g673(.A1(new_n852), .A2(new_n834), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(G902), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT56), .B1(new_n862), .B2(G210), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n355), .A2(new_n358), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(new_n356), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n865), .B(KEYINPUT55), .Z(new_n866));
  OAI22_X1  g680(.A1(new_n863), .A2(new_n866), .B1(G952), .B2(new_n285), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n863), .B2(new_n866), .ZN(G51));
  NOR2_X1   g682(.A1(new_n285), .A2(G952), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n860), .A2(KEYINPUT54), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n854), .ZN(new_n871));
  NAND2_X1  g685(.A1(G469), .A2(G902), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT57), .Z(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n295), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n862), .A2(G469), .A3(new_n740), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n869), .B1(new_n875), .B2(new_n876), .ZN(G54));
  AND3_X1   g691(.A1(new_n862), .A2(KEYINPUT58), .A3(G475), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n878), .A2(new_n421), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n421), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n879), .A2(new_n880), .A3(new_n869), .ZN(G60));
  NAND2_X1  g695(.A1(G478), .A2(G902), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT59), .Z(new_n883));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n884));
  AND4_X1   g698(.A1(KEYINPUT53), .A2(new_n833), .A3(new_n849), .A4(new_n841), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n885), .B1(new_n837), .B2(new_n852), .ZN(new_n886));
  INV_X1    g700(.A(new_n838), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n853), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n854), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n884), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n839), .A2(KEYINPUT118), .A3(new_n854), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n883), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT121), .B1(new_n892), .B2(new_n595), .ZN(new_n893));
  INV_X1    g707(.A(new_n883), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(new_n856), .B2(new_n855), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n896), .A3(new_n596), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n596), .A2(new_n883), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n869), .B1(new_n871), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n893), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT122), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n893), .A2(new_n897), .A3(new_n902), .A4(new_n899), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(G63));
  NAND2_X1  g718(.A1(G217), .A2(G902), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT60), .Z(new_n906));
  AND3_X1   g720(.A1(new_n860), .A2(new_n624), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n860), .A2(new_n906), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n567), .B(KEYINPUT123), .Z(new_n909));
  AOI211_X1 g723(.A(new_n869), .B(new_n907), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT61), .ZN(G66));
  NAND2_X1  g725(.A1(new_n798), .A2(new_n697), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n912), .A2(new_n816), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(G224), .A2(G953), .ZN(new_n915));
  OAI22_X1  g729(.A1(new_n914), .A2(G953), .B1(new_n468), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(G898), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n864), .B1(new_n917), .B2(G953), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n916), .B(new_n918), .ZN(G69));
  NAND3_X1  g733(.A1(new_n490), .A2(new_n494), .A3(new_n497), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(new_n411), .ZN(new_n921));
  INV_X1    g735(.A(new_n746), .ZN(new_n922));
  INV_X1    g736(.A(new_n751), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n922), .A2(new_n923), .A3(new_n730), .A4(new_n831), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n745), .A2(new_n822), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n728), .B(new_n924), .C1(new_n724), .C2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n926), .A2(G953), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n285), .A2(G900), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT126), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n921), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n921), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n813), .B(KEYINPUT125), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n675), .A2(new_n725), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n922), .B1(new_n647), .B2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n659), .A2(KEYINPUT124), .A3(KEYINPUT62), .A4(new_n831), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n659), .A2(new_n831), .ZN(new_n936));
  XOR2_X1   g750(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI211_X1 g752(.A(new_n751), .B(new_n934), .C1(new_n935), .C2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n931), .B1(new_n939), .B2(G953), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n930), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n285), .B1(G227), .B2(G900), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n942), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n930), .A2(new_n940), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n945), .ZN(G72));
  NOR2_X1   g760(.A1(new_n534), .A2(new_n517), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n533), .A2(new_n502), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(G472), .A2(G902), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT63), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n869), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  AOI22_X1  g766(.A1(new_n926), .A2(new_n948), .B1(new_n939), .B2(new_n947), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n952), .B1(new_n953), .B2(new_n914), .ZN(new_n954));
  AOI211_X1 g768(.A(new_n951), .B(new_n949), .C1(new_n886), .C2(new_n887), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT127), .Z(new_n956));
  NOR2_X1   g770(.A1(new_n954), .A2(new_n956), .ZN(G57));
endmodule


