//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(G101), .ZN(new_n191));
  INV_X1    g005(.A(G237), .ZN(new_n192));
  INV_X1    g006(.A(G953), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G210), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n191), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT11), .A3(G134), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G137), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n201), .B1(new_n198), .B2(G137), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n196), .A2(G134), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(new_n201), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n200), .A2(KEYINPUT68), .A3(new_n203), .A4(new_n206), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n207), .A2(G131), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n200), .A2(new_n203), .A3(new_n206), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(G131), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n200), .A2(new_n212), .A3(new_n203), .A4(new_n206), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n205), .B1(new_n204), .B2(new_n201), .ZN(new_n216));
  AOI211_X1 g030(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n196), .C2(G134), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n218), .A2(KEYINPUT67), .A3(new_n212), .A4(new_n200), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n208), .A2(new_n211), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G146), .ZN(new_n224));
  INV_X1    g038(.A(G143), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(G146), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  OR2_X1    g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n222), .A2(new_n224), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G143), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n221), .A2(G143), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n230), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n232), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT71), .B1(new_n220), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n215), .A2(new_n219), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n211), .A2(G131), .A3(new_n207), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n244));
  INV_X1    g058(.A(new_n239), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n240), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G116), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(G119), .ZN(new_n249));
  OR2_X1    g063(.A1(KEYINPUT70), .A2(G116), .ZN(new_n250));
  NAND2_X1  g064(.A1(KEYINPUT70), .A2(G116), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n249), .B1(new_n252), .B2(G119), .ZN(new_n253));
  XOR2_X1   g067(.A(KEYINPUT2), .B(G113), .Z(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n235), .B1(new_n233), .B2(G143), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT1), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(G128), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n261));
  INV_X1    g075(.A(new_n229), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OR2_X1    g077(.A1(new_n199), .A2(KEYINPUT69), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n199), .A2(KEYINPUT69), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(new_n204), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G131), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n241), .A2(new_n263), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n247), .A2(new_n256), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n243), .A2(new_n245), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT30), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n270), .A2(new_n271), .A3(new_n268), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n244), .B1(new_n243), .B2(new_n245), .ZN(new_n273));
  AOI211_X1 g087(.A(KEYINPUT71), .B(new_n239), .C1(new_n241), .C2(new_n242), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n268), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n272), .B1(new_n275), .B2(KEYINPUT30), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n195), .B(new_n269), .C1(new_n276), .C2(new_n256), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT31), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n268), .ZN(new_n280));
  AOI211_X1 g094(.A(new_n255), .B(new_n280), .C1(new_n240), .C2(new_n246), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n270), .A2(new_n271), .A3(new_n268), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n280), .B1(new_n240), .B2(new_n246), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n282), .B1(new_n283), .B2(new_n271), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n281), .B1(new_n284), .B2(new_n255), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(KEYINPUT31), .A3(new_n195), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n279), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n270), .A2(new_n268), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n255), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT28), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n290), .B1(new_n288), .B2(new_n255), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n289), .B(new_n291), .C1(new_n269), .C2(new_n290), .ZN(new_n292));
  INV_X1    g106(.A(new_n195), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n189), .B1(new_n287), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n187), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n294), .B1(new_n279), .B2(new_n286), .ZN(new_n299));
  OAI211_X1 g113(.A(KEYINPUT72), .B(KEYINPUT32), .C1(new_n299), .C2(new_n189), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G472), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n256), .B1(new_n247), .B2(new_n268), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT28), .B1(new_n303), .B2(new_n281), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n291), .A2(KEYINPUT74), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g120(.A(KEYINPUT74), .B(KEYINPUT28), .C1(new_n303), .C2(new_n281), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n306), .A2(KEYINPUT29), .A3(new_n195), .A4(new_n307), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT75), .B(G902), .Z(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT73), .B1(new_n285), .B2(new_n195), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n269), .B1(new_n276), .B2(new_n256), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT73), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(new_n293), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n292), .A2(new_n293), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n312), .A2(new_n315), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n302), .B1(new_n311), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n301), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  INV_X1    g136(.A(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(G125), .A2(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT16), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n322), .A2(KEYINPUT16), .A3(G140), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(G146), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n233), .A2(new_n326), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n260), .A2(G119), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n260), .A2(G119), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT23), .ZN(new_n334));
  OAI211_X1 g148(.A(KEYINPUT77), .B(new_n332), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n334), .A2(KEYINPUT77), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n335), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(G110), .ZN(new_n338));
  XOR2_X1   g152(.A(KEYINPUT24), .B(G110), .Z(new_n339));
  XNOR2_X1  g153(.A(new_n332), .B(KEYINPUT76), .ZN(new_n340));
  INV_X1    g154(.A(new_n333), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n330), .B(new_n331), .C1(new_n338), .C2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT16), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n344), .B1(new_n324), .B2(new_n325), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n221), .B1(new_n345), .B2(new_n328), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n330), .A2(new_n346), .A3(KEYINPUT78), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n340), .A2(new_n341), .A3(new_n339), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n337), .A2(G110), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n327), .A2(new_n350), .A3(G146), .A4(new_n329), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n347), .A2(new_n348), .A3(new_n349), .A4(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n343), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n193), .A2(G221), .A3(G234), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(KEYINPUT22), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(G137), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n343), .A2(new_n352), .A3(new_n356), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OR3_X1    g174(.A1(new_n360), .A2(KEYINPUT25), .A3(new_n309), .ZN(new_n361));
  INV_X1    g175(.A(G217), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(new_n310), .B2(G234), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT25), .B1(new_n360), .B2(new_n309), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n360), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n363), .A2(G902), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n347), .A2(new_n351), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n192), .A2(new_n193), .A3(G214), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n225), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n192), .A2(new_n193), .A3(G143), .A4(G214), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n212), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(KEYINPUT17), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n375), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT17), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n372), .A2(new_n212), .A3(new_n373), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n370), .A2(new_n376), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(KEYINPUT18), .A2(G131), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT87), .B1(new_n374), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n331), .B1(new_n221), .B2(new_n326), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n374), .A2(new_n383), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT87), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n372), .A2(new_n387), .A3(new_n373), .A4(new_n382), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n384), .A2(new_n385), .A3(new_n386), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n381), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(G113), .B(G122), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n381), .A2(new_n393), .A3(new_n389), .ZN(new_n396));
  AOI21_X1  g210(.A(G902), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G475), .ZN(new_n398));
  OR2_X1    g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G902), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(KEYINPUT88), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT19), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n326), .B(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT64), .B(G146), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n330), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n377), .A2(new_n379), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n389), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n394), .ZN(new_n409));
  AOI211_X1 g223(.A(KEYINPUT20), .B(new_n402), .C1(new_n396), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT89), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n402), .B1(new_n396), .B2(new_n409), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT20), .ZN(new_n413));
  OR2_X1    g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n410), .A2(KEYINPUT89), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n399), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT90), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(KEYINPUT90), .B(new_n399), .C1(new_n415), .C2(new_n416), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT96), .ZN(new_n422));
  INV_X1    g236(.A(G478), .ZN(new_n423));
  NOR2_X1   g237(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n225), .A2(G128), .ZN(new_n428));
  AND2_X1   g242(.A1(KEYINPUT92), .A2(KEYINPUT13), .ZN(new_n429));
  NOR2_X1   g243(.A1(KEYINPUT92), .A2(KEYINPUT13), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n225), .A2(G128), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n428), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n432), .B1(new_n429), .B2(new_n430), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT93), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT93), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n432), .B(new_n437), .C1(new_n429), .C2(new_n430), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n434), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G134), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n433), .A2(new_n428), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n198), .ZN(new_n442));
  NOR2_X1   g256(.A1(KEYINPUT91), .A2(G122), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(KEYINPUT91), .A2(G122), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n248), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G122), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n250), .B2(new_n251), .ZN(new_n448));
  OAI21_X1  g262(.A(G107), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n252), .A2(G122), .ZN(new_n450));
  INV_X1    g264(.A(new_n445), .ZN(new_n451));
  OAI21_X1  g265(.A(G116), .B1(new_n451), .B2(new_n443), .ZN(new_n452));
  INV_X1    g266(.A(G107), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n440), .A2(new_n442), .A3(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n441), .B(new_n198), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n453), .B1(new_n452), .B2(KEYINPUT14), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n448), .B2(new_n446), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n450), .B(new_n452), .C1(KEYINPUT14), .C2(new_n453), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n457), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT9), .B(G234), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n462), .A2(new_n362), .A3(G953), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n456), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n463), .B1(new_n456), .B2(new_n461), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n310), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT95), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n427), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n467), .ZN(new_n470));
  OAI211_X1 g284(.A(KEYINPUT95), .B(new_n310), .C1(new_n464), .C2(new_n465), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n427), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n422), .B(new_n469), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n470), .B2(new_n471), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT96), .B1(new_n475), .B2(new_n468), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n421), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(G214), .B1(G237), .B2(G902), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n193), .A2(G952), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(G234), .B2(G237), .ZN(new_n483));
  AOI211_X1 g297(.A(new_n193), .B(new_n310), .C1(G234), .C2(G237), .ZN(new_n484));
  XOR2_X1   g298(.A(KEYINPUT21), .B(G898), .Z(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n483), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n239), .A2(G125), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n488), .A2(KEYINPUT84), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(KEYINPUT84), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n259), .B(new_n322), .C1(new_n261), .C2(new_n262), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT85), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n492), .B(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G224), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(G953), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT7), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT86), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n497), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n495), .A2(KEYINPUT7), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT3), .B1(new_n392), .B2(G107), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT3), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n453), .A3(G104), .ZN(new_n505));
  INV_X1    g319(.A(G101), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n392), .A2(G107), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n503), .A2(new_n505), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n453), .A2(G104), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n392), .A2(G107), .ZN(new_n510));
  OAI21_X1  g324(.A(G101), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT81), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n253), .A2(new_n254), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n253), .A2(KEYINPUT5), .ZN(new_n516));
  OR3_X1    g330(.A1(new_n248), .A2(KEYINPUT5), .A3(G119), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(G113), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n514), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n503), .A2(new_n505), .A3(new_n507), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G101), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(KEYINPUT4), .A3(new_n508), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT79), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT79), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n521), .A2(new_n524), .A3(KEYINPUT4), .A4(new_n508), .ZN(new_n525));
  OR2_X1    g339(.A1(new_n521), .A2(KEYINPUT4), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n255), .A2(new_n523), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  XOR2_X1   g341(.A(G110), .B(G122), .Z(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n519), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n528), .B(KEYINPUT8), .Z(new_n532));
  NAND2_X1  g346(.A1(new_n518), .A2(new_n515), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(new_n512), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n531), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT86), .ZN(new_n536));
  OAI221_X1 g350(.A(new_n536), .B1(new_n498), .B2(new_n497), .C1(new_n491), .C2(new_n494), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n500), .A2(new_n502), .A3(new_n535), .A4(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n497), .B1(new_n491), .B2(new_n494), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n492), .B(KEYINPUT85), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n540), .A2(new_n501), .A3(new_n490), .A4(new_n489), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT6), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n519), .A2(new_n527), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n528), .B(KEYINPUT83), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n543), .B1(new_n546), .B2(new_n530), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT6), .B1(new_n544), .B2(new_n545), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n542), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n538), .A2(new_n400), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(G210), .B1(G237), .B2(G902), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n538), .A2(new_n400), .A3(new_n549), .A4(new_n551), .ZN(new_n554));
  AOI211_X1 g368(.A(new_n481), .B(new_n487), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G221), .B1(new_n462), .B2(G902), .ZN(new_n556));
  XNOR2_X1  g370(.A(G110), .B(G140), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n193), .A2(G227), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n557), .B(new_n558), .Z(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n523), .A2(new_n526), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT80), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n561), .A2(new_n562), .A3(new_n245), .A4(new_n525), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n245), .A2(new_n523), .A3(new_n525), .A4(new_n526), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT80), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n514), .A2(new_n263), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT10), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT10), .ZN(new_n569));
  INV_X1    g383(.A(new_n512), .ZN(new_n570));
  INV_X1    g384(.A(new_n259), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n260), .B1(new_n228), .B2(KEYINPUT1), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n257), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n566), .A2(new_n220), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n570), .B1(new_n571), .B2(new_n573), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n263), .B2(new_n570), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n578), .A2(KEYINPUT12), .A3(new_n243), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT12), .B1(new_n578), .B2(new_n243), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n560), .B1(new_n576), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n563), .A2(new_n565), .B1(new_n568), .B2(new_n574), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n560), .B1(new_n583), .B2(new_n220), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n566), .A2(new_n575), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n243), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(KEYINPUT82), .B(G469), .C1(new_n588), .C2(G902), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT82), .ZN(new_n590));
  AOI21_X1  g404(.A(G902), .B1(new_n582), .B2(new_n587), .ZN(new_n591));
  INV_X1    g405(.A(G469), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n576), .A2(new_n581), .A3(new_n560), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n583), .A2(new_n220), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n559), .B1(new_n586), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n592), .B(new_n310), .C1(new_n594), .C2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n589), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  AND4_X1   g412(.A1(new_n479), .A2(new_n555), .A3(new_n556), .A4(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n321), .A2(new_n369), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n556), .ZN(new_n602));
  OAI21_X1  g416(.A(G472), .B1(new_n299), .B2(new_n309), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n277), .A2(new_n278), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT31), .B1(new_n285), .B2(new_n195), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n295), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n188), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n369), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n602), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n466), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n423), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n464), .A2(new_n465), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT97), .B1(new_n456), .B2(new_n461), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n614), .B(new_n617), .Z(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n310), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n613), .B1(new_n619), .B2(G478), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n419), .B2(new_n420), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n555), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n610), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  NOR2_X1   g442(.A1(new_n412), .A2(new_n413), .ZN(new_n629));
  OAI22_X1  g443(.A1(new_n629), .A2(new_n410), .B1(new_n397), .B2(new_n398), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n624), .A2(new_n477), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n610), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT35), .B(G107), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT98), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n632), .B(new_n634), .ZN(G9));
  NOR2_X1   g449(.A1(new_n357), .A2(KEYINPUT36), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(new_n353), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n367), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n365), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n599), .A2(new_n607), .A3(new_n603), .A4(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n641), .B(KEYINPUT37), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G110), .ZN(G12));
  AOI211_X1 g457(.A(new_n481), .B(new_n639), .C1(new_n553), .C2(new_n554), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n556), .A3(new_n598), .ZN(new_n645));
  INV_X1    g459(.A(G900), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n483), .B1(new_n484), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n630), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n474), .A2(new_n648), .A3(new_n476), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(KEYINPUT99), .Z(new_n650));
  NOR2_X1   g464(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n321), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n319), .B1(new_n298), .B2(new_n300), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n649), .B(KEYINPUT99), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n655), .A2(new_n556), .A3(new_n598), .A4(new_n644), .ZN(new_n656));
  OAI21_X1  g470(.A(KEYINPUT100), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G128), .ZN(G30));
  NAND2_X1  g473(.A1(new_n553), .A2(new_n554), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n660), .B(KEYINPUT38), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n647), .B(KEYINPUT39), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n602), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n661), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n313), .A2(new_n195), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n303), .A2(new_n281), .ZN(new_n668));
  AOI21_X1  g482(.A(G902), .B1(new_n668), .B2(new_n293), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n302), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n298), .B2(new_n300), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT101), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n421), .A2(new_n478), .A3(new_n480), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n640), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n674), .B(KEYINPUT102), .Z(new_n675));
  NAND3_X1  g489(.A1(new_n666), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT103), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n225), .ZN(G45));
  AOI21_X1  g492(.A(new_n645), .B1(new_n301), .B2(new_n320), .ZN(new_n679));
  INV_X1    g493(.A(new_n647), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n622), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G146), .ZN(G48));
  NOR2_X1   g498(.A1(new_n594), .A2(new_n596), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n592), .B1(new_n686), .B2(new_n310), .ZN(new_n687));
  INV_X1    g501(.A(new_n597), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n556), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n321), .A2(new_n369), .A3(new_n625), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NAND4_X1  g508(.A1(new_n321), .A2(new_n631), .A3(new_n369), .A4(new_n691), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  INV_X1    g510(.A(new_n487), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n689), .A2(new_n697), .A3(new_n556), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n644), .A2(new_n479), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n321), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  INV_X1    g516(.A(new_n660), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n673), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT104), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n275), .A2(new_n255), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n290), .B1(new_n706), .B2(new_n269), .ZN(new_n707));
  INV_X1    g521(.A(new_n305), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n307), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n293), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n287), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n705), .B1(new_n711), .B2(new_n188), .ZN(new_n712));
  AOI211_X1 g526(.A(KEYINPUT104), .B(new_n189), .C1(new_n287), .C2(new_n710), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n714), .A2(KEYINPUT105), .A3(new_n369), .A4(new_n603), .ZN(new_n715));
  AOI22_X1  g529(.A1(new_n279), .A2(new_n286), .B1(new_n709), .B2(new_n293), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT104), .B1(new_n716), .B2(new_n189), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n711), .A2(new_n705), .A3(new_n188), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n717), .A2(new_n718), .A3(new_n369), .A4(new_n603), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI211_X1 g535(.A(new_n698), .B(new_n704), .C1(new_n715), .C2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n447), .ZN(G24));
  NAND4_X1  g537(.A1(new_n689), .A2(new_n622), .A3(new_n556), .A4(new_n680), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n644), .A2(new_n717), .A3(new_n718), .A4(new_n603), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT106), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n322), .ZN(G27));
  XNOR2_X1  g542(.A(new_n296), .B(new_n187), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n609), .B1(new_n729), .B2(new_n320), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n556), .A2(new_n480), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n660), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n597), .B1(new_n592), .B2(new_n591), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n622), .A2(new_n733), .A3(new_n680), .A4(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n730), .A2(KEYINPUT42), .A3(new_n736), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n654), .A2(new_n735), .A3(new_n609), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n738), .A2(KEYINPUT107), .ZN(new_n739));
  XOR2_X1   g553(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(new_n738), .B2(KEYINPUT107), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n737), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G131), .ZN(G33));
  NAND2_X1  g558(.A1(new_n321), .A2(new_n369), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n733), .A2(new_n734), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n745), .A2(new_n650), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n198), .ZN(G36));
  NAND2_X1  g562(.A1(new_n588), .A2(KEYINPUT45), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n582), .A2(new_n587), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(G469), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(G469), .A2(G902), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(KEYINPUT46), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n597), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n753), .A2(new_n754), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n759), .A2(KEYINPUT110), .A3(new_n760), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n755), .A2(KEYINPUT109), .A3(new_n597), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n758), .A2(new_n763), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n556), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n662), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n419), .A2(new_n620), .A3(new_n420), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n608), .A3(new_n640), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n660), .A2(new_n481), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n772), .B2(new_n773), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n768), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G137), .ZN(G39));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n767), .B(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n681), .A2(new_n369), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n321), .A2(new_n776), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n781), .A2(KEYINPUT111), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n767), .A2(new_n780), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT47), .B1(new_n766), .B2(new_n556), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n782), .B(new_n783), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT111), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT112), .Z(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G140), .ZN(G42));
  AOI22_X1  g606(.A1(new_n653), .A2(new_n657), .B1(new_n682), .B2(new_n679), .ZN(new_n793));
  INV_X1    g607(.A(new_n670), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT32), .B1(new_n607), .B2(KEYINPUT72), .ZN(new_n795));
  INV_X1    g609(.A(new_n300), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n556), .A3(new_n639), .A4(new_n734), .ZN(new_n798));
  INV_X1    g612(.A(new_n704), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n680), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT115), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n734), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n671), .A2(new_n640), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n704), .A2(new_n647), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n803), .A2(new_n804), .A3(new_n556), .A4(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n726), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n793), .A2(new_n801), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n475), .A2(new_n468), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n623), .B1(new_n421), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n602), .A2(new_n624), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n608), .A2(new_n609), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n695), .A2(new_n600), .A3(new_n641), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n692), .A2(new_n701), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n816), .A2(new_n722), .A3(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n714), .A2(new_n603), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n736), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n321), .A2(new_n811), .A3(new_n648), .A4(new_n775), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n820), .B1(new_n821), .B2(new_n602), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n747), .B1(new_n822), .B2(new_n640), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n818), .A2(new_n823), .A3(new_n743), .A4(KEYINPUT53), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT52), .B1(new_n808), .B2(KEYINPUT116), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n810), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n818), .A2(new_n743), .A3(new_n823), .ZN(new_n827));
  AOI221_X4 g641(.A(new_n726), .B1(new_n679), .B2(new_n682), .C1(new_n653), .C2(new_n657), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(KEYINPUT52), .A3(new_n801), .A4(new_n806), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n801), .A2(new_n806), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n658), .A2(new_n683), .A3(new_n807), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT53), .B1(new_n827), .B2(new_n834), .ZN(new_n835));
  OR3_X1    g649(.A1(new_n826), .A2(new_n835), .A3(KEYINPUT54), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n771), .A2(new_n483), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n689), .A2(new_n733), .ZN(new_n838));
  AND4_X1   g652(.A1(new_n640), .A2(new_n837), .A3(new_n819), .A4(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n672), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(new_n369), .A3(new_n483), .A4(new_n838), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n421), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n839), .B1(new_n842), .B2(new_n621), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n771), .A2(new_n483), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n715), .B2(new_n721), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n481), .A3(new_n661), .A4(new_n691), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT50), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n846), .B(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n689), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n556), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n775), .B(new_n845), .C1(new_n781), .C2(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n843), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n827), .A2(new_n834), .A3(KEYINPUT53), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n818), .A2(new_n743), .A3(new_n823), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n808), .A2(KEYINPUT116), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n830), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n818), .A2(new_n823), .A3(new_n743), .A4(KEYINPUT114), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n858), .A2(new_n860), .A3(new_n809), .A4(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n854), .B1(new_n855), .B2(new_n862), .ZN(new_n863));
  OAI221_X1 g677(.A(new_n836), .B1(KEYINPUT51), .B2(new_n852), .C1(new_n853), .C2(new_n863), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n841), .A2(new_n623), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT48), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n730), .A2(new_n837), .A3(new_n838), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n690), .A2(new_n481), .A3(new_n703), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n866), .A2(new_n867), .B1(new_n845), .B2(new_n868), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n867), .A2(new_n866), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n482), .B(KEYINPUT118), .Z(new_n871));
  NAND4_X1  g685(.A1(new_n865), .A2(new_n869), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT119), .Z(new_n873));
  NAND4_X1  g687(.A1(new_n843), .A2(KEYINPUT51), .A3(new_n848), .A4(new_n851), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n874), .A2(new_n875), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n873), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI22_X1  g692(.A1(new_n864), .A2(new_n878), .B1(G952), .B2(G953), .ZN(new_n879));
  OR2_X1    g693(.A1(KEYINPUT113), .A2(KEYINPUT49), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n732), .B1(new_n849), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(KEYINPUT113), .A2(KEYINPUT49), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n840), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n769), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n849), .A2(new_n880), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n884), .A2(new_n369), .A3(new_n661), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n879), .A2(new_n886), .ZN(G75));
  OAI211_X1 g701(.A(new_n309), .B(new_n552), .C1(new_n826), .C2(new_n835), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n547), .A2(new_n548), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(new_n542), .Z(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT55), .Z(new_n893));
  NAND2_X1  g707(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n193), .A2(G952), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n893), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n888), .A2(new_n889), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n894), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n894), .A2(KEYINPUT120), .A3(new_n896), .A4(new_n898), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(G51));
  AOI21_X1  g717(.A(new_n856), .B1(new_n833), .B2(new_n829), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n860), .A2(new_n809), .ZN(new_n905));
  OAI22_X1  g719(.A1(new_n904), .A2(KEYINPUT53), .B1(new_n905), .B2(new_n824), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT54), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n836), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n754), .A2(KEYINPUT57), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n754), .A2(KEYINPUT57), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n686), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n906), .A2(new_n309), .ZN(new_n913));
  INV_X1    g727(.A(new_n753), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n895), .B1(new_n912), .B2(new_n915), .ZN(G54));
  NAND3_X1  g730(.A1(new_n913), .A2(KEYINPUT58), .A3(G475), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(new_n396), .A3(new_n409), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n396), .A2(new_n409), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n913), .A2(KEYINPUT58), .A3(G475), .A4(new_n919), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n918), .A2(new_n896), .A3(new_n920), .ZN(G60));
  OAI21_X1  g735(.A(new_n836), .B1(new_n863), .B2(new_n853), .ZN(new_n922));
  NAND2_X1  g736(.A1(G478), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT59), .Z(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n618), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n908), .A2(new_n618), .A3(new_n925), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n895), .ZN(G63));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT60), .Z(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n826), .B2(new_n835), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n895), .B1(new_n931), .B2(new_n360), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n637), .B(KEYINPUT121), .Z(new_n933));
  OAI211_X1 g747(.A(new_n930), .B(new_n933), .C1(new_n826), .C2(new_n835), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(KEYINPUT122), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n906), .A2(new_n936), .A3(new_n930), .A4(new_n933), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n932), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT124), .ZN(new_n940));
  NAND2_X1  g754(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n938), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n940), .B1(new_n938), .B2(new_n941), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(G66));
  OAI21_X1  g758(.A(G953), .B1(new_n486), .B2(new_n496), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n818), .B2(G953), .ZN(new_n946));
  INV_X1    g760(.A(G898), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n891), .B1(new_n947), .B2(G953), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n946), .B(new_n948), .Z(G69));
  XNOR2_X1  g763(.A(new_n284), .B(new_n404), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(G900), .B2(G953), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n768), .A2(new_n799), .A3(new_n730), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n784), .B2(new_n789), .ZN(new_n953));
  INV_X1    g767(.A(new_n743), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT126), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n774), .A2(new_n777), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n956), .A2(new_n662), .A3(new_n767), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n955), .B1(new_n957), .B2(new_n832), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n778), .A2(KEYINPUT126), .A3(new_n828), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n954), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n747), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n953), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n951), .B1(new_n962), .B2(G953), .ZN(new_n963));
  INV_X1    g777(.A(new_n745), .ZN(new_n964));
  AND4_X1   g778(.A1(new_n964), .A2(new_n663), .A3(new_n775), .A4(new_n812), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n784), .B2(new_n789), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n828), .A2(new_n676), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT62), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n828), .A2(new_n676), .A3(KEYINPUT62), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n957), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(G953), .B1(new_n966), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n950), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n963), .B(KEYINPUT125), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n193), .B1(G227), .B2(G900), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n963), .B(KEYINPUT127), .C1(new_n972), .C2(new_n973), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n974), .A2(new_n975), .A3(new_n977), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(G72));
  NAND4_X1  g796(.A1(new_n953), .A2(new_n960), .A3(new_n961), .A4(new_n818), .ZN(new_n983));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  AOI211_X1 g799(.A(new_n195), .B(new_n313), .C1(new_n983), .C2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n966), .A2(new_n971), .A3(new_n818), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n987), .A2(new_n985), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n896), .B1(new_n988), .B2(new_n667), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n312), .A2(new_n315), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n863), .B1(new_n277), .B2(new_n990), .ZN(new_n991));
  AOI211_X1 g805(.A(new_n986), .B(new_n989), .C1(new_n985), .C2(new_n991), .ZN(G57));
endmodule


