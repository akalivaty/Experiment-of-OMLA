//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n538, new_n539, new_n540, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n559,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n587, new_n588,
    new_n589, new_n590, new_n593, new_n595, new_n596, new_n597, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1147, new_n1148;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n458));
  OAI21_X1  g033(.A(KEYINPUT64), .B1(new_n458), .B2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT3), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n465), .B1(new_n461), .B2(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n458), .A2(KEYINPUT65), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n463), .A2(new_n464), .A3(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  XOR2_X1   g047(.A(KEYINPUT3), .B(G2104), .Z(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n461), .A2(G2105), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n475), .A2(G2105), .B1(G101), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT66), .ZN(G160));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n468), .A2(G2105), .A3(new_n459), .A4(new_n462), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  OAI221_X1 g059(.A(new_n481), .B1(new_n482), .B2(new_n483), .C1(new_n469), .C2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  NOR4_X1   g062(.A1(new_n473), .A2(KEYINPUT4), .A3(new_n487), .A4(G2105), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n487), .A2(G2105), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n468), .A2(new_n459), .A3(new_n462), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT67), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n490), .A2(new_n493), .A3(KEYINPUT4), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n488), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G114), .C2(new_n464), .ZN(new_n497));
  INV_X1    g072(.A(G126), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n482), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n495), .A2(new_n499), .ZN(G164));
  AND2_X1   g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n504), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n508));
  XOR2_X1   g083(.A(KEYINPUT6), .B(G651), .Z(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n507), .A2(new_n510), .ZN(G166));
  NOR2_X1   g086(.A1(new_n509), .A2(new_n503), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G89), .ZN(new_n513));
  NAND3_X1  g088(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT7), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n509), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT68), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n519), .A2(G543), .A3(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n517), .B1(new_n523), .B2(G51), .ZN(G168));
  NAND2_X1  g099(.A1(new_n523), .A2(G52), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n526), .A2(new_n506), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n512), .A2(G90), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(G171));
  NAND2_X1  g105(.A1(new_n512), .A2(G81), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G43), .ZN(new_n533));
  OAI221_X1 g108(.A(new_n531), .B1(new_n532), .B2(new_n506), .C1(new_n522), .C2(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT69), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G860), .ZN(G153));
  NAND4_X1  g111(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g112(.A1(G1), .A2(G3), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT70), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT8), .ZN(new_n540));
  NAND4_X1  g115(.A1(G319), .A2(G483), .A3(G661), .A4(new_n540), .ZN(G188));
  NAND2_X1  g116(.A1(new_n523), .A2(G53), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT9), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT71), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT9), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n542), .B(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(G78), .A2(G543), .ZN(new_n550));
  XOR2_X1   g125(.A(new_n550), .B(KEYINPUT72), .Z(new_n551));
  INV_X1    g126(.A(G65), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n503), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g128(.A(G651), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n512), .A2(G91), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n549), .A2(new_n557), .ZN(G299));
  XNOR2_X1  g133(.A(new_n529), .B(KEYINPUT73), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(G301));
  INV_X1    g135(.A(G168), .ZN(G286));
  INV_X1    g136(.A(G166), .ZN(G303));
  NAND2_X1  g137(.A1(new_n512), .A2(G87), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n564));
  INV_X1    g139(.A(G49), .ZN(new_n565));
  OAI211_X1 g140(.A(new_n563), .B(new_n564), .C1(new_n522), .C2(new_n565), .ZN(G288));
  AOI22_X1  g141(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n567), .A2(new_n506), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n504), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(new_n509), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G305));
  NAND2_X1  g147(.A1(new_n512), .A2(G85), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  XOR2_X1   g149(.A(KEYINPUT74), .B(G47), .Z(new_n575));
  OAI221_X1 g150(.A(new_n573), .B1(new_n574), .B2(new_n506), .C1(new_n522), .C2(new_n575), .ZN(G290));
  NAND2_X1  g151(.A1(new_n512), .A2(G92), .ZN(new_n577));
  XOR2_X1   g152(.A(new_n577), .B(KEYINPUT10), .Z(new_n578));
  NAND2_X1  g153(.A1(new_n523), .A2(G54), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n506), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(G868), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(G868), .B2(new_n559), .ZN(G284));
  AOI21_X1  g160(.A(new_n584), .B1(G868), .B2(new_n559), .ZN(G321));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NOR2_X1   g162(.A1(G168), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT75), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n556), .B1(new_n544), .B2(new_n548), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n590), .B2(G868), .ZN(G297));
  XOR2_X1   g166(.A(G297), .B(KEYINPUT76), .Z(G280));
  INV_X1    g167(.A(G559), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n582), .B1(new_n593), .B2(G860), .ZN(G148));
  INV_X1    g169(.A(new_n535), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(new_n587), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n583), .A2(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n587), .ZN(G323));
  XNOR2_X1  g173(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g174(.A(new_n482), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G123), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT78), .Z(new_n602));
  NAND2_X1  g177(.A1(new_n470), .A2(G135), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n464), .A2(G111), .ZN(new_n604));
  OAI21_X1  g179(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n602), .B(new_n603), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT79), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(G2096), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(G2096), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT13), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n612), .A2(new_n613), .B1(new_n614), .B2(G2100), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n613), .B2(new_n612), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n614), .A2(G2100), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n609), .A2(new_n610), .A3(new_n618), .ZN(G156));
  XNOR2_X1  g194(.A(G2427), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT15), .B(G2435), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n623), .A2(KEYINPUT14), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(G1341), .B(G1348), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n625), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G2451), .B(G2454), .Z(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G14), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n629), .A2(new_n632), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n634), .A2(new_n635), .ZN(G401));
  XOR2_X1   g211(.A(G2072), .B(G2078), .Z(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2067), .B(G2678), .ZN(new_n639));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT18), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT81), .B(KEYINPUT17), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n637), .B(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n639), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI211_X1 g221(.A(new_n640), .B(new_n646), .C1(new_n645), .C2(new_n637), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n645), .A2(new_n640), .ZN(new_n648));
  AOI211_X1 g223(.A(new_n642), .B(new_n647), .C1(new_n644), .C2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2096), .B(G2100), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G227));
  XOR2_X1   g227(.A(G1971), .B(G1976), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT19), .ZN(new_n654));
  XOR2_X1   g229(.A(G1956), .B(G2474), .Z(new_n655));
  XOR2_X1   g230(.A(G1961), .B(G1966), .Z(new_n656));
  AND2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT20), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n655), .A2(new_n656), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT82), .ZN(new_n662));
  OR3_X1    g237(.A1(new_n654), .A2(new_n657), .A3(new_n660), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n659), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT83), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT84), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1991), .B(G1996), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1981), .B(G1986), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(G229));
  NAND2_X1  g250(.A1(new_n470), .A2(G141), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT92), .Z(new_n677));
  NAND2_X1  g252(.A1(new_n600), .A2(G129), .ZN(new_n678));
  NAND3_X1  g253(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT26), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  AOI22_X1  g257(.A1(new_n681), .A2(new_n682), .B1(G105), .B2(new_n476), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n677), .A2(new_n678), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT93), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n687), .B2(G32), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT27), .B(G1996), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT94), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT95), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n687), .A2(G26), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT28), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n470), .A2(G140), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n600), .A2(G128), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n464), .A2(G116), .ZN(new_n698));
  OAI21_X1  g273(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n696), .B(new_n697), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT89), .Z(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n695), .B1(new_n702), .B2(G29), .ZN(new_n703));
  INV_X1    g278(.A(G2067), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G19), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(new_n535), .B2(new_n706), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT88), .Z(new_n709));
  OAI22_X1  g284(.A1(new_n689), .A2(new_n691), .B1(G1341), .B2(new_n709), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n693), .A2(new_n705), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n706), .A2(G6), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n571), .B2(new_n706), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT86), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT32), .B(G1981), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(G166), .A2(new_n706), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n706), .B2(G22), .ZN(new_n718));
  INV_X1    g293(.A(G1971), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n706), .A2(G23), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G288), .B2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT33), .B(G1976), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT87), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n722), .A2(new_n724), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n718), .A2(new_n719), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n720), .A2(new_n725), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  OR3_X1    g303(.A1(new_n716), .A2(new_n728), .A3(KEYINPUT34), .ZN(new_n729));
  OAI21_X1  g304(.A(KEYINPUT34), .B1(new_n716), .B2(new_n728), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n687), .A2(G25), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n470), .A2(G131), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n600), .A2(G119), .ZN(new_n733));
  OR2_X1    g308(.A1(G95), .A2(G2105), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n734), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n732), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n731), .B1(new_n737), .B2(new_n687), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT35), .B(G1991), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(G16), .A2(G24), .ZN(new_n741));
  XNOR2_X1  g316(.A(G290), .B(KEYINPUT85), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(G16), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(G1986), .Z(new_n744));
  NAND4_X1  g319(.A1(new_n729), .A2(new_n730), .A3(new_n740), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT36), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n709), .A2(G1341), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n706), .A2(G4), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n582), .B2(new_n706), .ZN(new_n749));
  INV_X1    g324(.A(G1348), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n607), .A2(G29), .ZN(new_n752));
  INV_X1    g327(.A(G34), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n753), .B2(KEYINPUT24), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(KEYINPUT24), .B2(new_n753), .ZN(new_n755));
  INV_X1    g330(.A(G160), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(new_n687), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2084), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n747), .A2(new_n751), .A3(new_n752), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n706), .A2(G20), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT23), .Z(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G299), .B2(G16), .ZN(new_n762));
  INV_X1    g337(.A(G1956), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n470), .A2(G139), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT25), .Z(new_n767));
  INV_X1    g342(.A(G127), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n473), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G115), .B2(G2104), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n765), .B(new_n767), .C1(new_n464), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(new_n687), .ZN(new_n772));
  NOR2_X1   g347(.A1(G29), .A2(G33), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT90), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(G2072), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT31), .B(G11), .Z(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT96), .B(G28), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n778), .A2(KEYINPUT30), .ZN(new_n779));
  AOI21_X1  g354(.A(G29), .B1(new_n778), .B2(KEYINPUT30), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n777), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n775), .A2(G2072), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT91), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n776), .B(new_n781), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n706), .A2(G21), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G168), .B2(new_n706), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1966), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n706), .A2(G5), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G171), .B2(new_n706), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1961), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n784), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G29), .A2(G35), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G162), .B2(G29), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT29), .B(G2090), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  AOI211_X1 g371(.A(new_n795), .B(new_n796), .C1(new_n782), .C2(new_n783), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n687), .A2(G27), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT97), .ZN(new_n799));
  INV_X1    g374(.A(G164), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G29), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2078), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n791), .A2(new_n797), .A3(new_n802), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n759), .A2(new_n764), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n711), .A2(new_n746), .A3(new_n804), .ZN(G150));
  INV_X1    g380(.A(G150), .ZN(G311));
  AOI22_X1  g381(.A1(new_n523), .A2(G55), .B1(G93), .B2(new_n512), .ZN(new_n807));
  NAND2_X1  g382(.A1(G80), .A2(G543), .ZN(new_n808));
  INV_X1    g383(.A(G67), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n503), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT99), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n506), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n811), .B2(new_n810), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n807), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT101), .B(G860), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT102), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT37), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n535), .A2(new_n814), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(KEYINPUT100), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(KEYINPUT100), .ZN(new_n821));
  INV_X1    g396(.A(new_n814), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(new_n534), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n582), .A2(G559), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT39), .Z(new_n829));
  OAI21_X1  g404(.A(new_n818), .B1(new_n829), .B2(new_n815), .ZN(G145));
  NAND2_X1  g405(.A1(new_n470), .A2(G142), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n600), .A2(G130), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n464), .A2(G118), .ZN(new_n833));
  OAI21_X1  g408(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n831), .B(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT106), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n612), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n736), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n685), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT105), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n499), .A2(KEYINPUT104), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n463), .A2(G126), .A3(G2105), .A4(new_n468), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT104), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n842), .A2(new_n843), .A3(new_n497), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n840), .B1(new_n845), .B2(new_n495), .ZN(new_n846));
  INV_X1    g421(.A(new_n844), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n843), .B1(new_n842), .B2(new_n497), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n488), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n490), .A2(new_n493), .A3(KEYINPUT4), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n493), .B1(new_n490), .B2(KEYINPUT4), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n849), .A2(KEYINPUT105), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n846), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n771), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n701), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n839), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(G160), .B(KEYINPUT103), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(G162), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n608), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n858), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(KEYINPUT107), .B(G37), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g440(.A1(new_n590), .A2(new_n583), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT108), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(G299), .A2(new_n582), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n824), .B(new_n597), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n870), .A2(KEYINPUT41), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n869), .A2(new_n866), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n873), .B1(new_n878), .B2(new_n872), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n879), .A2(KEYINPUT42), .ZN(new_n880));
  XNOR2_X1  g455(.A(G290), .B(new_n571), .ZN(new_n881));
  XNOR2_X1  g456(.A(G166), .B(G288), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n881), .B(new_n882), .Z(new_n883));
  NAND2_X1  g458(.A1(new_n879), .A2(KEYINPUT42), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n880), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n883), .B1(new_n880), .B2(new_n884), .ZN(new_n886));
  OAI21_X1  g461(.A(G868), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(G868), .B2(new_n822), .ZN(G295));
  OAI21_X1  g463(.A(new_n887), .B1(G868), .B2(new_n822), .ZN(G331));
  AND2_X1   g464(.A1(new_n875), .A2(KEYINPUT41), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT111), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(G171), .A2(G168), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n893), .B1(new_n559), .B2(G168), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT109), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n824), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n824), .A2(new_n896), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n897), .A2(new_n898), .A3(new_n895), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n890), .A2(new_n891), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n892), .A2(new_n900), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n897), .A2(new_n898), .A3(new_n895), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n904), .A2(new_n899), .A3(new_n876), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n905), .B2(new_n871), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n883), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n870), .B1(new_n904), .B2(new_n899), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT110), .ZN(new_n909));
  INV_X1    g484(.A(new_n883), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n900), .A2(new_n874), .A3(new_n877), .A4(new_n901), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT110), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n912), .B(new_n870), .C1(new_n904), .C2(new_n899), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n909), .A2(new_n910), .A3(new_n911), .A4(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n907), .A2(new_n863), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n909), .A2(new_n911), .A3(new_n913), .ZN(new_n918));
  AOI21_X1  g493(.A(G37), .B1(new_n918), .B2(new_n883), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT43), .B1(new_n919), .B2(new_n914), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT44), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n915), .A2(KEYINPUT43), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n916), .B1(new_n919), .B2(new_n914), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n921), .A2(new_n925), .ZN(G397));
  INV_X1    g501(.A(G1996), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n686), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n685), .A2(G1996), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n701), .B(G2067), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n737), .A2(new_n739), .ZN(new_n932));
  OAI22_X1  g507(.A1(new_n931), .A2(new_n932), .B1(G2067), .B2(new_n702), .ZN(new_n933));
  INV_X1    g508(.A(G1384), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n846), .A2(new_n854), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n471), .A2(G40), .A3(new_n477), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n933), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n930), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n939), .B1(new_n941), .B2(new_n685), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n939), .A2(new_n927), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n943), .A2(KEYINPUT46), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n943), .A2(KEYINPUT46), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n946), .B(KEYINPUT47), .Z(new_n947));
  NOR4_X1   g522(.A1(new_n937), .A2(G1986), .A3(G290), .A4(new_n938), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT48), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(KEYINPUT48), .ZN(new_n950));
  INV_X1    g525(.A(new_n931), .ZN(new_n951));
  OR2_X1    g526(.A1(new_n737), .A2(new_n739), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n952), .A3(new_n932), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n950), .B1(new_n953), .B2(new_n939), .ZN(new_n954));
  AOI211_X1 g529(.A(new_n940), .B(new_n947), .C1(new_n949), .C2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G1384), .B1(new_n849), .B2(new_n853), .ZN(new_n956));
  INV_X1    g531(.A(new_n938), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(KEYINPUT114), .B(G8), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g535(.A(KEYINPUT115), .B(G1981), .Z(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n571), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1981), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(new_n571), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT49), .ZN(new_n966));
  AOI211_X1 g541(.A(G1976), .B(G288), .C1(new_n960), .C2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n963), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n960), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G1976), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n960), .B1(new_n970), .B2(G288), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT52), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT52), .B1(G288), .B2(new_n970), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n960), .B(new_n973), .C1(new_n970), .C2(G288), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n960), .A2(new_n966), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT116), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(G303), .A2(G8), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n981), .B1(new_n982), .B2(KEYINPUT55), .ZN(new_n983));
  XNOR2_X1  g558(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n983), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n934), .B1(new_n495), .B2(new_n499), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(KEYINPUT45), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n936), .A2(G1384), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n846), .A2(new_n854), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT112), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n846), .A2(new_n854), .A3(new_n992), .A4(new_n989), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n988), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(G1971), .B1(new_n994), .B2(new_n957), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n986), .A2(KEYINPUT50), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n853), .A2(new_n841), .A3(new_n844), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n998), .A3(new_n934), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n999), .A3(new_n957), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(G2090), .ZN(new_n1001));
  OAI211_X1 g576(.A(G8), .B(new_n985), .C1(new_n995), .C2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n969), .B1(new_n980), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n959), .ZN(new_n1004));
  INV_X1    g579(.A(G2090), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n956), .A2(new_n998), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT117), .B1(new_n1006), .B2(new_n938), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n987), .A2(new_n998), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT117), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1009), .B(new_n957), .C1(new_n956), .C2(new_n998), .ZN(new_n1010));
  AND4_X1   g585(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1004), .B1(new_n995), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n985), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n976), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n991), .A2(new_n993), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1016), .A2(G2078), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n957), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1018), .B1(new_n935), .B2(new_n936), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1015), .A2(KEYINPUT125), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1961), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1000), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT125), .B1(new_n1015), .B2(new_n1019), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G2078), .ZN(new_n1026));
  INV_X1    g601(.A(new_n988), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1015), .A2(new_n1026), .A3(new_n957), .A4(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n1016), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n529), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n989), .B1(new_n495), .B2(new_n499), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n957), .B(new_n1031), .C1(new_n956), .C2(KEYINPUT45), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n1033), .A2(new_n1017), .B1(new_n1000), .B2(new_n1021), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1029), .A2(G301), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT54), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1002), .B(new_n1014), .C1(new_n1030), .C2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n1038));
  INV_X1    g613(.A(G1966), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT45), .B1(new_n997), .B2(new_n934), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1031), .A2(new_n957), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1038), .B(new_n1039), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G2084), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n996), .A2(new_n999), .A3(new_n1043), .A4(new_n957), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1038), .B1(new_n1032), .B2(new_n1039), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(G168), .A2(new_n959), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n1051));
  OAI21_X1  g626(.A(G8), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1048), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1004), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1048), .A2(KEYINPUT51), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT123), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1055), .A2(KEYINPUT123), .A3(new_n1056), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1050), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT124), .B(KEYINPUT54), .ZN(new_n1061));
  AOI21_X1  g636(.A(G301), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1023), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1024), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1064), .A2(G301), .A3(new_n1029), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1061), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1037), .A2(new_n1060), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n543), .A2(new_n1069), .A3(new_n557), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n590), .B2(new_n1069), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1071), .B1(new_n1072), .B2(new_n763), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT56), .B(G2072), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n994), .A2(new_n957), .A3(new_n1074), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1072), .A2(new_n763), .ZN(new_n1078));
  NAND2_X1  g653(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1078), .A2(new_n1075), .B1(new_n1079), .B2(new_n1070), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1000), .A2(new_n750), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n958), .A2(new_n704), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n583), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1077), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT61), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT60), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1081), .A2(KEYINPUT60), .A3(new_n1082), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n582), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1081), .A2(KEYINPUT60), .A3(new_n583), .A4(new_n1082), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1087), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1085), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1078), .A2(new_n1075), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1071), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1091), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1086), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n956), .A2(new_n957), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT58), .B(G1341), .Z(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1097), .A2(KEYINPUT121), .A3(new_n1098), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n938), .A2(G1996), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n994), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT122), .B1(new_n1105), .B2(new_n595), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n994), .A2(new_n1104), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1107), .B(new_n535), .C1(new_n1108), .C2(new_n1103), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1106), .A2(KEYINPUT59), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n1111));
  OAI211_X1 g686(.A(KEYINPUT122), .B(new_n1111), .C1(new_n1105), .C2(new_n595), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1084), .B1(new_n1096), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1003), .B1(new_n1068), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n978), .A2(new_n979), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1047), .A2(G168), .A3(new_n1004), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1118), .A2(KEYINPUT63), .ZN(new_n1119));
  OAI21_X1  g694(.A(G8), .B1(new_n995), .B2(new_n1001), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1013), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1116), .A2(new_n1119), .A3(new_n1002), .A4(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1014), .A2(new_n1118), .A3(new_n1002), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT119), .B(KEYINPUT63), .Z(new_n1125));
  AND3_X1   g700(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1124), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1122), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1059), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1129), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT62), .B1(new_n1130), .B2(new_n1050), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1132), .B(new_n1049), .C1(new_n1133), .C2(new_n1129), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1014), .A2(new_n1002), .A3(new_n1062), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT126), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1131), .A2(new_n1134), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1131), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT126), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1115), .A2(new_n1128), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(G290), .B(G1986), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n939), .B1(new_n953), .B2(new_n1141), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1140), .A2(KEYINPUT127), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT127), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n955), .B1(new_n1143), .B2(new_n1144), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g720(.A(new_n651), .B(G319), .C1(new_n635), .C2(new_n634), .ZN(new_n1147));
  AOI21_X1  g721(.A(new_n1147), .B1(new_n673), .B2(new_n674), .ZN(new_n1148));
  OAI211_X1 g722(.A(new_n864), .B(new_n1148), .C1(new_n923), .C2(new_n924), .ZN(G225));
  INV_X1    g723(.A(G225), .ZN(G308));
endmodule


