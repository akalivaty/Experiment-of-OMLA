

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785;

  OR2_X1 U377 ( .A1(n743), .A2(n500), .ZN(n499) );
  XNOR2_X1 U378 ( .A(n769), .B(n559), .ZN(n595) );
  XNOR2_X1 U379 ( .A(G134), .B(n357), .ZN(n533) );
  BUF_X1 U380 ( .A(G122), .Z(n357) );
  BUF_X1 U381 ( .A(G143), .Z(n356) );
  INV_X1 U382 ( .A(G953), .ZN(n776) );
  NOR2_X2 U383 ( .A1(n602), .A2(n623), .ZN(n597) );
  XOR2_X1 U384 ( .A(G116), .B(G107), .Z(n550) );
  XNOR2_X2 U385 ( .A(n415), .B(KEYINPUT41), .ZN(n643) );
  NOR2_X2 U386 ( .A1(n388), .A2(n390), .ZN(n387) );
  NOR2_X2 U387 ( .A1(n757), .A2(n517), .ZN(n662) );
  NOR2_X2 U388 ( .A1(n757), .A2(n774), .ZN(n733) );
  XNOR2_X2 U389 ( .A(n385), .B(n373), .ZN(n757) );
  XNOR2_X2 U390 ( .A(n446), .B(n445), .ZN(n785) );
  NOR2_X1 U391 ( .A1(n681), .A2(n676), .ZN(n714) );
  NOR2_X2 U392 ( .A1(n610), .A2(n611), .ZN(n681) );
  XNOR2_X1 U393 ( .A(n595), .B(n560), .ZN(n575) );
  NOR2_X1 U394 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X2 U395 ( .A1(n642), .A2(n606), .ZN(n636) );
  INV_X1 U396 ( .A(n681), .ZN(n684) );
  INV_X1 U397 ( .A(n609), .ZN(n611) );
  AND2_X1 U398 ( .A1(n616), .A2(n492), .ZN(n490) );
  NOR2_X1 U399 ( .A1(n436), .A2(KEYINPUT44), .ZN(n510) );
  NAND2_X1 U400 ( .A1(n497), .A2(n495), .ZN(n700) );
  NOR2_X1 U401 ( .A1(n684), .A2(n630), .ZN(n652) );
  XNOR2_X1 U402 ( .A(n485), .B(n416), .ZN(n713) );
  XNOR2_X1 U403 ( .A(n745), .B(n744), .ZN(n746) );
  XNOR2_X1 U404 ( .A(n548), .B(n547), .ZN(n609) );
  XOR2_X1 U405 ( .A(n748), .B(n747), .Z(n374) );
  XNOR2_X1 U406 ( .A(n440), .B(n575), .ZN(n743) );
  NOR2_X1 U407 ( .A1(G902), .A2(n748), .ZN(n548) );
  XOR2_X1 U408 ( .A(n751), .B(KEYINPUT122), .Z(n376) );
  XOR2_X1 U409 ( .A(n664), .B(n529), .Z(n375) );
  XNOR2_X1 U410 ( .A(n546), .B(n358), .ZN(n748) );
  XNOR2_X1 U411 ( .A(n768), .B(n545), .ZN(n358) );
  XNOR2_X1 U412 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U413 ( .A(n451), .B(G125), .ZN(n555) );
  XOR2_X1 U414 ( .A(KEYINPUT3), .B(G119), .Z(n588) );
  NAND2_X1 U415 ( .A1(n750), .A2(G210), .ZN(n742) );
  AND2_X2 U416 ( .A1(n459), .A2(n460), .ZN(n750) );
  NOR2_X1 U417 ( .A1(n609), .A2(n610), .ZN(n600) );
  NAND2_X1 U418 ( .A1(n359), .A2(n371), .ZN(n414) );
  NAND2_X1 U419 ( .A1(n410), .A2(n413), .ZN(n359) );
  NAND2_X2 U420 ( .A1(n783), .A2(n675), .ZN(n622) );
  XNOR2_X2 U421 ( .A(n621), .B(n620), .ZN(n783) );
  INV_X1 U422 ( .A(G472), .ZN(n422) );
  NOR2_X1 U423 ( .A1(G902), .A2(n664), .ZN(n596) );
  NOR2_X1 U424 ( .A1(n457), .A2(n498), .ZN(n497) );
  INV_X1 U425 ( .A(KEYINPUT84), .ZN(n432) );
  NAND2_X1 U426 ( .A1(G234), .A2(G237), .ZN(n569) );
  XNOR2_X1 U427 ( .A(KEYINPUT73), .B(G110), .ZN(n560) );
  NAND2_X1 U428 ( .A1(n576), .A2(n501), .ZN(n500) );
  INV_X1 U429 ( .A(G902), .ZN(n501) );
  XNOR2_X1 U430 ( .A(n480), .B(n479), .ZN(n660) );
  INV_X1 U431 ( .A(KEYINPUT39), .ZN(n479) );
  AND2_X1 U432 ( .A1(n512), .A2(n700), .ZN(n619) );
  XNOR2_X1 U433 ( .A(n481), .B(n449), .ZN(n383) );
  INV_X1 U434 ( .A(KEYINPUT22), .ZN(n449) );
  INV_X1 U435 ( .A(n531), .ZN(n431) );
  INV_X1 U436 ( .A(n647), .ZN(n425) );
  XNOR2_X1 U437 ( .A(n682), .B(n649), .ZN(n450) );
  NAND2_X1 U438 ( .A1(n427), .A2(n365), .ZN(n426) );
  INV_X1 U439 ( .A(n785), .ZN(n410) );
  NAND2_X1 U440 ( .A1(n413), .A2(n412), .ZN(n411) );
  NOR2_X1 U441 ( .A1(n785), .A2(n371), .ZN(n412) );
  NOR2_X1 U442 ( .A1(n492), .A2(n439), .ZN(n435) );
  NAND2_X1 U443 ( .A1(n504), .A2(n503), .ZN(n494) );
  NAND2_X1 U444 ( .A1(n505), .A2(G902), .ZN(n503) );
  INV_X1 U445 ( .A(KEYINPUT48), .ZN(n452) );
  XNOR2_X1 U446 ( .A(n573), .B(G134), .ZN(n773) );
  XNOR2_X1 U447 ( .A(n572), .B(n508), .ZN(n767) );
  INV_X1 U448 ( .A(KEYINPUT97), .ZN(n508) );
  INV_X1 U449 ( .A(G146), .ZN(n451) );
  XNOR2_X1 U450 ( .A(n516), .B(n515), .ZN(n584) );
  INV_X1 U451 ( .A(KEYINPUT8), .ZN(n515) );
  NAND2_X1 U452 ( .A1(n776), .A2(G234), .ZN(n516) );
  XNOR2_X1 U453 ( .A(n444), .B(n574), .ZN(n443) );
  INV_X1 U454 ( .A(G107), .ZN(n574) );
  NAND2_X1 U455 ( .A1(n776), .A2(G227), .ZN(n444) );
  XNOR2_X1 U456 ( .A(n442), .B(G104), .ZN(n441) );
  INV_X1 U457 ( .A(G140), .ZN(n442) );
  INV_X1 U458 ( .A(n767), .ZN(n507) );
  INV_X1 U459 ( .A(KEYINPUT67), .ZN(n558) );
  XNOR2_X1 U460 ( .A(n773), .B(G146), .ZN(n594) );
  XOR2_X1 U461 ( .A(KEYINPUT9), .B(KEYINPUT105), .Z(n534) );
  XNOR2_X1 U462 ( .A(n544), .B(n543), .ZN(n545) );
  NAND2_X1 U463 ( .A1(n700), .A2(n699), .ZN(n602) );
  NAND2_X1 U464 ( .A1(n721), .A2(n712), .ZN(n415) );
  NAND2_X1 U465 ( .A1(n382), .A2(n571), .ZN(n384) );
  XOR2_X1 U466 ( .A(G478), .B(n537), .Z(n610) );
  NOR2_X1 U467 ( .A1(n637), .A2(n638), .ZN(n403) );
  BUF_X1 U468 ( .A(n645), .Z(n485) );
  AND2_X1 U469 ( .A1(n521), .A2(n520), .ZN(n648) );
  INV_X1 U470 ( .A(n642), .ZN(n520) );
  XNOR2_X1 U471 ( .A(n706), .B(KEYINPUT6), .ZN(n623) );
  OR2_X1 U472 ( .A1(n754), .A2(G902), .ZN(n522) );
  INV_X1 U473 ( .A(n700), .ZN(n448) );
  NAND2_X1 U474 ( .A1(n425), .A2(n432), .ZN(n424) );
  XOR2_X1 U475 ( .A(n714), .B(KEYINPUT85), .Z(n650) );
  AND2_X1 U476 ( .A1(n409), .A2(n408), .ZN(n407) );
  NAND2_X1 U477 ( .A1(n406), .A2(n405), .ZN(n404) );
  NOR2_X1 U478 ( .A1(n659), .A2(KEYINPUT71), .ZN(n405) );
  INV_X1 U479 ( .A(KEYINPUT4), .ZN(n556) );
  INV_X1 U480 ( .A(KEYINPUT16), .ZN(n526) );
  XNOR2_X1 U481 ( .A(G137), .B(KEYINPUT70), .ZN(n586) );
  XNOR2_X1 U482 ( .A(KEYINPUT15), .B(G902), .ZN(n577) );
  XNOR2_X1 U483 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n540) );
  INV_X1 U484 ( .A(KEYINPUT103), .ZN(n543) );
  XNOR2_X1 U485 ( .A(n555), .B(n367), .ZN(n524) );
  NOR2_X1 U486 ( .A1(G902), .A2(G237), .ZN(n561) );
  AND2_X1 U487 ( .A1(n717), .A2(n713), .ZN(n721) );
  AND2_X1 U488 ( .A1(n499), .A2(KEYINPUT1), .ZN(n496) );
  AND2_X1 U489 ( .A1(n494), .A2(n493), .ZN(n457) );
  XNOR2_X1 U490 ( .A(n600), .B(KEYINPUT106), .ZN(n717) );
  NAND2_X1 U491 ( .A1(n697), .A2(n454), .ZN(n453) );
  INV_X1 U492 ( .A(n638), .ZN(n454) );
  XNOR2_X1 U493 ( .A(G116), .B(G113), .ZN(n591) );
  NOR2_X1 U494 ( .A1(n694), .A2(n519), .ZN(n518) );
  INV_X1 U495 ( .A(n693), .ZN(n519) );
  XNOR2_X1 U496 ( .A(n587), .B(n360), .ZN(n397) );
  XOR2_X1 U497 ( .A(KEYINPUT86), .B(KEYINPUT79), .Z(n587) );
  XNOR2_X1 U498 ( .A(n586), .B(KEYINPUT23), .ZN(n395) );
  XNOR2_X1 U499 ( .A(n392), .B(n538), .ZN(n768) );
  XOR2_X1 U500 ( .A(KEYINPUT68), .B(KEYINPUT10), .Z(n538) );
  XNOR2_X1 U501 ( .A(n555), .B(G140), .ZN(n392) );
  INV_X1 U502 ( .A(KEYINPUT87), .ZN(n468) );
  XNOR2_X1 U503 ( .A(n506), .B(n594), .ZN(n440) );
  XNOR2_X1 U504 ( .A(n509), .B(n507), .ZN(n506) );
  XNOR2_X1 U505 ( .A(n443), .B(n441), .ZN(n509) );
  NOR2_X1 U506 ( .A1(n602), .A2(n421), .ZN(n708) );
  INV_X1 U507 ( .A(KEYINPUT96), .ZN(n475) );
  XNOR2_X1 U508 ( .A(n419), .B(n418), .ZN(n664) );
  XNOR2_X1 U509 ( .A(n514), .B(n420), .ZN(n418) );
  XNOR2_X1 U510 ( .A(n595), .B(n594), .ZN(n419) );
  XNOR2_X1 U511 ( .A(n588), .B(KEYINPUT76), .ZN(n420) );
  BUF_X1 U512 ( .A(n776), .Z(n471) );
  XNOR2_X1 U513 ( .A(n393), .B(n768), .ZN(n754) );
  XNOR2_X1 U514 ( .A(n396), .B(n394), .ZN(n393) );
  XNOR2_X1 U515 ( .A(n585), .B(n395), .ZN(n394) );
  XNOR2_X1 U516 ( .A(n398), .B(n397), .ZN(n396) );
  XNOR2_X1 U517 ( .A(n484), .B(n458), .ZN(n751) );
  XNOR2_X1 U518 ( .A(n535), .B(n366), .ZN(n484) );
  XNOR2_X1 U519 ( .A(n536), .B(n532), .ZN(n458) );
  XNOR2_X1 U520 ( .A(n597), .B(KEYINPUT33), .ZN(n723) );
  INV_X1 U521 ( .A(n643), .ZN(n711) );
  INV_X1 U522 ( .A(KEYINPUT42), .ZN(n445) );
  INV_X1 U523 ( .A(KEYINPUT40), .ZN(n391) );
  XNOR2_X1 U524 ( .A(n646), .B(KEYINPUT107), .ZN(n434) );
  AND2_X1 U525 ( .A1(n618), .A2(n456), .ZN(n666) );
  INV_X1 U526 ( .A(KEYINPUT60), .ZN(n464) );
  XOR2_X1 U527 ( .A(G128), .B(G119), .Z(n360) );
  XOR2_X1 U528 ( .A(n583), .B(n582), .Z(n361) );
  XOR2_X1 U529 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n362) );
  XOR2_X1 U530 ( .A(n524), .B(n554), .Z(n363) );
  XNOR2_X1 U531 ( .A(KEYINPUT82), .B(n619), .ZN(n364) );
  AND2_X1 U532 ( .A1(n647), .A2(n432), .ZN(n365) );
  XNOR2_X1 U533 ( .A(KEYINPUT104), .B(KEYINPUT7), .ZN(n366) );
  AND2_X1 U534 ( .A1(G224), .A2(n776), .ZN(n367) );
  OR2_X1 U535 ( .A1(n733), .A2(KEYINPUT2), .ZN(n368) );
  AND2_X1 U536 ( .A1(n531), .A2(KEYINPUT84), .ZN(n369) );
  INV_X1 U537 ( .A(n696), .ZN(n513) );
  XOR2_X1 U538 ( .A(KEYINPUT66), .B(KEYINPUT0), .Z(n370) );
  XNOR2_X1 U539 ( .A(n644), .B(KEYINPUT64), .ZN(n371) );
  XOR2_X1 U540 ( .A(KEYINPUT89), .B(KEYINPUT35), .Z(n372) );
  INV_X1 U541 ( .A(n756), .ZN(n483) );
  XOR2_X1 U542 ( .A(KEYINPUT88), .B(KEYINPUT45), .Z(n373) );
  XOR2_X1 U543 ( .A(n740), .B(n741), .Z(n377) );
  NAND2_X1 U544 ( .A1(n663), .A2(KEYINPUT2), .ZN(n378) );
  XOR2_X1 U545 ( .A(KEYINPUT90), .B(KEYINPUT56), .Z(n379) );
  XOR2_X1 U546 ( .A(n357), .B(KEYINPUT126), .Z(n380) );
  NAND2_X1 U547 ( .A1(n381), .A2(KEYINPUT44), .ZN(n447) );
  INV_X1 U548 ( .A(n511), .ZN(n381) );
  XNOR2_X2 U549 ( .A(n622), .B(KEYINPUT93), .ZN(n511) );
  AND2_X1 U550 ( .A1(n382), .A2(n648), .ZN(n682) );
  XNOR2_X2 U551 ( .A(n654), .B(KEYINPUT19), .ZN(n382) );
  NAND2_X1 U552 ( .A1(n383), .A2(n364), .ZN(n621) );
  AND2_X1 U553 ( .A1(n383), .A2(n448), .ZN(n618) );
  XNOR2_X2 U554 ( .A(n384), .B(n370), .ZN(n603) );
  NAND2_X2 U555 ( .A1(n645), .A2(n712), .ZN(n654) );
  NAND2_X1 U556 ( .A1(n387), .A2(n386), .ZN(n385) );
  XNOR2_X1 U557 ( .A(n389), .B(KEYINPUT74), .ZN(n386) );
  NAND2_X1 U558 ( .A1(n489), .A2(n447), .ZN(n388) );
  NAND2_X1 U559 ( .A1(n510), .A2(n511), .ZN(n389) );
  NAND2_X1 U560 ( .A1(n487), .A2(n486), .ZN(n390) );
  XNOR2_X1 U561 ( .A(n413), .B(G131), .ZN(G33) );
  XNOR2_X2 U562 ( .A(n639), .B(n391), .ZN(n413) );
  NAND2_X1 U563 ( .A1(n584), .A2(G221), .ZN(n398) );
  NAND2_X2 U564 ( .A1(n399), .A2(n518), .ZN(n774) );
  XNOR2_X2 U565 ( .A(n400), .B(n452), .ZN(n399) );
  NAND2_X1 U566 ( .A1(n402), .A2(n401), .ZN(n400) );
  NAND2_X1 U567 ( .A1(n407), .A2(n404), .ZN(n401) );
  NAND2_X1 U568 ( .A1(n414), .A2(n411), .ZN(n402) );
  NAND2_X1 U569 ( .A1(n403), .A2(n713), .ZN(n480) );
  NAND2_X1 U570 ( .A1(n403), .A2(n485), .ZN(n646) );
  INV_X1 U571 ( .A(n658), .ZN(n406) );
  NAND2_X1 U572 ( .A1(n659), .A2(KEYINPUT71), .ZN(n408) );
  NAND2_X1 U573 ( .A1(n658), .A2(KEYINPUT71), .ZN(n409) );
  INV_X1 U574 ( .A(KEYINPUT38), .ZN(n416) );
  BUF_X1 U575 ( .A(n436), .Z(n417) );
  AND2_X1 U576 ( .A1(n623), .A2(n696), .ZN(n456) );
  BUF_X1 U577 ( .A(n706), .Z(n478) );
  AND2_X1 U578 ( .A1(n623), .A2(n513), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n417), .B(n380), .ZN(G24) );
  XNOR2_X2 U580 ( .A(n476), .B(n372), .ZN(n436) );
  XNOR2_X2 U581 ( .A(n557), .B(n556), .ZN(n769) );
  INV_X1 U582 ( .A(n706), .ZN(n421) );
  XNOR2_X2 U583 ( .A(n596), .B(n422), .ZN(n706) );
  NAND2_X1 U584 ( .A1(n424), .A2(n423), .ZN(n429) );
  NAND2_X1 U585 ( .A1(n647), .A2(n430), .ZN(n423) );
  NAND2_X1 U586 ( .A1(n434), .A2(n369), .ZN(n433) );
  NAND2_X1 U587 ( .A1(n434), .A2(n531), .ZN(n679) );
  NAND2_X1 U588 ( .A1(n428), .A2(n426), .ZN(n659) );
  INV_X1 U589 ( .A(n434), .ZN(n427) );
  AND2_X1 U590 ( .A1(n433), .A2(n429), .ZN(n428) );
  NAND2_X1 U591 ( .A1(n431), .A2(n432), .ZN(n430) );
  NAND2_X1 U592 ( .A1(n436), .A2(KEYINPUT44), .ZN(n491) );
  NAND2_X1 U593 ( .A1(n436), .A2(n435), .ZN(n486) );
  XNOR2_X2 U594 ( .A(n437), .B(n363), .ZN(n523) );
  XNOR2_X1 U595 ( .A(n437), .B(G101), .ZN(n762) );
  XNOR2_X2 U596 ( .A(n525), .B(n438), .ZN(n437) );
  INV_X1 U597 ( .A(n551), .ZN(n438) );
  INV_X1 U598 ( .A(KEYINPUT44), .ZN(n439) );
  NOR2_X1 U599 ( .A1(n499), .A2(KEYINPUT1), .ZN(n498) );
  NAND2_X1 U600 ( .A1(n643), .A2(n648), .ZN(n446) );
  NAND2_X1 U601 ( .A1(n651), .A2(n450), .ZN(n455) );
  NOR2_X1 U602 ( .A1(n696), .A2(n453), .ZN(n640) );
  XNOR2_X2 U603 ( .A(n522), .B(n361), .ZN(n696) );
  AND2_X1 U604 ( .A1(n460), .A2(n368), .ZN(n734) );
  XNOR2_X1 U605 ( .A(n461), .B(KEYINPUT78), .ZN(n460) );
  NAND2_X1 U606 ( .A1(n603), .A2(n601), .ZN(n481) );
  NAND2_X1 U607 ( .A1(n455), .A2(n691), .ZN(n658) );
  NOR2_X2 U608 ( .A1(n607), .A2(n723), .ZN(n598) );
  NOR2_X1 U609 ( .A1(n653), .A2(n654), .ZN(n656) );
  XNOR2_X1 U610 ( .A(n774), .B(n661), .ZN(n517) );
  NAND2_X1 U611 ( .A1(n467), .A2(n378), .ZN(n459) );
  XNOR2_X1 U612 ( .A(n528), .B(n746), .ZN(n462) );
  NAND2_X1 U613 ( .A1(n733), .A2(KEYINPUT2), .ZN(n461) );
  NAND2_X1 U614 ( .A1(n462), .A2(n483), .ZN(n527) );
  XNOR2_X1 U615 ( .A(n463), .B(n379), .ZN(G51) );
  NAND2_X1 U616 ( .A1(n474), .A2(n483), .ZN(n463) );
  XNOR2_X1 U617 ( .A(n465), .B(n464), .ZN(G60) );
  NAND2_X1 U618 ( .A1(n472), .A2(n483), .ZN(n465) );
  XNOR2_X1 U619 ( .A(n466), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U620 ( .A1(n473), .A2(n483), .ZN(n466) );
  XNOR2_X1 U621 ( .A(n469), .B(n468), .ZN(n467) );
  NAND2_X1 U622 ( .A1(n662), .A2(n663), .ZN(n469) );
  NAND2_X1 U623 ( .A1(n470), .A2(n483), .ZN(n482) );
  XNOR2_X1 U624 ( .A(n752), .B(n376), .ZN(n470) );
  XNOR2_X1 U625 ( .A(n641), .B(KEYINPUT28), .ZN(n521) );
  XNOR2_X1 U626 ( .A(n749), .B(n374), .ZN(n472) );
  XNOR2_X1 U627 ( .A(n665), .B(n375), .ZN(n473) );
  XNOR2_X1 U628 ( .A(n742), .B(n377), .ZN(n474) );
  XNOR2_X1 U629 ( .A(n603), .B(n475), .ZN(n607) );
  NAND2_X1 U630 ( .A1(n599), .A2(n531), .ZN(n476) );
  NAND2_X1 U631 ( .A1(n477), .A2(n636), .ZN(n637) );
  XNOR2_X1 U632 ( .A(n635), .B(n634), .ZN(n477) );
  XOR2_X2 U633 ( .A(G131), .B(KEYINPUT69), .Z(n573) );
  NAND2_X1 U634 ( .A1(n696), .A2(n697), .ZN(n606) );
  XNOR2_X1 U635 ( .A(n482), .B(KEYINPUT123), .ZN(G63) );
  XNOR2_X2 U636 ( .A(n523), .B(n575), .ZN(n740) );
  NAND2_X1 U637 ( .A1(n488), .A2(KEYINPUT92), .ZN(n487) );
  INV_X1 U638 ( .A(n616), .ZN(n488) );
  NAND2_X1 U639 ( .A1(n491), .A2(n490), .ZN(n489) );
  INV_X1 U640 ( .A(KEYINPUT92), .ZN(n492) );
  INV_X1 U641 ( .A(n494), .ZN(n502) );
  INV_X1 U642 ( .A(KEYINPUT1), .ZN(n493) );
  NAND2_X1 U643 ( .A1(n502), .A2(n499), .ZN(n642) );
  NAND2_X1 U644 ( .A1(n496), .A2(n502), .ZN(n495) );
  NAND2_X1 U645 ( .A1(n743), .A2(n505), .ZN(n504) );
  INV_X1 U646 ( .A(n576), .ZN(n505) );
  XNOR2_X1 U647 ( .A(n593), .B(n590), .ZN(n514) );
  XNOR2_X2 U648 ( .A(n549), .B(n526), .ZN(n525) );
  XNOR2_X1 U649 ( .A(n527), .B(KEYINPUT121), .ZN(G54) );
  NAND2_X1 U650 ( .A1(n750), .A2(G469), .ZN(n528) );
  XNOR2_X2 U651 ( .A(n539), .B(G104), .ZN(n549) );
  XNOR2_X2 U652 ( .A(G113), .B(G122), .ZN(n539) );
  XNOR2_X1 U653 ( .A(KEYINPUT62), .B(KEYINPUT108), .ZN(n529) );
  AND2_X1 U654 ( .A1(G214), .A2(n589), .ZN(n530) );
  AND2_X1 U655 ( .A1(n609), .A2(n610), .ZN(n531) );
  INV_X1 U656 ( .A(KEYINPUT47), .ZN(n649) );
  INV_X1 U657 ( .A(KEYINPUT30), .ZN(n634) );
  XNOR2_X1 U658 ( .A(n558), .B(G101), .ZN(n559) );
  INV_X1 U659 ( .A(KEYINPUT83), .ZN(n562) );
  XNOR2_X1 U660 ( .A(KEYINPUT36), .B(KEYINPUT94), .ZN(n655) );
  XNOR2_X1 U661 ( .A(n656), .B(n655), .ZN(n657) );
  NOR2_X1 U662 ( .A1(G952), .A2(n471), .ZN(n756) );
  INV_X1 U663 ( .A(n577), .ZN(n663) );
  NAND2_X1 U664 ( .A1(G217), .A2(n584), .ZN(n532) );
  XNOR2_X1 U665 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X2 U666 ( .A(G143), .B(G128), .Z(n557) );
  XNOR2_X1 U667 ( .A(n557), .B(n550), .ZN(n536) );
  NOR2_X1 U668 ( .A1(G902), .A2(n751), .ZN(n537) );
  NOR2_X1 U669 ( .A1(G953), .A2(G237), .ZN(n589) );
  XNOR2_X1 U670 ( .A(n549), .B(n530), .ZN(n542) );
  XNOR2_X1 U671 ( .A(n362), .B(n540), .ZN(n541) );
  XNOR2_X1 U672 ( .A(n542), .B(n541), .ZN(n546) );
  XNOR2_X1 U673 ( .A(n573), .B(n356), .ZN(n544) );
  XNOR2_X1 U674 ( .A(KEYINPUT13), .B(G475), .ZN(n547) );
  XNOR2_X1 U675 ( .A(n588), .B(n550), .ZN(n551) );
  XOR2_X1 U676 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n553) );
  XNOR2_X1 U677 ( .A(KEYINPUT81), .B(KEYINPUT80), .ZN(n552) );
  XNOR2_X1 U678 ( .A(n553), .B(n552), .ZN(n554) );
  NOR2_X2 U679 ( .A1(n740), .A2(n663), .ZN(n565) );
  XNOR2_X1 U680 ( .A(n561), .B(KEYINPUT75), .ZN(n566) );
  NAND2_X1 U681 ( .A1(G210), .A2(n566), .ZN(n563) );
  XNOR2_X2 U682 ( .A(n565), .B(n564), .ZN(n645) );
  NAND2_X1 U683 ( .A1(G214), .A2(n566), .ZN(n712) );
  NOR2_X1 U684 ( .A1(G898), .A2(n471), .ZN(n567) );
  XOR2_X1 U685 ( .A(KEYINPUT95), .B(n567), .Z(n764) );
  NAND2_X1 U686 ( .A1(n764), .A2(G902), .ZN(n568) );
  NAND2_X1 U687 ( .A1(G952), .A2(n471), .ZN(n625) );
  AND2_X1 U688 ( .A1(n568), .A2(n625), .ZN(n570) );
  XNOR2_X1 U689 ( .A(KEYINPUT14), .B(n569), .ZN(n627) );
  INV_X1 U690 ( .A(n627), .ZN(n729) );
  NOR2_X1 U691 ( .A1(n570), .A2(n729), .ZN(n571) );
  INV_X1 U692 ( .A(n586), .ZN(n572) );
  XNOR2_X1 U693 ( .A(KEYINPUT72), .B(G469), .ZN(n576) );
  NAND2_X1 U694 ( .A1(n577), .A2(G234), .ZN(n578) );
  XNOR2_X1 U695 ( .A(n578), .B(KEYINPUT20), .ZN(n579) );
  XNOR2_X1 U696 ( .A(KEYINPUT98), .B(n579), .ZN(n581) );
  NAND2_X1 U697 ( .A1(n581), .A2(G221), .ZN(n580) );
  XOR2_X1 U698 ( .A(n580), .B(KEYINPUT21), .Z(n697) );
  XOR2_X1 U699 ( .A(KEYINPUT25), .B(KEYINPUT99), .Z(n583) );
  NAND2_X1 U700 ( .A1(G217), .A2(n581), .ZN(n582) );
  XOR2_X1 U701 ( .A(KEYINPUT24), .B(G110), .Z(n585) );
  INV_X1 U702 ( .A(n606), .ZN(n699) );
  NAND2_X1 U703 ( .A1(n589), .A2(G210), .ZN(n590) );
  XOR2_X1 U704 ( .A(KEYINPUT5), .B(G137), .Z(n592) );
  XNOR2_X1 U705 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U706 ( .A(n598), .B(KEYINPUT34), .ZN(n599) );
  AND2_X1 U707 ( .A1(n717), .A2(n697), .ZN(n601) );
  INV_X1 U708 ( .A(n666), .ZN(n615) );
  XOR2_X1 U709 ( .A(KEYINPUT100), .B(KEYINPUT31), .Z(n605) );
  NAND2_X1 U710 ( .A1(n708), .A2(n603), .ZN(n604) );
  XNOR2_X1 U711 ( .A(n605), .B(n604), .ZN(n687) );
  NOR2_X1 U712 ( .A1(n478), .A2(n607), .ZN(n608) );
  NAND2_X1 U713 ( .A1(n636), .A2(n608), .ZN(n670) );
  NAND2_X1 U714 ( .A1(n687), .A2(n670), .ZN(n613) );
  NAND2_X1 U715 ( .A1(n611), .A2(n610), .ZN(n686) );
  INV_X1 U716 ( .A(n686), .ZN(n676) );
  INV_X1 U717 ( .A(n650), .ZN(n612) );
  NAND2_X1 U718 ( .A1(n613), .A2(n612), .ZN(n614) );
  AND2_X1 U719 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U720 ( .A1(n478), .A2(n696), .ZN(n617) );
  NAND2_X1 U721 ( .A1(n618), .A2(n617), .ZN(n675) );
  XOR2_X1 U722 ( .A(KEYINPUT32), .B(KEYINPUT65), .Z(n620) );
  INV_X1 U723 ( .A(KEYINPUT77), .ZN(n661) );
  INV_X1 U724 ( .A(n623), .ZN(n629) );
  NOR2_X1 U725 ( .A1(G900), .A2(n471), .ZN(n624) );
  NAND2_X1 U726 ( .A1(n624), .A2(G902), .ZN(n626) );
  NAND2_X1 U727 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U728 ( .A1(n628), .A2(n627), .ZN(n638) );
  NAND2_X1 U729 ( .A1(n629), .A2(n640), .ZN(n630) );
  NAND2_X1 U730 ( .A1(n652), .A2(n712), .ZN(n631) );
  NOR2_X1 U731 ( .A1(n700), .A2(n631), .ZN(n632) );
  XNOR2_X1 U732 ( .A(n632), .B(KEYINPUT43), .ZN(n633) );
  NOR2_X1 U733 ( .A1(n485), .A2(n633), .ZN(n694) );
  NAND2_X1 U734 ( .A1(n706), .A2(n712), .ZN(n635) );
  NOR2_X2 U735 ( .A1(n660), .A2(n684), .ZN(n639) );
  AND2_X1 U736 ( .A1(n706), .A2(n640), .ZN(n641) );
  XNOR2_X1 U737 ( .A(KEYINPUT46), .B(KEYINPUT91), .ZN(n644) );
  NAND2_X1 U738 ( .A1(n714), .A2(KEYINPUT47), .ZN(n647) );
  NAND2_X1 U739 ( .A1(n682), .A2(n650), .ZN(n651) );
  INV_X1 U740 ( .A(n652), .ZN(n653) );
  NAND2_X1 U741 ( .A1(n700), .A2(n657), .ZN(n691) );
  OR2_X1 U742 ( .A1(n686), .A2(n660), .ZN(n693) );
  NAND2_X1 U743 ( .A1(n750), .A2(G472), .ZN(n665) );
  XOR2_X1 U744 ( .A(n666), .B(G101), .Z(G3) );
  NOR2_X1 U745 ( .A1(n684), .A2(n670), .ZN(n667) );
  XOR2_X1 U746 ( .A(G104), .B(n667), .Z(G6) );
  XOR2_X1 U747 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n669) );
  XNOR2_X1 U748 ( .A(KEYINPUT109), .B(KEYINPUT27), .ZN(n668) );
  XNOR2_X1 U749 ( .A(n669), .B(n668), .ZN(n674) );
  NOR2_X1 U750 ( .A1(n686), .A2(n670), .ZN(n672) );
  XNOR2_X1 U751 ( .A(G107), .B(KEYINPUT26), .ZN(n671) );
  XNOR2_X1 U752 ( .A(n672), .B(n671), .ZN(n673) );
  XOR2_X1 U753 ( .A(n674), .B(n673), .Z(G9) );
  XNOR2_X1 U754 ( .A(G110), .B(n675), .ZN(G12) );
  XOR2_X1 U755 ( .A(G128), .B(KEYINPUT29), .Z(n678) );
  NAND2_X1 U756 ( .A1(n682), .A2(n676), .ZN(n677) );
  XNOR2_X1 U757 ( .A(n678), .B(n677), .ZN(G30) );
  XNOR2_X1 U758 ( .A(n356), .B(KEYINPUT112), .ZN(n680) );
  XNOR2_X1 U759 ( .A(n680), .B(n679), .ZN(G45) );
  NAND2_X1 U760 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U761 ( .A(n683), .B(G146), .ZN(G48) );
  NOR2_X1 U762 ( .A1(n687), .A2(n684), .ZN(n685) );
  XOR2_X1 U763 ( .A(G113), .B(n685), .Z(G15) );
  NOR2_X1 U764 ( .A1(n687), .A2(n686), .ZN(n689) );
  XNOR2_X1 U765 ( .A(G116), .B(KEYINPUT113), .ZN(n688) );
  XNOR2_X1 U766 ( .A(n689), .B(n688), .ZN(G18) );
  XOR2_X1 U767 ( .A(KEYINPUT37), .B(KEYINPUT114), .Z(n690) );
  XNOR2_X1 U768 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U769 ( .A(G125), .B(n692), .ZN(G27) );
  XNOR2_X1 U770 ( .A(G134), .B(n693), .ZN(G36) );
  XNOR2_X1 U771 ( .A(G140), .B(n694), .ZN(n695) );
  XNOR2_X1 U772 ( .A(n695), .B(KEYINPUT115), .ZN(G42) );
  OR2_X1 U773 ( .A1(n711), .A2(n723), .ZN(n737) );
  NOR2_X1 U774 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U775 ( .A(KEYINPUT49), .B(n698), .ZN(n704) );
  XOR2_X1 U776 ( .A(KEYINPUT50), .B(n701), .Z(n702) );
  XNOR2_X1 U777 ( .A(KEYINPUT116), .B(n702), .ZN(n703) );
  NAND2_X1 U778 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U779 ( .A1(n478), .A2(n705), .ZN(n707) );
  NOR2_X1 U780 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U781 ( .A(KEYINPUT51), .B(n709), .Z(n710) );
  NOR2_X1 U782 ( .A1(n711), .A2(n710), .ZN(n725) );
  INV_X1 U783 ( .A(n712), .ZN(n719) );
  INV_X1 U784 ( .A(n713), .ZN(n715) );
  NOR2_X1 U785 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U786 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U787 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U788 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U789 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U790 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U791 ( .A(n726), .B(KEYINPUT52), .Z(n727) );
  XNOR2_X1 U792 ( .A(KEYINPUT117), .B(n727), .ZN(n728) );
  NOR2_X1 U793 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U794 ( .A1(n730), .A2(G952), .ZN(n731) );
  XNOR2_X1 U795 ( .A(n731), .B(KEYINPUT118), .ZN(n732) );
  NAND2_X1 U796 ( .A1(n732), .A2(n471), .ZN(n735) );
  NOR2_X1 U797 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U798 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U799 ( .A(n738), .B(KEYINPUT53), .ZN(n739) );
  XNOR2_X1 U800 ( .A(KEYINPUT119), .B(n739), .ZN(G75) );
  XOR2_X1 U801 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n741) );
  XNOR2_X1 U802 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n745) );
  XNOR2_X1 U803 ( .A(n743), .B(KEYINPUT57), .ZN(n744) );
  NAND2_X1 U804 ( .A1(n750), .A2(G475), .ZN(n749) );
  INV_X1 U805 ( .A(KEYINPUT59), .ZN(n747) );
  NAND2_X1 U806 ( .A1(n750), .A2(G478), .ZN(n752) );
  NAND2_X1 U807 ( .A1(G217), .A2(n750), .ZN(n753) );
  XNOR2_X1 U808 ( .A(n754), .B(n753), .ZN(n755) );
  NOR2_X1 U809 ( .A1(n756), .A2(n755), .ZN(G66) );
  OR2_X1 U810 ( .A1(n757), .A2(G953), .ZN(n761) );
  NAND2_X1 U811 ( .A1(G953), .A2(G224), .ZN(n758) );
  XNOR2_X1 U812 ( .A(KEYINPUT61), .B(n758), .ZN(n759) );
  NAND2_X1 U813 ( .A1(n759), .A2(G898), .ZN(n760) );
  NAND2_X1 U814 ( .A1(n761), .A2(n760), .ZN(n766) );
  XNOR2_X1 U815 ( .A(G110), .B(n762), .ZN(n763) );
  NOR2_X1 U816 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U817 ( .A(n766), .B(n765), .ZN(G69) );
  XOR2_X1 U818 ( .A(KEYINPUT124), .B(n767), .Z(n771) );
  XNOR2_X1 U819 ( .A(n768), .B(n769), .ZN(n770) );
  XNOR2_X1 U820 ( .A(n771), .B(n770), .ZN(n772) );
  XOR2_X1 U821 ( .A(n773), .B(n772), .Z(n778) );
  XNOR2_X1 U822 ( .A(KEYINPUT125), .B(n778), .ZN(n775) );
  XOR2_X1 U823 ( .A(n775), .B(n774), .Z(n777) );
  NAND2_X1 U824 ( .A1(n777), .A2(n471), .ZN(n782) );
  XNOR2_X1 U825 ( .A(G227), .B(n778), .ZN(n779) );
  NAND2_X1 U826 ( .A1(n779), .A2(G900), .ZN(n780) );
  NAND2_X1 U827 ( .A1(n780), .A2(G953), .ZN(n781) );
  NAND2_X1 U828 ( .A1(n782), .A2(n781), .ZN(G72) );
  XOR2_X1 U829 ( .A(n783), .B(G119), .Z(n784) );
  XNOR2_X1 U830 ( .A(KEYINPUT127), .B(n784), .ZN(G21) );
  XOR2_X1 U831 ( .A(n785), .B(G137), .Z(G39) );
endmodule

