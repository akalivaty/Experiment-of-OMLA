//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT67), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT68), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT69), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT70), .Z(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n466), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n477), .A2(new_n467), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  OAI211_X1 g060(.A(G138), .B(new_n467), .C1(new_n475), .C2(new_n476), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n488), .A2(new_n467), .A3(G138), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT71), .B1(new_n477), .B2(new_n489), .ZN(new_n490));
  AND3_X1   g065(.A1(new_n488), .A2(new_n467), .A3(G138), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n466), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n487), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n480), .B2(G126), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n494), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n495), .B1(new_n494), .B2(new_n499), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(G164));
  OR2_X1    g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n512), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n513), .A2(new_n514), .B1(G651), .B2(new_n520), .ZN(G166));
  NAND3_X1  g096(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT74), .Z(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  OR2_X1    g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT75), .B(G89), .Z(new_n531));
  OAI211_X1 g106(.A(new_n528), .B(new_n530), .C1(new_n507), .C2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n523), .A2(new_n532), .ZN(G168));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n518), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT76), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n534), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n539), .B1(new_n538), .B2(new_n537), .ZN(new_n540));
  INV_X1    g115(.A(new_n507), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n541), .A2(G90), .B1(new_n527), .B2(G52), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  AOI22_X1  g119(.A1(new_n541), .A2(G81), .B1(new_n527), .B2(G43), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n534), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(new_n507), .A2(KEYINPUT78), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT78), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n505), .A2(new_n506), .A3(new_n555), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G91), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n559));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n509), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n527), .A2(KEYINPUT77), .A3(G53), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n561), .A2(KEYINPUT9), .A3(new_n562), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n565), .A2(new_n534), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n558), .A2(new_n563), .A3(new_n564), .A4(new_n566), .ZN(G299));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  NAND3_X1  g144(.A1(new_n554), .A2(G87), .A3(new_n556), .ZN(new_n570));
  INV_X1    g145(.A(G74), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n534), .B1(new_n518), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(G49), .B2(new_n527), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(G288));
  INV_X1    g149(.A(KEYINPUT79), .ZN(new_n575));
  INV_X1    g150(.A(G73), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n576), .B2(new_n524), .ZN(new_n577));
  NAND3_X1  g152(.A1(KEYINPUT79), .A2(G73), .A3(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n577), .B(new_n578), .C1(new_n518), .C2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(new_n527), .B2(G48), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n554), .A2(G86), .A3(new_n556), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n534), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  INV_X1    g161(.A(G47), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n507), .A2(new_n586), .B1(new_n509), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n505), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G54), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n592), .A2(new_n534), .B1(new_n593), .B2(new_n509), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n557), .A2(G92), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n557), .A2(KEYINPUT10), .A3(G92), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n591), .B1(new_n599), .B2(G868), .ZN(G284));
  XOR2_X1   g175(.A(G284), .B(KEYINPUT80), .Z(G321));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NOR2_X1   g177(.A1(G168), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT81), .ZN(new_n604));
  INV_X1    g179(.A(G299), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n605), .A2(KEYINPUT82), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n602), .B1(new_n605), .B2(KEYINPUT82), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(G297));
  OAI21_X1  g183(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n599), .B1(new_n610), .B2(G860), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT83), .ZN(G148));
  OAI21_X1  g187(.A(KEYINPUT84), .B1(new_n548), .B2(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n599), .A2(new_n610), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  MUX2_X1   g190(.A(KEYINPUT84), .B(new_n613), .S(new_n615), .Z(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n466), .A2(new_n464), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  INV_X1    g195(.A(G2100), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  AOI22_X1  g198(.A1(G123), .A2(new_n480), .B1(new_n478), .B2(G135), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n467), .A2(G111), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n463), .B1(new_n625), .B2(KEYINPUT85), .ZN(new_n626));
  OAI21_X1  g201(.A(KEYINPUT85), .B1(G99), .B2(G2105), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n626), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(G2096), .Z(new_n631));
  NAND3_X1  g206(.A1(new_n622), .A2(new_n623), .A3(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  INV_X1    g208(.A(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G2427), .B(G2430), .Z(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT86), .B(KEYINPUT14), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n635), .A2(new_n636), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT87), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(G14), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n645), .B2(new_n646), .ZN(new_n651));
  AND2_X1   g226(.A1(new_n649), .A2(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT17), .Z(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  INV_X1    g233(.A(new_n655), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(new_n653), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n657), .B(new_n658), .C1(new_n656), .C2(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n653), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2096), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT88), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(KEYINPUT90), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  OR3_X1    g249(.A1(new_n668), .A2(new_n669), .A3(KEYINPUT90), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n674), .A2(new_n668), .A3(new_n669), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n668), .B(new_n669), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n677), .B(new_n678), .C1(new_n674), .C2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1991), .B(G1996), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G229));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  NOR2_X1   g263(.A1(G162), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n688), .B2(G35), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n691));
  INV_X1    g266(.A(G2090), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G2084), .ZN(new_n695));
  NAND2_X1  g270(.A1(G160), .A2(G29), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT24), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n697), .A2(G34), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n688), .B1(new_n697), .B2(G34), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n694), .B1(new_n695), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n695), .B2(new_n700), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n688), .A2(G26), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n478), .A2(G140), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n480), .A2(G128), .ZN(new_n706));
  OR2_X1    g281(.A1(G104), .A2(G2105), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n707), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n704), .B1(new_n710), .B2(new_n688), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G2067), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G21), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G168), .B2(new_n713), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1966), .ZN(new_n716));
  NOR2_X1   g291(.A1(G16), .A2(G19), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n548), .B2(G16), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT93), .B(G1341), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT30), .B(G28), .ZN(new_n721));
  OR2_X1    g296(.A1(KEYINPUT31), .A2(G11), .ZN(new_n722));
  NAND2_X1  g297(.A1(KEYINPUT31), .A2(G11), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n721), .A2(new_n688), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n630), .B2(new_n688), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n690), .B2(new_n693), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  NOR4_X1   g302(.A1(new_n702), .A2(new_n712), .A3(new_n716), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n688), .A2(G27), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G164), .B2(new_n688), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(G2078), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n688), .A2(G32), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n478), .A2(G141), .B1(G105), .B2(new_n464), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n480), .A2(G129), .ZN(new_n734));
  NAND3_X1  g309(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT26), .Z(new_n736));
  NAND3_X1  g311(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT97), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n732), .B1(new_n742), .B2(new_n688), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT27), .B(G1996), .Z(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G2078), .B2(new_n730), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n713), .A2(G5), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G171), .B2(new_n713), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1961), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT25), .Z(new_n751));
  INV_X1    g326(.A(G139), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(new_n468), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT94), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(new_n467), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT95), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  MUX2_X1   g333(.A(G33), .B(new_n758), .S(G29), .Z(new_n759));
  AOI21_X1  g334(.A(new_n749), .B1(G2072), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n728), .A2(new_n731), .A3(new_n746), .A4(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n759), .A2(G2072), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT96), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n713), .A2(G4), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n599), .B2(new_n713), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1348), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n713), .A2(G20), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT23), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n605), .B2(new_n713), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1956), .ZN(new_n770));
  NOR4_X1   g345(.A1(new_n761), .A2(new_n763), .A3(new_n766), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(G166), .A2(G16), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G16), .B2(G22), .ZN(new_n773));
  INV_X1    g348(.A(G1971), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n713), .A2(G23), .ZN(new_n776));
  INV_X1    g351(.A(G288), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(new_n713), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT33), .B(G1976), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G6), .B(G305), .S(G16), .Z(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT32), .B(G1981), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n781), .B(new_n782), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n773), .A2(new_n774), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n775), .A2(new_n780), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(KEYINPUT34), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(KEYINPUT34), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n688), .A2(G25), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n480), .A2(G119), .ZN(new_n789));
  INV_X1    g364(.A(G131), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n468), .ZN(new_n791));
  OR2_X1    g366(.A1(G95), .A2(G2105), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n792), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT91), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n788), .B1(new_n795), .B2(new_n688), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT35), .B(G1991), .Z(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n796), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n589), .A2(G16), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G16), .B2(G24), .ZN(new_n801));
  INV_X1    g376(.A(G1986), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(KEYINPUT92), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n801), .A2(new_n802), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n799), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n786), .A2(new_n787), .A3(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT36), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n771), .A2(new_n809), .A3(new_n810), .ZN(G150));
  XOR2_X1   g386(.A(G150), .B(KEYINPUT99), .Z(G311));
  NAND2_X1  g387(.A1(new_n599), .A2(G559), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT102), .B(G93), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n541), .A2(new_n816), .B1(new_n527), .B2(G55), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  OAI21_X1  g393(.A(KEYINPUT101), .B1(new_n818), .B2(new_n534), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n818), .A2(KEYINPUT101), .A3(new_n534), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(new_n548), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n815), .B(new_n823), .Z(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(KEYINPUT39), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT103), .ZN(new_n826));
  AOI21_X1  g401(.A(G860), .B1(new_n824), .B2(KEYINPUT39), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(G860), .B1(new_n820), .B2(new_n821), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT37), .Z(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(G145));
  NAND2_X1  g406(.A1(new_n494), .A2(new_n499), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT104), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n758), .B(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n795), .B(new_n619), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n741), .B(new_n709), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n480), .A2(G130), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n467), .A2(G118), .ZN(new_n839));
  OAI21_X1  g414(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(G142), .B2(new_n478), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n837), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n836), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n630), .B(G160), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G162), .ZN(new_n846));
  AOI21_X1  g421(.A(G37), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n846), .B2(new_n844), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g424(.A(new_n823), .B(new_n614), .Z(new_n850));
  INV_X1    g425(.A(KEYINPUT105), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n599), .B(new_n605), .ZN(new_n852));
  OR3_X1    g427(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(KEYINPUT41), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n850), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT42), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n858), .A2(KEYINPUT106), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(G166), .B(new_n777), .ZN(new_n861));
  XNOR2_X1  g436(.A(G305), .B(new_n589), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(KEYINPUT106), .B2(new_n858), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n857), .A2(new_n859), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n860), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n864), .B1(new_n860), .B2(new_n865), .ZN(new_n867));
  OAI21_X1  g442(.A(G868), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(G868), .B2(new_n822), .ZN(G295));
  OAI21_X1  g444(.A(new_n868), .B1(G868), .B2(new_n822), .ZN(G331));
  NAND2_X1  g445(.A1(G301), .A2(KEYINPUT107), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n823), .B(new_n871), .Z(new_n872));
  OAI21_X1  g447(.A(G168), .B1(G301), .B2(KEYINPUT107), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n823), .B(new_n871), .ZN(new_n875));
  INV_X1    g450(.A(new_n873), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n854), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT108), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n874), .A2(new_n852), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n863), .ZN(new_n883));
  AOI21_X1  g458(.A(G37), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n880), .A2(new_n863), .A3(new_n881), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n885), .B1(new_n884), .B2(new_n886), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n889));
  OAI22_X1  g464(.A1(new_n887), .A2(new_n888), .B1(KEYINPUT109), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n884), .A2(new_n886), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT43), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n893));
  XOR2_X1   g468(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n890), .A2(new_n895), .ZN(G397));
  AOI22_X1  g471(.A1(new_n478), .A2(G137), .B1(G101), .B2(new_n464), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n471), .A2(new_n472), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n897), .B(G40), .C1(new_n467), .C2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(G1384), .B1(new_n494), .B2(new_n499), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT45), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n709), .B(G2067), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n901), .B1(new_n741), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n901), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n904), .A2(G1996), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n905), .B2(KEYINPUT46), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n906), .B1(KEYINPUT46), .B2(new_n905), .ZN(new_n907));
  XNOR2_X1  g482(.A(KEYINPUT124), .B(KEYINPUT47), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n907), .B(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n909), .A2(KEYINPUT125), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(KEYINPUT125), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n742), .A2(G1996), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n742), .A2(G1996), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n902), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n795), .A2(new_n797), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n791), .A2(new_n794), .A3(new_n798), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(new_n904), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n901), .A2(new_n802), .A3(new_n589), .ZN(new_n921));
  XOR2_X1   g496(.A(new_n921), .B(KEYINPUT48), .Z(new_n922));
  NOR2_X1   g497(.A1(new_n709), .A2(G2067), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n914), .B2(new_n916), .ZN(new_n924));
  OAI22_X1  g499(.A1(new_n920), .A2(new_n922), .B1(new_n904), .B2(new_n924), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n910), .A2(new_n911), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G40), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n470), .A2(new_n473), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n900), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(G8), .ZN(new_n930));
  INV_X1    g505(.A(G1981), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n581), .A2(new_n582), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n577), .A2(new_n578), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n579), .B1(new_n503), .B2(new_n504), .ZN(new_n934));
  OAI21_X1  g509(.A(G651), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n527), .A2(G48), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n505), .A2(new_n506), .A3(G86), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(G1981), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT49), .B1(new_n932), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n930), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n932), .A2(new_n939), .A3(KEYINPUT49), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n942), .A2(KEYINPUT113), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(KEYINPUT113), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G1976), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n946), .A3(new_n777), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n930), .B1(new_n947), .B2(new_n932), .ZN(new_n948));
  XNOR2_X1  g523(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n949));
  NAND3_X1  g524(.A1(G303), .A2(G8), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n949), .ZN(new_n951));
  INV_X1    g526(.A(G8), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(G166), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n900), .A2(KEYINPUT45), .ZN(new_n955));
  INV_X1    g530(.A(G1384), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(new_n500), .B2(new_n501), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(G1971), .B1(new_n959), .B2(new_n928), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n899), .B1(new_n900), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n832), .A2(KEYINPUT72), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n494), .A2(new_n499), .A3(new_n495), .ZN(new_n964));
  AOI21_X1  g539(.A(G1384), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n692), .B(new_n962), .C1(new_n965), .C2(new_n961), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  OAI211_X1 g542(.A(G8), .B(new_n954), .C1(new_n960), .C2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n952), .B1(new_n928), .B2(new_n900), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT52), .B1(G288), .B2(new_n946), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n570), .A2(new_n573), .A3(G1976), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT112), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n970), .A2(new_n971), .A3(new_n975), .A4(new_n972), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n929), .A2(G8), .A3(new_n972), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT111), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n970), .A2(new_n980), .A3(new_n972), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n979), .A2(new_n981), .A3(KEYINPUT52), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n977), .A2(new_n982), .A3(new_n945), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n948), .B1(new_n969), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n954), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n900), .A2(KEYINPUT45), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n986), .B(new_n928), .C1(new_n965), .C2(KEYINPUT45), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n928), .B1(new_n900), .B2(new_n961), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n965), .B2(new_n961), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n987), .A2(new_n774), .B1(new_n989), .B2(new_n692), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n985), .B1(new_n990), .B2(new_n952), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n832), .A2(new_n956), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n899), .B1(new_n992), .B2(new_n958), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n957), .B2(new_n958), .ZN(new_n994));
  INV_X1    g569(.A(G1966), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n695), .B(new_n962), .C1(new_n965), .C2(new_n961), .ZN(new_n997));
  AOI211_X1 g572(.A(new_n952), .B(G286), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n991), .A2(new_n983), .A3(new_n998), .A4(new_n968), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT63), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n928), .B1(new_n992), .B2(KEYINPUT50), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(KEYINPUT50), .B2(new_n957), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n1003), .A2(new_n695), .B1(new_n994), .B2(new_n995), .ZN(new_n1004));
  NOR4_X1   g579(.A1(new_n1004), .A2(new_n1000), .A3(new_n952), .A4(G286), .ZN(new_n1005));
  OAI21_X1  g580(.A(G8), .B1(new_n960), .B2(new_n967), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n985), .ZN(new_n1007));
  AND4_X1   g582(.A1(new_n968), .A2(new_n1005), .A3(new_n983), .A4(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n984), .B1(new_n1001), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n996), .A2(G168), .A3(new_n997), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(new_n952), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT51), .ZN(new_n1014));
  AOI21_X1  g589(.A(G168), .B1(new_n996), .B2(new_n997), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1011), .A2(KEYINPUT51), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n1010), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1014), .B1(new_n1017), .B2(new_n952), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT122), .B1(new_n1018), .B2(KEYINPUT62), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n991), .A2(new_n968), .A3(new_n983), .ZN(new_n1020));
  INV_X1    g595(.A(G1961), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n962), .B1(new_n965), .B2(new_n961), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n928), .B1(new_n900), .B2(KEYINPUT45), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n965), .B2(KEYINPUT45), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(G2078), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1021), .A2(new_n1022), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1025), .B1(new_n987), .B2(G2078), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(G171), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1020), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT62), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1032), .B(new_n1014), .C1(new_n1017), .C2(new_n952), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1019), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1018), .A2(KEYINPUT122), .A3(KEYINPUT62), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1009), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1016), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1038), .B1(new_n1004), .B2(G168), .ZN(new_n1039));
  OAI21_X1  g614(.A(G8), .B1(new_n1039), .B2(new_n1015), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1020), .B1(new_n1040), .B2(new_n1014), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT120), .B1(new_n1003), .B2(G1961), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1022), .A2(new_n1043), .A3(new_n1021), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n993), .A2(new_n986), .A3(new_n1026), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1042), .A2(new_n1028), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1030), .B1(G171), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1048), .B1(new_n1046), .B2(G171), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1027), .A2(G301), .A3(new_n1028), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT121), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1050), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1041), .A2(new_n1049), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT61), .ZN(new_n1057));
  XOR2_X1   g632(.A(G299), .B(KEYINPUT57), .Z(new_n1058));
  INV_X1    g633(.A(new_n988), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(new_n957), .B2(KEYINPUT50), .ZN(new_n1060));
  INV_X1    g635(.A(G1956), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT56), .B(G2072), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n959), .A2(new_n928), .A3(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1058), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1058), .B1(new_n1064), .B2(new_n1062), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1057), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n929), .A2(G2067), .ZN(new_n1069));
  INV_X1    g644(.A(G1348), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1069), .B1(new_n1022), .B2(new_n1070), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n597), .A2(new_n598), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1071), .A2(new_n1072), .A3(new_n594), .ZN(new_n1073));
  AOI211_X1 g648(.A(new_n599), .B(new_n1069), .C1(new_n1022), .C2(new_n1070), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT60), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1076));
  XNOR2_X1  g651(.A(G299), .B(KEYINPUT57), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1078), .A2(KEYINPUT61), .A3(new_n1065), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT60), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1071), .A2(new_n1080), .A3(new_n599), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1068), .A2(new_n1075), .A3(new_n1079), .A4(new_n1081), .ZN(new_n1082));
  OR2_X1    g657(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT58), .B(G1341), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(new_n928), .B2(new_n900), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n899), .A2(G1996), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n986), .B(new_n1086), .C1(new_n965), .C2(KEYINPUT45), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n957), .A2(new_n958), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1090), .A2(KEYINPUT115), .A3(new_n986), .A4(new_n1086), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1085), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n548), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI211_X1 g669(.A(KEYINPUT116), .B(new_n1085), .C1(new_n1089), .C2(new_n1091), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1083), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1097));
  XOR2_X1   g672(.A(new_n1097), .B(KEYINPUT118), .Z(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1083), .B(new_n1098), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1082), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1065), .B1(new_n1073), .B2(new_n1067), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1103), .B(KEYINPUT114), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1056), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1037), .A2(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n589), .B(G1986), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n904), .B1(new_n919), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT123), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n1111));
  AOI211_X1 g686(.A(new_n1111), .B(new_n1108), .C1(new_n1037), .C2(new_n1105), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n926), .B1(new_n1110), .B2(new_n1112), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g688(.A1(G227), .A2(new_n461), .ZN(new_n1115));
  AOI21_X1  g689(.A(new_n1115), .B1(new_n649), .B2(new_n651), .ZN(new_n1116));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n1117));
  AND3_X1   g691(.A1(new_n1116), .A2(new_n686), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g692(.A(new_n1117), .B1(new_n1116), .B2(new_n686), .ZN(new_n1119));
  OAI21_X1  g693(.A(new_n848), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g694(.A(new_n1120), .B1(new_n892), .B2(new_n893), .ZN(G308));
  OAI221_X1 g695(.A(new_n848), .B1(new_n1118), .B2(new_n1119), .C1(new_n887), .C2(new_n888), .ZN(G225));
endmodule


