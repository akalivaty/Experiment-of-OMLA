//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT0), .Z(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT65), .B(G68), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n212), .B1(G238), .B2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT66), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(new_n214), .A2(new_n215), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G87), .A2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G58), .A2(G232), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(G97), .A2(G257), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n205), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n227), .A2(G50), .A3(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n208), .B(new_n223), .C1(new_n226), .C2(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT68), .B(KEYINPUT69), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n236), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT70), .B(G107), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(G33), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n252), .A2(new_n253), .A3(new_n224), .A4(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G97), .ZN(new_n256));
  INV_X1    g0056(.A(G97), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  AND3_X1   g0058(.A1(new_n256), .A2(KEYINPUT83), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(KEYINPUT83), .B1(new_n256), .B2(new_n258), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(new_n225), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT7), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n264), .A2(KEYINPUT7), .A3(new_n225), .A4(new_n265), .ZN(new_n269));
  AOI21_X1  g0069(.A(KEYINPUT79), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT79), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n271), .B1(new_n266), .B2(new_n267), .ZN(new_n272));
  OAI21_X1  g0072(.A(G107), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(G97), .B(G107), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT82), .A2(KEYINPUT6), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT6), .A2(G107), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n277), .B1(KEYINPUT82), .B2(KEYINPUT6), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n276), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G20), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G77), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n273), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n254), .A2(new_n224), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n261), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  AND2_X1   g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  OAI211_X1 g0088(.A(G244), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT4), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n264), .A2(new_n265), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n292), .A2(KEYINPUT4), .A3(G244), .A4(new_n286), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G283), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(G250), .A3(G1698), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n291), .A2(new_n293), .A3(new_n294), .A4(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G41), .ZN(new_n297));
  OAI211_X1 g0097(.A(G1), .B(G13), .C1(new_n263), .C2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(KEYINPUT5), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT5), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G41), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n251), .A2(G45), .ZN(new_n306));
  OAI211_X1 g0106(.A(G257), .B(new_n298), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G274), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(new_n302), .A3(new_n304), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n300), .A2(new_n301), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n311), .B1(new_n296), .B2(new_n299), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n313), .B1(G169), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT84), .B1(new_n285), .B2(new_n315), .ZN(new_n316));
  AOI211_X1 g0116(.A(G179), .B(new_n311), .C1(new_n296), .C2(new_n299), .ZN(new_n317));
  AOI21_X1  g0117(.A(G169), .B1(new_n300), .B2(new_n312), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G107), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n287), .A2(new_n288), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT7), .B1(new_n321), .B2(new_n225), .ZN(new_n322));
  INV_X1    g0122(.A(new_n269), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n271), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n272), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n320), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n280), .A2(new_n282), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n284), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n261), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT84), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n319), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n316), .A2(new_n332), .ZN(new_n333));
  OR2_X1    g0133(.A1(G238), .A2(G1698), .ZN(new_n334));
  OAI221_X1 g0134(.A(new_n334), .B1(G244), .B2(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G33), .A2(G116), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n298), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n298), .A2(G250), .A3(new_n306), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n337), .A2(new_n339), .A3(new_n309), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n301), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n263), .A2(G20), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT19), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n343), .A3(G97), .ZN(new_n344));
  NOR2_X1   g0144(.A1(G97), .A2(G107), .ZN(new_n345));
  INV_X1    g0145(.A(G87), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G97), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n345), .A2(new_n346), .B1(new_n347), .B2(new_n225), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n344), .B1(new_n348), .B2(new_n343), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n225), .B(G68), .C1(new_n287), .C2(new_n288), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT85), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n292), .A2(KEYINPUT85), .A3(new_n225), .A4(G68), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n349), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n284), .ZN(new_n355));
  INV_X1    g0155(.A(new_n255), .ZN(new_n356));
  XOR2_X1   g0156(.A(KEYINPUT15), .B(G87), .Z(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT15), .B(G87), .ZN(new_n359));
  INV_X1    g0159(.A(new_n252), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n355), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n309), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n264), .A2(new_n265), .B1(new_n211), .B2(G1698), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(new_n334), .B1(G33), .B2(G116), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n338), .B(new_n363), .C1(new_n365), .C2(new_n298), .ZN(new_n366));
  INV_X1    g0166(.A(G169), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n341), .A2(new_n362), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n366), .A2(G200), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n335), .A2(new_n336), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n299), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n372), .A2(G190), .A3(new_n338), .A4(new_n363), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n354), .A2(new_n284), .B1(new_n360), .B2(new_n359), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n356), .A2(G87), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n370), .A2(new_n373), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n369), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n314), .A2(G190), .ZN(new_n378));
  INV_X1    g0178(.A(G200), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n285), .B(new_n378), .C1(new_n379), .C2(new_n314), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n333), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  XNOR2_X1  g0181(.A(KEYINPUT8), .B(G58), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n360), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n284), .B1(new_n251), .B2(G20), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n384), .B1(new_n386), .B2(new_n383), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  XNOR2_X1  g0188(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n213), .B1(new_n270), .B2(new_n272), .ZN(new_n390));
  INV_X1    g0190(.A(G68), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT65), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT65), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G68), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G58), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n202), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(G20), .B1(G159), .B2(new_n281), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n389), .B1(new_n390), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(G68), .B1(new_n322), .B2(new_n323), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n400), .A3(KEYINPUT16), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n284), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n388), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n404), .A2(new_n308), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n298), .A2(new_n404), .ZN(new_n407));
  INV_X1    g0207(.A(G232), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI211_X1 g0209(.A(G226), .B(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT80), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT80), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n292), .A2(new_n412), .A3(G226), .A4(G1698), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n292), .A2(G223), .A3(new_n286), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G87), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n411), .A2(new_n413), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n409), .B1(new_n416), .B2(new_n299), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G179), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n367), .B2(new_n417), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n403), .A2(KEYINPUT18), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT18), .B1(new_n403), .B2(new_n419), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT81), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT18), .ZN(new_n423));
  INV_X1    g0223(.A(new_n389), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n395), .B1(new_n324), .B2(new_n325), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n201), .B1(new_n213), .B2(G58), .ZN(new_n426));
  INV_X1    g0226(.A(G159), .ZN(new_n427));
  INV_X1    g0227(.A(new_n281), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n426), .A2(new_n225), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n424), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n284), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n391), .B1(new_n268), .B2(new_n269), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n431), .B1(new_n433), .B2(KEYINPUT16), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n387), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  AOI211_X1 g0235(.A(new_n301), .B(new_n409), .C1(new_n416), .C2(new_n299), .ZN(new_n436));
  INV_X1    g0236(.A(new_n417), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n436), .B1(G169), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n423), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT81), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n403), .A2(KEYINPUT18), .A3(new_n419), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n430), .A2(new_n434), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n417), .A2(G190), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n437), .A2(G200), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n443), .A2(new_n444), .A3(new_n388), .A4(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT17), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n435), .A2(KEYINPUT17), .A3(new_n444), .A4(new_n445), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n422), .A2(new_n442), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n292), .A2(G238), .A3(G1698), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n292), .A2(G232), .A3(new_n286), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n452), .B(new_n453), .C1(new_n320), .C2(new_n292), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n405), .B1(new_n454), .B2(new_n299), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n211), .B2(new_n407), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G169), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(new_n301), .B2(new_n456), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n360), .A2(new_n210), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n385), .A2(G77), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n357), .A2(KEYINPUT71), .A3(new_n342), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT71), .ZN(new_n462));
  INV_X1    g0262(.A(new_n342), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n359), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  OAI22_X1  g0265(.A1(new_n382), .A2(new_n428), .B1(new_n225), .B2(new_n210), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n284), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT72), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n467), .A2(new_n468), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n459), .B(new_n460), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n458), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n471), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n456), .A2(G200), .ZN(new_n474));
  INV_X1    g0274(.A(G190), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(new_n456), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n451), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(G226), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n478));
  OAI211_X1 g0278(.A(G232), .B(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n478), .A2(new_n479), .A3(new_n347), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n299), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT74), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n407), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n405), .B1(new_n484), .B2(G238), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n480), .A2(KEYINPUT74), .A3(new_n299), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT13), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT75), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT13), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n483), .A2(new_n490), .A3(new_n485), .A4(new_n486), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  OR3_X1    g0292(.A1(new_n487), .A2(new_n489), .A3(KEYINPUT13), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G179), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n367), .B1(new_n488), .B2(new_n491), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT14), .ZN(new_n497));
  OR2_X1    g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n497), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n495), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n281), .A2(G50), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n501), .B(KEYINPUT76), .ZN(new_n502));
  OAI22_X1  g0302(.A1(new_n225), .A2(new_n213), .B1(new_n463), .B2(new_n210), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n284), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n504), .B(KEYINPUT11), .ZN(new_n505));
  XNOR2_X1  g0305(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n395), .B2(new_n360), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n386), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n252), .A2(KEYINPUT12), .ZN(new_n510));
  OAI221_X1 g0310(.A(new_n505), .B1(new_n391), .B2(new_n509), .C1(new_n507), .C2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n494), .B2(G190), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n488), .A2(new_n491), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G200), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n500), .A2(new_n511), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(G222), .A2(G1698), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n286), .A2(G223), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n292), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n518), .B(new_n299), .C1(G77), .C2(new_n292), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n484), .A2(G226), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n406), .A3(new_n520), .ZN(new_n521));
  OR2_X1    g0321(.A1(new_n521), .A2(G179), .ZN(new_n522));
  OAI21_X1  g0322(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n523));
  INV_X1    g0323(.A(G150), .ZN(new_n524));
  OAI221_X1 g0324(.A(new_n523), .B1(new_n524), .B2(new_n428), .C1(new_n463), .C2(new_n382), .ZN(new_n525));
  INV_X1    g0325(.A(G50), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n525), .A2(new_n284), .B1(new_n526), .B2(new_n360), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n385), .A2(G50), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n521), .A2(new_n367), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n522), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT9), .ZN(new_n533));
  OR2_X1    g0333(.A1(new_n533), .A2(KEYINPUT73), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(KEYINPUT73), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n529), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n527), .A2(KEYINPUT73), .A3(new_n533), .A4(new_n528), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n521), .A2(new_n475), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(G200), .B2(new_n521), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT10), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT10), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n538), .A2(new_n543), .A3(new_n540), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n532), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n515), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n477), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT95), .ZN(new_n548));
  INV_X1    g0348(.A(new_n310), .ZN(new_n549));
  OAI211_X1 g0349(.A(G250), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT93), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n292), .A2(KEYINPUT93), .A3(G250), .A4(new_n286), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G33), .A2(G294), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n292), .A2(G257), .A3(G1698), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n552), .A2(new_n553), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n549), .B1(new_n556), .B2(new_n299), .ZN(new_n557));
  OAI211_X1 g0357(.A(G264), .B(new_n298), .C1(new_n305), .C2(new_n306), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n558), .B(KEYINPUT94), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n557), .A2(G179), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n367), .B1(new_n557), .B2(new_n558), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n548), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OR3_X1    g0362(.A1(new_n336), .A2(KEYINPUT91), .A3(G20), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT91), .B1(new_n336), .B2(G20), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT23), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n225), .B2(G107), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n320), .A2(KEYINPUT23), .A3(G20), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n563), .A2(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n292), .A2(new_n225), .A3(G87), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n569), .A2(KEYINPUT22), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n569), .A2(KEYINPUT22), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n568), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT24), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(KEYINPUT24), .B(new_n568), .C1(new_n570), .C2(new_n571), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(new_n575), .A3(new_n284), .ZN(new_n576));
  OR3_X1    g0376(.A1(new_n252), .A2(KEYINPUT25), .A3(G107), .ZN(new_n577));
  OAI21_X1  g0377(.A(KEYINPUT25), .B1(new_n252), .B2(G107), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n577), .B(new_n578), .C1(new_n320), .C2(new_n255), .ZN(new_n579));
  XNOR2_X1  g0379(.A(new_n579), .B(KEYINPUT92), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n557), .A2(G179), .A3(new_n559), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n556), .A2(new_n299), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n583), .A2(new_n310), .A3(new_n558), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n582), .B(KEYINPUT95), .C1(new_n584), .C2(new_n367), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n562), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n557), .A2(new_n475), .A3(new_n558), .ZN(new_n587));
  AOI21_X1  g0387(.A(G200), .B1(new_n557), .B2(new_n559), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n576), .B(new_n580), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(G264), .B(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT87), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n292), .A2(KEYINPUT87), .A3(G264), .A4(G1698), .ZN(new_n594));
  XOR2_X1   g0394(.A(KEYINPUT88), .B(G303), .Z(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n321), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n292), .A2(G257), .A3(new_n286), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n593), .A2(new_n594), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n598), .A2(KEYINPUT89), .A3(new_n299), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(G270), .B(new_n298), .C1(new_n305), .C2(new_n306), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT86), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n601), .A2(new_n602), .A3(new_n310), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n602), .B1(new_n601), .B2(new_n310), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT89), .B1(new_n598), .B2(new_n299), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n600), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(G116), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n255), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n294), .B(new_n225), .C1(G33), .C2(new_n257), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n610), .B(new_n284), .C1(new_n225), .C2(G116), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT20), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n609), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n360), .A2(new_n608), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n607), .A2(KEYINPUT90), .A3(G179), .A4(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT90), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n598), .A2(new_n299), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT89), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n604), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n601), .A2(new_n602), .A3(new_n310), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n622), .A2(new_n625), .A3(G179), .A4(new_n599), .ZN(new_n626));
  INV_X1    g0426(.A(new_n617), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n619), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n622), .A2(new_n625), .A3(new_n599), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n367), .B1(new_n615), .B2(new_n616), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT21), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n631), .B1(new_n629), .B2(new_n630), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n618), .B(new_n628), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n607), .A2(new_n379), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n629), .A2(new_n475), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n635), .A2(new_n636), .A3(new_n617), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n381), .A2(new_n547), .A3(new_n590), .A4(new_n638), .ZN(G372));
  NAND2_X1  g0439(.A1(new_n439), .A2(new_n441), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n512), .A2(new_n514), .ZN(new_n641));
  INV_X1    g0441(.A(new_n511), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n496), .B(KEYINPUT14), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n642), .B1(new_n643), .B2(new_n495), .ZN(new_n644));
  INV_X1    g0444(.A(new_n472), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n448), .A2(new_n449), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n640), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n542), .A2(new_n544), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n532), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n547), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n581), .B1(new_n561), .B2(new_n560), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n634), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n333), .A2(new_n380), .A3(new_n377), .A4(new_n589), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT96), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n369), .B(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n316), .A2(new_n332), .A3(new_n377), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n658), .B1(new_n659), .B2(KEYINPUT26), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n285), .A2(new_n315), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n377), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n656), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n650), .B1(new_n651), .B2(new_n665), .ZN(G369));
  INV_X1    g0466(.A(G13), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G20), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n251), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n590), .A2(new_n634), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n653), .A2(new_n675), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n627), .A2(new_n675), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n634), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n634), .A2(new_n637), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n679), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n581), .A2(new_n674), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n562), .A2(new_n581), .A3(new_n585), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n590), .A2(new_n684), .B1(new_n685), .B2(new_n674), .ZN(new_n686));
  INV_X1    g0486(.A(new_n634), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n686), .B1(new_n687), .B2(new_n674), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n678), .B1(new_n683), .B2(new_n688), .ZN(new_n689));
  XOR2_X1   g0489(.A(new_n689), .B(KEYINPUT97), .Z(G399));
  INV_X1    g0490(.A(new_n206), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G41), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n345), .A2(new_n346), .A3(new_n608), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n693), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n229), .B2(new_n693), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n316), .A2(new_n332), .A3(new_n377), .A4(new_n662), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n377), .A2(new_n661), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n658), .B1(KEYINPUT26), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n634), .A2(new_n685), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n699), .B(new_n701), .C1(new_n702), .C2(new_n655), .ZN(new_n703));
  AND4_X1   g0503(.A1(KEYINPUT99), .A2(new_n703), .A3(KEYINPUT29), .A4(new_n675), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n675), .B1(new_n656), .B2(new_n664), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT29), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT99), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n703), .A2(KEYINPUT29), .A3(new_n675), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n704), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n314), .A2(new_n340), .A3(new_n559), .A4(new_n583), .ZN(new_n711));
  OR3_X1    g0511(.A1(new_n626), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(G179), .B1(new_n557), .B2(new_n559), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n300), .A2(new_n312), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n629), .A2(new_n366), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n710), .B1(new_n626), .B2(new_n711), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n712), .B(new_n715), .C1(KEYINPUT98), .C2(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n716), .A2(KEYINPUT98), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n674), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n381), .A2(new_n638), .A3(new_n590), .A4(new_n675), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n712), .A2(new_n716), .A3(new_n715), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G330), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n709), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n698), .B1(new_n728), .B2(G1), .ZN(G364));
  INV_X1    g0529(.A(new_n683), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n251), .B1(new_n668), .B2(G45), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n693), .A2(new_n731), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n682), .A2(G330), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n730), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  XOR2_X1   g0534(.A(new_n734), .B(KEYINPUT100), .Z(new_n735));
  NOR2_X1   g0535(.A1(G13), .A2(G33), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n682), .A2(G20), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n732), .B(KEYINPUT101), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n224), .B1(G20), .B2(new_n367), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n475), .A2(G20), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G179), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT103), .Z(new_n746));
  INV_X1    g0546(.A(G329), .ZN(new_n747));
  INV_X1    g0547(.A(G303), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n379), .A2(G179), .ZN(new_n749));
  NAND2_X1  g0549(.A1(G20), .A2(G190), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n746), .A2(new_n747), .B1(new_n748), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n301), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n751), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n753), .B1(G322), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n743), .A2(new_n749), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G283), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n225), .B1(new_n744), .B2(G190), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G294), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n742), .A2(new_n301), .A3(new_n379), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(KEYINPUT33), .B(G317), .Z(new_n766));
  NOR3_X1   g0566(.A1(new_n750), .A2(new_n301), .A3(new_n379), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G326), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n765), .A2(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n743), .A2(new_n754), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n292), .B(new_n770), .C1(G311), .C2(new_n772), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n757), .A2(new_n760), .A3(new_n763), .A4(new_n773), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n765), .A2(new_n391), .B1(new_n346), .B2(new_n752), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(G77), .B2(new_n772), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n745), .A2(new_n427), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT32), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n759), .A2(G107), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n762), .A2(G97), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n768), .A2(new_n526), .B1(new_n755), .B2(new_n396), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n321), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n776), .A2(new_n778), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n741), .B1(new_n774), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n737), .A2(G20), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n740), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n691), .A2(new_n292), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(new_n249), .B2(G45), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(G45), .B2(new_n229), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n691), .A2(new_n321), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT102), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G355), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n791), .B(new_n794), .C1(G116), .C2(new_n206), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n739), .B(new_n785), .C1(new_n787), .C2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT104), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n735), .B1(new_n738), .B2(new_n797), .ZN(G396));
  OAI21_X1  g0598(.A(KEYINPUT106), .B1(new_n473), .B2(new_n675), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT106), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n471), .A2(new_n800), .A3(new_n674), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n476), .A2(new_n799), .A3(new_n472), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(KEYINPUT107), .B1(new_n645), .B2(new_n674), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT107), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n472), .A2(new_n804), .A3(new_n675), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n802), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n705), .B(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(new_n726), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n732), .ZN(new_n809));
  INV_X1    g0609(.A(G311), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n321), .B1(new_n746), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G283), .B2(new_n764), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n758), .A2(new_n346), .ZN(new_n813));
  INV_X1    g0613(.A(G294), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n780), .B1(new_n320), .B2(new_n752), .C1(new_n814), .C2(new_n755), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n813), .B(new_n815), .C1(G303), .C2(new_n767), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n812), .B(new_n816), .C1(new_n608), .C2(new_n771), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT105), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n772), .A2(G159), .B1(new_n756), .B2(G143), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n767), .A2(G137), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n819), .B(new_n820), .C1(new_n524), .C2(new_n765), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT34), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n758), .A2(new_n391), .B1(new_n761), .B2(new_n396), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n321), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n822), .B(new_n824), .C1(new_n526), .C2(new_n752), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n746), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n740), .B1(new_n818), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n740), .A2(new_n736), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n739), .B1(new_n210), .B2(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n829), .B(new_n831), .C1(new_n806), .C2(new_n737), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n809), .A2(new_n832), .ZN(G384));
  INV_X1    g0633(.A(G330), .ZN(new_n834));
  OAI211_X1 g0634(.A(KEYINPUT31), .B(new_n674), .C1(new_n717), .C2(new_n718), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n721), .A2(new_n722), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n500), .A2(new_n511), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n511), .A2(new_n674), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n837), .A2(new_n641), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n644), .A2(new_n674), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n836), .A2(new_n841), .A3(new_n806), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT38), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n433), .A2(new_n389), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n388), .B1(new_n845), .B2(new_n402), .ZN(new_n846));
  INV_X1    g0646(.A(new_n672), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n420), .A2(new_n421), .A3(KEYINPUT81), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n440), .B1(new_n439), .B2(new_n441), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n647), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n848), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n403), .B1(new_n419), .B2(new_n847), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n854), .A2(new_n446), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n846), .B1(new_n419), .B2(new_n847), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n855), .B1(new_n857), .B2(new_n446), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n844), .B1(new_n853), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n848), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n859), .B1(new_n450), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT38), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT40), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n843), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n448), .B(new_n449), .C1(new_n420), .C2(new_n421), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n435), .A2(new_n672), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n854), .A2(new_n446), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n854), .A2(new_n446), .A3(new_n855), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT38), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(KEYINPUT38), .B2(new_n862), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT40), .B1(new_n842), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n834), .B1(new_n866), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n547), .A2(G330), .A3(new_n836), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n866), .A2(new_n876), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n547), .A2(new_n836), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n878), .A2(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n515), .A2(new_n838), .B1(new_n644), .B2(new_n674), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n806), .B(new_n675), .C1(new_n656), .C2(new_n664), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n472), .A2(new_n674), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n883), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n864), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n640), .B2(new_n847), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n644), .A2(new_n675), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n875), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n862), .A2(KEYINPUT38), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n844), .B(new_n859), .C1(new_n450), .C2(new_n861), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT39), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n890), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n889), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n882), .B(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n648), .A2(new_n649), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n531), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT99), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n660), .A2(new_n663), .ZN(new_n902));
  INV_X1    g0702(.A(new_n633), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n905), .A2(new_n628), .A3(new_n618), .A4(new_n652), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n381), .A2(new_n906), .A3(new_n589), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n674), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n901), .B(new_n708), .C1(new_n908), .C2(KEYINPUT29), .ZN(new_n909));
  INV_X1    g0709(.A(new_n704), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n900), .B1(new_n911), .B2(new_n547), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n898), .B(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n251), .B2(new_n668), .ZN(new_n914));
  OAI211_X1 g0714(.A(G116), .B(new_n226), .C1(new_n279), .C2(KEYINPUT35), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT108), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n279), .A2(KEYINPUT35), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT36), .ZN(new_n919));
  OAI21_X1  g0719(.A(G77), .B1(new_n395), .B2(new_n396), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n229), .A2(new_n920), .B1(G50), .B2(new_n391), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(G1), .A3(new_n667), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n914), .A2(new_n919), .A3(new_n922), .ZN(G367));
  NAND2_X1  g0723(.A1(new_n374), .A2(new_n375), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n658), .A2(new_n924), .A3(new_n674), .ZN(new_n925));
  INV_X1    g0725(.A(new_n924), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n377), .B1(new_n926), .B2(new_n675), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT43), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n333), .B(new_n380), .C1(new_n285), .C2(new_n675), .ZN(new_n933));
  OR3_X1    g0733(.A1(new_n676), .A2(KEYINPUT42), .A3(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT109), .Z(new_n935));
  NAND2_X1  g0735(.A1(new_n661), .A2(new_n674), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n333), .B1(new_n937), .B2(new_n586), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n675), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT42), .B1(new_n676), .B2(new_n933), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n931), .B(new_n932), .C1(new_n935), .C2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n683), .A2(new_n688), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(new_n937), .ZN(new_n944));
  INV_X1    g0744(.A(new_n941), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n934), .B(KEYINPUT109), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n945), .A2(new_n946), .A3(new_n930), .A4(new_n929), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n942), .A2(new_n944), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT110), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT111), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n678), .B(new_n937), .C1(new_n950), .C2(KEYINPUT44), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(KEYINPUT44), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n678), .A2(new_n937), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT45), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n953), .A2(new_n955), .A3(new_n943), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n683), .A2(new_n688), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n957), .A2(new_n943), .A3(new_n676), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n727), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n692), .B(KEYINPUT41), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n731), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n942), .A2(new_n947), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n962), .B1(new_n963), .B2(new_n944), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n949), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n739), .B1(new_n929), .B2(new_n786), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n787), .B1(new_n206), .B2(new_n359), .C1(new_n241), .C2(new_n789), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n772), .A2(G283), .B1(new_n767), .B2(G311), .ZN(new_n968));
  INV_X1    g0768(.A(new_n752), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(KEYINPUT46), .A3(G116), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT46), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n752), .B2(new_n608), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n970), .B(new_n972), .C1(new_n814), .C2(new_n765), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n968), .B1(new_n973), .B2(KEYINPUT112), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n759), .A2(G97), .ZN(new_n975));
  INV_X1    g0775(.A(G317), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n975), .B(new_n321), .C1(new_n976), .C2(new_n745), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT113), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n977), .A2(new_n978), .B1(G107), .B2(new_n762), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n973), .A2(KEYINPUT112), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n979), .B(new_n980), .C1(new_n978), .C2(new_n977), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n974), .B(new_n981), .C1(new_n595), .C2(new_n756), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n292), .B1(new_n758), .B2(new_n210), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT114), .ZN(new_n984));
  INV_X1    g0784(.A(new_n745), .ZN(new_n985));
  XNOR2_X1  g0785(.A(KEYINPUT115), .B(G137), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n985), .A2(new_n986), .B1(new_n764), .B2(G159), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G58), .A2(new_n969), .B1(new_n756), .B2(G150), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n762), .A2(G68), .B1(new_n767), .B2(G143), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n984), .A2(new_n987), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G50), .B2(new_n772), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n982), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT47), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n966), .B(new_n967), .C1(new_n993), .C2(new_n741), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n965), .A2(new_n994), .ZN(G387));
  INV_X1    g0795(.A(new_n731), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n958), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n686), .A2(new_n786), .ZN(new_n998));
  INV_X1    g0798(.A(new_n236), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n789), .B1(new_n999), .B2(G45), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n694), .B2(new_n793), .ZN(new_n1001));
  AOI21_X1  g0801(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n383), .A2(new_n526), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n695), .B(new_n1002), .C1(new_n1003), .C2(KEYINPUT50), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(KEYINPUT50), .B2(new_n1003), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n1001), .A2(new_n1005), .B1(G107), .B2(new_n206), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n739), .B1(new_n1006), .B2(new_n787), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n761), .A2(new_n359), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n391), .B2(new_n771), .C1(new_n524), .C2(new_n745), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n755), .A2(new_n526), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n765), .A2(new_n382), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n752), .A2(new_n210), .ZN(new_n1013));
  NOR4_X1   g0813(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n767), .A2(G159), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1014), .A2(new_n292), .A3(new_n975), .A4(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n772), .A2(new_n595), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n764), .A2(G311), .B1(new_n767), .B2(G322), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(new_n976), .C2(new_n755), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT48), .ZN(new_n1020));
  INV_X1    g0820(.A(G283), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1020), .B1(new_n1021), .B2(new_n761), .C1(new_n814), .C2(new_n752), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT49), .Z(new_n1023));
  OAI221_X1 g0823(.A(new_n321), .B1(new_n745), .B2(new_n769), .C1(new_n608), .C2(new_n758), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1016), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT116), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n998), .B(new_n1007), .C1(new_n1026), .C2(new_n741), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n728), .A2(new_n958), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n692), .B1(new_n728), .B2(new_n958), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n997), .B(new_n1027), .C1(new_n1028), .C2(new_n1029), .ZN(G393));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n956), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n953), .A2(new_n955), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(new_n943), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1031), .B(new_n692), .C1(new_n1028), .C2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n996), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n739), .B1(new_n937), .B2(new_n786), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n768), .A2(new_n524), .B1(new_n755), .B2(new_n427), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT51), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n761), .A2(new_n210), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n771), .A2(new_n382), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(G143), .C2(new_n985), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n526), .B2(new_n765), .C1(new_n395), .C2(new_n752), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n1043), .A2(new_n321), .A3(new_n813), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n756), .A2(G311), .B1(new_n767), .B2(G317), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT52), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n752), .A2(new_n1021), .B1(new_n761), .B2(new_n608), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n772), .A2(G294), .B1(new_n595), .B2(new_n764), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n292), .B1(new_n985), .B2(G322), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1048), .A2(new_n1049), .A3(new_n779), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n1046), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n740), .B1(new_n1044), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n246), .A2(new_n788), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1053), .B(new_n787), .C1(new_n257), .C2(new_n206), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT117), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1036), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1034), .A2(new_n1035), .A3(new_n1056), .ZN(G390));
  AOI21_X1  g0857(.A(new_n891), .B1(new_n860), .B2(new_n863), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n894), .A2(KEYINPUT39), .A3(new_n874), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n739), .B1(new_n1060), .B2(new_n736), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n830), .A2(new_n382), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n321), .B1(new_n746), .B2(new_n814), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1039), .B(new_n1063), .C1(G283), .C2(new_n767), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n756), .A2(G116), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n759), .A2(G68), .B1(new_n969), .B2(G87), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n772), .A2(G97), .B1(G107), .B2(new_n764), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(G125), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n746), .A2(new_n1069), .B1(new_n526), .B2(new_n758), .ZN(new_n1070));
  XOR2_X1   g0870(.A(KEYINPUT54), .B(G143), .Z(new_n1071));
  AOI211_X1 g0871(.A(new_n321), .B(new_n1070), .C1(new_n772), .C2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n752), .A2(new_n524), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT53), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n762), .A2(G159), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n756), .A2(G132), .B1(new_n764), .B2(new_n986), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(G128), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n768), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1068), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n740), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1061), .A2(new_n1062), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n890), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n892), .B(new_n895), .C1(new_n887), .C2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n890), .B1(new_n894), .B2(new_n874), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n703), .A2(new_n806), .A3(new_n675), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n883), .B1(new_n1086), .B2(new_n886), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n725), .A2(new_n841), .A3(G330), .A4(new_n806), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1084), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n885), .B1(new_n908), .B2(new_n806), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n890), .B1(new_n1092), .B2(new_n883), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1091), .B1(new_n1060), .B2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n836), .A2(new_n841), .A3(G330), .A4(new_n806), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1090), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1082), .B1(new_n1096), .B2(new_n731), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1084), .A2(new_n1088), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1095), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n725), .A2(G330), .A3(new_n806), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n883), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n1095), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1092), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n836), .A2(G330), .A3(new_n806), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n883), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1086), .A2(new_n886), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1107), .A2(new_n1089), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n650), .B(new_n879), .C1(new_n709), .C2(new_n651), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1100), .A2(new_n1090), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1109), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1092), .B1(new_n1102), .B2(new_n1095), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n912), .B(new_n879), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(KEYINPUT118), .B1(new_n1096), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1111), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1118), .A2(new_n1119), .A3(new_n1090), .A4(new_n1100), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1113), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1097), .B1(new_n1121), .B2(new_n692), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(G378));
  XNOR2_X1  g0923(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n544), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n543), .B1(new_n538), .B2(new_n540), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n531), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n529), .A2(new_n847), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n545), .A2(new_n1128), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1124), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1130), .A2(new_n1131), .A3(new_n1124), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(KEYINPUT119), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT119), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1134), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1136), .B1(new_n1137), .B2(new_n1132), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n736), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n755), .A2(new_n320), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n746), .A2(new_n1021), .ZN(new_n1142));
  NOR3_X1   g0942(.A1(new_n1142), .A2(G41), .A3(new_n292), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n759), .A2(G58), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(new_n359), .C2(new_n771), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1141), .B(new_n1145), .C1(G97), .C2(new_n764), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1013), .B1(G68), .B2(new_n762), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1146), .B(new_n1147), .C1(new_n608), .C2(new_n768), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT58), .Z(new_n1149));
  INV_X1    g0949(.A(G124), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n297), .B1(new_n745), .B2(new_n1150), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n768), .A2(new_n1069), .B1(new_n761), .B2(new_n524), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n772), .A2(G137), .B1(G132), .B2(new_n764), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n1078), .B2(new_n755), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1152), .B(new_n1154), .C1(new_n969), .C2(new_n1071), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT59), .ZN(new_n1156));
  AOI211_X1 g0956(.A(G33), .B(new_n1151), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n1156), .B2(new_n1155), .C1(new_n427), .C2(new_n758), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n526), .B1(new_n287), .B2(G41), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n740), .B1(new_n1149), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n732), .B1(new_n526), .B2(new_n830), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1140), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n897), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n877), .A2(new_n1166), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n834), .B(new_n1139), .C1(new_n866), .C2(new_n876), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1165), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n880), .A2(G330), .A3(new_n1135), .A4(new_n1138), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1170), .B(new_n897), .C1(new_n877), .C2(new_n1166), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1164), .B1(new_n1172), .B2(new_n996), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT57), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1111), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n692), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1169), .A2(new_n1171), .A3(KEYINPUT120), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT120), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n1181), .A3(new_n897), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n1183), .A2(new_n1175), .A3(new_n1174), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1173), .B1(new_n1178), .B2(new_n1184), .ZN(G375));
  OAI21_X1  g0985(.A(new_n996), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(KEYINPUT121), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT121), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1110), .A2(new_n1188), .A3(new_n996), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n739), .B1(new_n883), .B2(new_n736), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n830), .A2(new_n391), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1008), .B1(G107), .B2(new_n772), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n210), .B2(new_n758), .C1(new_n814), .C2(new_n768), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n321), .B1(new_n746), .B2(new_n748), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n755), .A2(new_n1021), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n765), .A2(new_n608), .B1(new_n257), .B2(new_n752), .ZN(new_n1197));
  NOR4_X1   g0997(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n746), .A2(new_n1078), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n756), .A2(new_n986), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(G50), .A2(new_n762), .B1(new_n764), .B2(new_n1071), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n767), .A2(G132), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1201), .A2(new_n1144), .A3(new_n292), .A4(new_n1202), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n771), .A2(new_n524), .B1(new_n752), .B2(new_n427), .ZN(new_n1204));
  NOR4_X1   g1004(.A1(new_n1199), .A2(new_n1200), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n740), .B1(new_n1198), .B2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1191), .A2(new_n1192), .A3(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n1111), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1209), .A2(new_n1116), .A3(new_n960), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1190), .A2(new_n1207), .A3(new_n1210), .ZN(G381));
  NAND2_X1  g1011(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1112), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT57), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n692), .B(new_n1177), .C1(new_n1214), .C2(new_n1183), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1215), .A2(new_n1122), .A3(new_n1173), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1216), .A2(G381), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT122), .Z(new_n1219));
  INV_X1    g1019(.A(G390), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1220), .A2(new_n965), .A3(new_n994), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1217), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT123), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1217), .A2(new_n1222), .A3(KEYINPUT123), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1225), .A2(new_n1226), .ZN(G407));
  INV_X1    g1027(.A(G213), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1228), .A2(G343), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1216), .A2(new_n1230), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1231), .A2(KEYINPUT124), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1228), .B1(new_n1231), .B2(KEYINPUT124), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(new_n1225), .C2(new_n1226), .ZN(G409));
  NAND2_X1  g1034(.A1(G375), .A2(G378), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1213), .A2(new_n960), .A3(new_n1172), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1179), .A2(new_n996), .A3(new_n1182), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1236), .A2(new_n1122), .A3(new_n1163), .A4(new_n1237), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1238), .A2(new_n1230), .ZN(new_n1239));
  INV_X1    g1039(.A(G384), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1111), .A2(new_n1105), .A3(KEYINPUT60), .A4(new_n1109), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1116), .A2(new_n1241), .A3(new_n692), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT60), .B1(new_n1208), .B2(new_n1111), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1187), .A2(new_n1189), .A3(new_n1207), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1240), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT60), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1248), .A2(new_n692), .A3(new_n1116), .A4(new_n1241), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1249), .A2(new_n1190), .A3(G384), .A4(new_n1207), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1246), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1235), .A2(new_n1239), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(KEYINPUT62), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1229), .A2(G2897), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1229), .A2(KEYINPUT125), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1246), .A2(new_n1250), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(KEYINPUT126), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT126), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1246), .A2(new_n1250), .A3(new_n1259), .A4(new_n1256), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1255), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1258), .A2(new_n1255), .A3(new_n1260), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1122), .B1(new_n1215), .B2(new_n1173), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1238), .A2(new_n1230), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1262), .B(new_n1263), .C1(new_n1264), .C2(new_n1265), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT62), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1235), .A2(new_n1239), .A3(new_n1268), .A4(new_n1252), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1254), .A2(new_n1266), .A3(new_n1267), .A4(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G387), .A2(G390), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1221), .ZN(new_n1272));
  XOR2_X1   g1072(.A(G393), .B(G396), .Z(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1273), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1271), .A2(new_n1221), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1270), .A2(new_n1277), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1264), .A2(new_n1265), .A3(new_n1251), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1277), .B1(new_n1279), .B2(KEYINPUT63), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT61), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT63), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1263), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1283), .A2(new_n1261), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1235), .A2(new_n1239), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1282), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1280), .B(new_n1281), .C1(new_n1286), .C2(new_n1279), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1278), .A2(new_n1287), .ZN(G405));
  NAND2_X1  g1088(.A1(new_n1235), .A2(new_n1216), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1252), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1235), .A2(new_n1216), .A3(new_n1251), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1277), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1292), .B(new_n1293), .ZN(G402));
endmodule


