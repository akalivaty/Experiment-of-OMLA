//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G228gat), .ZN(new_n206));
  INV_X1    g005(.A(G233gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G197gat), .B(G204gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT22), .ZN(new_n210));
  INV_X1    g009(.A(G211gat), .ZN(new_n211));
  INV_X1    g010(.A(G218gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G211gat), .B(G218gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT73), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n215), .A2(new_n209), .A3(new_n213), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n214), .A2(KEYINPUT73), .A3(new_n216), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT76), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(G155gat), .B2(G162gat), .ZN(new_n224));
  OR2_X1    g023(.A1(G141gat), .A2(G148gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(G141gat), .A2(G148gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n228), .B1(G155gat), .B2(G162gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n224), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G155gat), .B(G162gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G155gat), .ZN(new_n234));
  INV_X1    g033(.A(G162gat), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT2), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(new_n225), .A3(new_n226), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(new_n231), .A3(new_n224), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT3), .B1(new_n233), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n222), .B1(new_n239), .B2(KEYINPUT29), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT29), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n220), .A2(new_n241), .A3(new_n221), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n233), .A2(new_n238), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n208), .B(new_n240), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT79), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n230), .A2(new_n232), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n231), .B1(new_n237), .B2(new_n224), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT29), .B1(new_n217), .B2(new_n219), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n250), .B1(KEYINPUT3), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n240), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n208), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n247), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AOI211_X1 g054(.A(KEYINPUT79), .B(new_n208), .C1(new_n240), .C2(new_n252), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n246), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G22gat), .ZN(new_n258));
  INV_X1    g057(.A(G78gat), .ZN(new_n259));
  INV_X1    g058(.A(G22gat), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n246), .B(new_n260), .C1(new_n255), .C2(new_n256), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n258), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n259), .B1(new_n258), .B2(new_n261), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n205), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n258), .A2(new_n261), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G78gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n258), .A2(new_n259), .A3(new_n261), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(new_n267), .A3(new_n204), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(G15gat), .B(G43gat), .Z(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT70), .ZN(new_n272));
  XNOR2_X1  g071(.A(G71gat), .B(G99gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G227gat), .A2(G233gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT23), .ZN(new_n277));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT23), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(G169gat), .B2(G176gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  AND2_X1   g081(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT64), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n284), .A3(G190gat), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT64), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n285), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n282), .A2(new_n291), .A3(KEYINPUT25), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT25), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n287), .A2(new_n286), .B1(new_n283), .B2(G190gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n293), .B1(new_n281), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G183gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT27), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT27), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(G190gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n298), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT65), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT66), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n299), .A2(G183gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n297), .A2(KEYINPUT27), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n298), .A2(new_n300), .A3(KEYINPUT66), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n303), .A2(G190gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n302), .A2(KEYINPUT65), .A3(new_n303), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n306), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n276), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT26), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n287), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n318), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n315), .A2(KEYINPUT67), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT67), .B1(new_n315), .B2(new_n320), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n296), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G113gat), .B(G120gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(KEYINPUT1), .ZN(new_n325));
  XNOR2_X1  g124(.A(G127gat), .B(G134gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n326), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n328), .B1(KEYINPUT1), .B2(new_n324), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n323), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n330), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n332), .B(new_n296), .C1(new_n321), .C2(new_n322), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n275), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT68), .B(KEYINPUT33), .ZN(new_n335));
  OAI211_X1 g134(.A(KEYINPUT69), .B(new_n274), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT32), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n274), .A2(new_n335), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n334), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT69), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n341), .B(new_n274), .C1(new_n334), .C2(new_n335), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n331), .A2(new_n333), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT32), .B1(new_n343), .B2(new_n275), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n275), .A3(new_n333), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT71), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT34), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT34), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n346), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT72), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT34), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT34), .B1(new_n347), .B2(new_n348), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n351), .A2(KEYINPUT72), .A3(new_n352), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n359), .A2(new_n360), .A3(new_n345), .A4(new_n340), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT30), .ZN(new_n364));
  XNOR2_X1  g163(.A(G8gat), .B(G36gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n365), .B(new_n366), .Z(new_n367));
  XOR2_X1   g166(.A(new_n367), .B(KEYINPUT75), .Z(new_n368));
  AND2_X1   g167(.A1(G226gat), .A2(G233gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n369), .A2(KEYINPUT29), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n323), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT74), .ZN(new_n372));
  AOI221_X4 g171(.A(new_n372), .B1(new_n292), .B2(new_n295), .C1(new_n315), .C2(new_n320), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n315), .A2(new_n320), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT74), .B1(new_n374), .B2(new_n296), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n369), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n371), .A2(new_n376), .A3(new_n222), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n374), .A2(new_n296), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n372), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n374), .A2(KEYINPUT74), .A3(new_n296), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(new_n380), .A3(new_n370), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n296), .B(new_n369), .C1(new_n321), .C2(new_n322), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n222), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n368), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n222), .ZN(new_n385));
  INV_X1    g184(.A(new_n370), .ZN(new_n386));
  NOR3_X1   g185(.A1(new_n373), .A2(new_n375), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n382), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n371), .A2(new_n376), .A3(new_n222), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n367), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n364), .B1(new_n384), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n377), .A2(new_n383), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT30), .B1(new_n393), .B2(new_n367), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n332), .A2(new_n245), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n243), .B1(new_n248), .B2(new_n249), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n233), .A2(KEYINPUT3), .A3(new_n238), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n330), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(G225gat), .A2(G233gat), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n332), .A2(KEYINPUT4), .A3(new_n245), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n398), .A2(new_n401), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT5), .ZN(new_n405));
  OR2_X1    g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G1gat), .B(G29gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n407), .B(KEYINPUT0), .ZN(new_n408));
  XNOR2_X1  g207(.A(G57gat), .B(G85gat), .ZN(new_n409));
  XOR2_X1   g208(.A(new_n408), .B(new_n409), .Z(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n250), .A2(new_n330), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n402), .B1(new_n412), .B2(new_n396), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n404), .B1(new_n405), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT77), .B(KEYINPUT6), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n406), .A2(new_n411), .A3(new_n414), .A4(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n406), .A2(new_n411), .A3(new_n414), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n415), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n411), .B1(new_n406), .B2(new_n414), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n363), .B1(new_n395), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n367), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n377), .A2(new_n383), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n368), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n389), .B2(new_n390), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT30), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n391), .A2(new_n364), .ZN(new_n428));
  AND4_X1   g227(.A1(new_n363), .A2(new_n421), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n270), .B(new_n362), .C1(new_n422), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT35), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n353), .A2(new_n340), .A3(new_n345), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n353), .B1(new_n345), .B2(new_n340), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n432), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n355), .A2(KEYINPUT82), .A3(new_n433), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n269), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n395), .A2(new_n421), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n439), .A2(KEYINPUT35), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n431), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(KEYINPUT78), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n395), .A2(new_n363), .A3(new_n421), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n444), .A3(new_n269), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT40), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n398), .A2(new_n401), .A3(new_n403), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT39), .ZN(new_n448));
  INV_X1    g247(.A(new_n402), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n410), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n412), .A2(new_n396), .A3(new_n402), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT39), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n453), .B1(new_n449), .B2(new_n447), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n446), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n447), .A2(new_n449), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n456), .A2(KEYINPUT39), .A3(new_n452), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n457), .A2(KEYINPUT40), .A3(new_n410), .A4(new_n450), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n455), .A2(new_n458), .A3(new_n418), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(new_n392), .B2(new_n394), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n460), .A2(new_n268), .A3(new_n264), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT81), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT37), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n393), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n389), .A2(new_n463), .A3(new_n390), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT81), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(KEYINPUT80), .B(KEYINPUT38), .Z(new_n468));
  NAND2_X1  g267(.A1(new_n368), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n371), .A2(new_n376), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n463), .B1(new_n470), .B2(new_n385), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n222), .B1(new_n387), .B2(new_n388), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n421), .A2(new_n424), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n423), .B1(new_n393), .B2(new_n463), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n476), .B1(new_n466), .B2(new_n464), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n474), .B(new_n475), .C1(new_n477), .C2(new_n468), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT36), .B1(new_n355), .B2(new_n433), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n355), .A2(KEYINPUT36), .A3(new_n361), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n445), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n442), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(G15gat), .B(G22gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT87), .ZN(new_n485));
  INV_X1    g284(.A(G1gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(KEYINPUT87), .A3(G1gat), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT16), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  XOR2_X1   g290(.A(new_n491), .B(G8gat), .Z(new_n492));
  XOR2_X1   g291(.A(KEYINPUT84), .B(G29gat), .Z(new_n493));
  INV_X1    g292(.A(G36gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(G29gat), .A2(G36gat), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n496), .A2(KEYINPUT14), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(KEYINPUT14), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G43gat), .B(G50gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT83), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OR2_X1    g302(.A1(G43gat), .A2(G50gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(G43gat), .A2(G50gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(KEYINPUT83), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(KEYINPUT15), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n501), .A2(KEYINPUT15), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n500), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n503), .A2(KEYINPUT15), .A3(new_n506), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n497), .B(new_n498), .C1(new_n493), .C2(new_n494), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n510), .A2(KEYINPUT17), .A3(new_n513), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n492), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT86), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n511), .A2(new_n508), .A3(new_n512), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n500), .A2(new_n507), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT85), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT85), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n510), .A2(new_n520), .A3(new_n513), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT17), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n516), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI211_X1 g323(.A(KEYINPUT86), .B(KEYINPUT17), .C1(new_n519), .C2(new_n521), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n515), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n492), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n522), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT18), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(G229gat), .B2(G233gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n526), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT88), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT88), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n526), .A2(new_n533), .A3(new_n528), .A4(new_n530), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G113gat), .B(G141gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(G197gat), .ZN(new_n537));
  XOR2_X1   g336(.A(KEYINPUT11), .B(G169gat), .Z(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n539), .B(KEYINPUT12), .Z(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT13), .ZN(new_n543));
  INV_X1    g342(.A(new_n522), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n492), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n543), .B1(new_n545), .B2(new_n528), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n526), .A2(new_n528), .A3(new_n542), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(new_n529), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n535), .A2(new_n541), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n541), .B1(new_n535), .B2(new_n548), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n483), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT89), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT90), .B(G57gat), .ZN(new_n555));
  MUX2_X1   g354(.A(G57gat), .B(new_n555), .S(G64gat), .Z(new_n556));
  AOI21_X1  g355(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(G71gat), .B(G78gat), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n558), .B2(KEYINPUT91), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n556), .B(new_n559), .C1(KEYINPUT91), .C2(new_n558), .ZN(new_n560));
  XOR2_X1   g359(.A(G57gat), .B(G64gat), .Z(new_n561));
  AND2_X1   g360(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n560), .B1(new_n558), .B2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(KEYINPUT92), .B(KEYINPUT21), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G127gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT21), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n492), .B1(new_n569), .B2(new_n563), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n568), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G183gat), .B(G211gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT93), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(new_n234), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n571), .A2(new_n577), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT95), .B(KEYINPUT7), .ZN(new_n581));
  NAND2_X1  g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n582), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  INV_X1    g384(.A(G85gat), .ZN(new_n586));
  INV_X1    g385(.A(G92gat), .ZN(new_n587));
  AOI22_X1  g386(.A1(KEYINPUT8), .A2(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n583), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G99gat), .B(G106gat), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n514), .ZN(new_n592));
  INV_X1    g391(.A(new_n521), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n520), .B1(new_n510), .B2(new_n513), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n523), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT86), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n522), .A2(new_n516), .A3(new_n523), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n592), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n599), .B1(new_n544), .B2(new_n591), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G190gat), .B(G218gat), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT94), .ZN(new_n607));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n601), .A2(new_n603), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n605), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n609), .B1(new_n605), .B2(new_n610), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n580), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n591), .A2(new_n563), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT10), .B1(new_n619), .B2(KEYINPUT96), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n591), .A2(new_n563), .ZN(new_n622));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT97), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n619), .A2(KEYINPUT96), .A3(KEYINPUT10), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n621), .A2(new_n622), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n623), .B1(new_n619), .B2(new_n622), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n618), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n621), .A2(new_n622), .A3(new_n623), .A4(new_n626), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n629), .A2(new_n618), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n615), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n554), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n421), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(KEYINPUT98), .B(G1gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(G1324gat));
  INV_X1    g441(.A(new_n395), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(G8gat), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT42), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT16), .B(G8gat), .Z(new_n647));
  NAND3_X1  g446(.A1(new_n638), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(new_n649), .A3(new_n646), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n649), .B1(new_n648), .B2(new_n646), .ZN(new_n652));
  OAI221_X1 g451(.A(new_n645), .B1(new_n646), .B2(new_n648), .C1(new_n651), .C2(new_n652), .ZN(G1325gat));
  INV_X1    g452(.A(G15gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n436), .A2(new_n437), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n638), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(KEYINPUT100), .B1(new_n481), .B2(new_n480), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT36), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(new_n434), .B2(new_n435), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n355), .A2(new_n361), .A3(KEYINPUT36), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT100), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n638), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n656), .B1(new_n666), .B2(new_n654), .ZN(G1326gat));
  NAND2_X1  g466(.A1(new_n638), .A2(new_n269), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT101), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT43), .B(G22gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  INV_X1    g470(.A(new_n580), .ZN(new_n672));
  INV_X1    g471(.A(new_n614), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n672), .A2(new_n673), .A3(new_n634), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n554), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(new_n639), .A3(new_n493), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT45), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n678), .B1(new_n483), .B2(new_n614), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n657), .A2(new_n445), .A3(new_n479), .A4(new_n662), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n422), .A2(new_n429), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n683), .A2(new_n269), .B1(new_n478), .B2(new_n461), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n684), .A2(KEYINPUT103), .A3(new_n657), .A4(new_n662), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT104), .B1(new_n686), .B2(new_n442), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n688));
  AOI22_X1  g487(.A1(new_n430), .A2(KEYINPUT35), .B1(new_n438), .B2(new_n440), .ZN(new_n689));
  AOI211_X1 g488(.A(new_n688), .B(new_n689), .C1(new_n682), .C2(new_n685), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n612), .B2(new_n613), .ZN(new_n693));
  INV_X1    g492(.A(new_n609), .ZN(new_n694));
  INV_X1    g493(.A(new_n610), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(new_n604), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n696), .A2(KEYINPUT105), .A3(new_n611), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n698), .A2(KEYINPUT44), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n679), .B1(new_n691), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n549), .B2(new_n550), .ZN(new_n702));
  INV_X1    g501(.A(new_n528), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n596), .A2(new_n597), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n703), .B1(new_n704), .B2(new_n515), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n533), .B1(new_n705), .B2(new_n530), .ZN(new_n706));
  INV_X1    g505(.A(new_n534), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n548), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n540), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n535), .A2(new_n541), .A3(new_n548), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n709), .A2(KEYINPUT102), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n702), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n713), .A2(new_n580), .A3(new_n635), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n700), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n421), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n677), .B1(new_n493), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT106), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n677), .B(new_n720), .C1(new_n493), .C2(new_n717), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(G1328gat));
  NAND3_X1  g521(.A1(new_n675), .A2(new_n494), .A3(new_n643), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT46), .Z(new_n724));
  OAI21_X1  g523(.A(G36gat), .B1(new_n716), .B2(new_n395), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(G1329gat));
  OAI21_X1  g525(.A(G43gat), .B1(new_n716), .B2(new_n663), .ZN(new_n727));
  AOI21_X1  g526(.A(G43gat), .B1(new_n436), .B2(new_n437), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n675), .A2(new_n728), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n727), .B(new_n729), .C1(KEYINPUT107), .C2(KEYINPUT47), .ZN(new_n730));
  NAND2_X1  g529(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1330gat));
  INV_X1    g531(.A(G50gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n715), .A2(new_n269), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n733), .B1(new_n734), .B2(KEYINPUT108), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(KEYINPUT108), .B2(new_n734), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n675), .A2(new_n733), .A3(new_n269), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n736), .A2(KEYINPUT48), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n737), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(G50gat), .B2(new_n734), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(KEYINPUT48), .B2(new_n740), .ZN(G1331gat));
  NAND3_X1  g540(.A1(new_n615), .A2(new_n634), .A3(new_n712), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT109), .Z(new_n743));
  NOR3_X1   g542(.A1(new_n743), .A2(new_n687), .A3(new_n690), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n639), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT110), .Z(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(new_n555), .ZN(G1332gat));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n643), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT49), .B(G64gat), .Z(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n748), .B2(new_n750), .ZN(G1333gat));
  INV_X1    g550(.A(G71gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n744), .A2(new_n752), .A3(new_n655), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n744), .A2(new_n664), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n754), .B2(new_n752), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g555(.A1(new_n744), .A2(new_n269), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g557(.A1(new_n686), .A2(new_n442), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n759), .A2(KEYINPUT112), .A3(new_n614), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n713), .A2(new_n672), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n689), .B1(new_n682), .B2(new_n685), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n763), .B2(new_n673), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n760), .A2(new_n761), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n760), .A2(new_n764), .A3(KEYINPUT51), .A4(new_n761), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n634), .A2(new_n586), .A3(new_n639), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(KEYINPUT113), .Z(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n761), .A2(new_n634), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n700), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n774), .ZN(new_n777));
  INV_X1    g576(.A(new_n699), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n687), .A2(new_n690), .A3(new_n778), .ZN(new_n779));
  OAI211_X1 g578(.A(KEYINPUT111), .B(new_n777), .C1(new_n779), .C2(new_n679), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n776), .A2(new_n781), .A3(new_n421), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n772), .B1(new_n782), .B2(new_n586), .ZN(G1336gat));
  NAND3_X1  g582(.A1(new_n775), .A2(new_n643), .A3(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G92gat), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n769), .A2(new_n587), .A3(new_n643), .A4(new_n634), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n700), .A2(new_n774), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n587), .B1(new_n789), .B2(new_n643), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n786), .A2(new_n788), .ZN(new_n791));
  OAI22_X1  g590(.A1(new_n787), .A2(new_n788), .B1(new_n790), .B2(new_n791), .ZN(G1337gat));
  INV_X1    g591(.A(G99gat), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n769), .A2(new_n793), .A3(new_n655), .A4(new_n634), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n776), .A2(new_n781), .A3(new_n663), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(new_n793), .ZN(G1338gat));
  NOR3_X1   g595(.A1(new_n270), .A2(G106gat), .A3(new_n635), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n798), .B1(new_n767), .B2(new_n768), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(KEYINPUT53), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n700), .A2(new_n270), .A3(new_n774), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n203), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n775), .A2(new_n269), .A3(new_n780), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n799), .B1(new_n803), .B2(G106gat), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT114), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n802), .B(new_n808), .C1(new_n804), .C2(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(G1339gat));
  NOR2_X1   g609(.A1(new_n636), .A2(new_n713), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n705), .A2(new_n542), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n545), .A2(new_n528), .A3(new_n543), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n539), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n710), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n813), .B1(new_n710), .B2(new_n816), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n626), .A2(new_n622), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n624), .B1(new_n820), .B2(new_n620), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n821), .A2(new_n631), .A3(KEYINPUT54), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n618), .B1(new_n627), .B2(KEYINPUT54), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n819), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n627), .A2(KEYINPUT54), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n821), .A2(new_n631), .A3(KEYINPUT54), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n825), .A2(new_n826), .A3(KEYINPUT55), .A4(new_n618), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n824), .A2(new_n827), .A3(new_n633), .ZN(new_n828));
  NOR4_X1   g627(.A1(new_n698), .A2(new_n817), .A3(new_n818), .A4(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n693), .A2(new_n697), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n824), .A2(new_n633), .A3(new_n827), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n702), .A2(new_n711), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n710), .A2(new_n634), .A3(new_n816), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n830), .B1(new_n834), .B2(KEYINPUT116), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n832), .A2(new_n836), .A3(new_n833), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n829), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n812), .B1(new_n838), .B2(new_n672), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n421), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n270), .A2(new_n362), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(new_n643), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g643(.A(new_n844), .B(KEYINPUT117), .Z(new_n845));
  INV_X1    g644(.A(G113gat), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n846), .A3(new_n713), .ZN(new_n847));
  INV_X1    g646(.A(new_n438), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n395), .A2(new_n639), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n840), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n552), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n847), .B1(new_n846), .B2(new_n852), .ZN(G1340gat));
  INV_X1    g652(.A(G120gat), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n845), .A2(new_n854), .A3(new_n634), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n850), .A2(new_n634), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n855), .B1(new_n854), .B2(new_n857), .ZN(G1341gat));
  INV_X1    g657(.A(new_n844), .ZN(new_n859));
  INV_X1    g658(.A(G127gat), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n860), .A3(new_n672), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n850), .A2(new_n672), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n860), .B2(new_n863), .ZN(G1342gat));
  OR3_X1    g663(.A1(new_n844), .A2(G134gat), .A3(new_n673), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n614), .ZN(new_n866));
  AOI22_X1  g665(.A1(new_n865), .A2(KEYINPUT56), .B1(G134gat), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n867), .B1(KEYINPUT56), .B2(new_n865), .ZN(G1343gat));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n664), .A2(new_n849), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n270), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n829), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n833), .B1(new_n551), .B2(new_n828), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n673), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n672), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n873), .B1(new_n877), .B2(new_n811), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n839), .B2(new_n269), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI211_X1 g680(.A(KEYINPUT118), .B(KEYINPUT57), .C1(new_n839), .C2(new_n269), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n713), .B(new_n871), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(G141gat), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n663), .A2(new_n269), .ZN(new_n885));
  XOR2_X1   g684(.A(new_n885), .B(KEYINPUT119), .Z(new_n886));
  NAND3_X1  g685(.A1(new_n839), .A2(new_n886), .A3(new_n639), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n551), .A2(G141gat), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n395), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n870), .B1(new_n884), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n887), .A2(KEYINPUT120), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n839), .A2(new_n886), .A3(new_n895), .A4(new_n639), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n395), .A3(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n889), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n870), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n552), .B(new_n871), .C1(new_n881), .C2(new_n882), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(G141gat), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n869), .B1(new_n893), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(G141gat), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n894), .A2(new_n395), .A3(new_n896), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT58), .B1(new_n904), .B2(new_n889), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  AOI22_X1  g705(.A1(new_n883), .A2(G141gat), .B1(new_n888), .B2(new_n891), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n906), .B(KEYINPUT121), .C1(new_n870), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n902), .A2(new_n908), .ZN(G1344gat));
  NOR2_X1   g708(.A1(new_n817), .A2(new_n818), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n614), .A3(new_n831), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n672), .B1(new_n911), .B2(new_n876), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n636), .A2(new_n552), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n269), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n872), .ZN(new_n915));
  XOR2_X1   g714(.A(new_n915), .B(KEYINPUT122), .Z(new_n916));
  AND2_X1   g715(.A1(new_n839), .A2(new_n873), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n871), .A2(new_n634), .ZN(new_n919));
  OAI21_X1  g718(.A(G148gat), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT59), .ZN(new_n921));
  INV_X1    g720(.A(G148gat), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(KEYINPUT59), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n871), .B1(new_n881), .B2(new_n882), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n924), .B2(new_n635), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n904), .A2(new_n922), .A3(new_n634), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1345gat));
  OAI21_X1  g727(.A(G155gat), .B1(new_n924), .B2(new_n580), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n904), .A2(new_n234), .A3(new_n672), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1346gat));
  OAI21_X1  g730(.A(G162gat), .B1(new_n924), .B2(new_n698), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n904), .A2(new_n235), .A3(new_n614), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1347gat));
  NAND2_X1  g733(.A1(new_n643), .A2(new_n421), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n840), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n438), .ZN(new_n937));
  INV_X1    g736(.A(G169gat), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n937), .A2(new_n938), .A3(new_n551), .ZN(new_n939));
  INV_X1    g738(.A(new_n842), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n713), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n939), .B1(new_n938), .B2(new_n943), .ZN(G1348gat));
  AOI21_X1  g743(.A(G176gat), .B1(new_n942), .B2(new_n634), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n936), .A2(G176gat), .A3(new_n438), .A4(new_n634), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n945), .A2(new_n948), .A3(new_n949), .ZN(G1349gat));
  NAND3_X1  g749(.A1(new_n936), .A2(new_n438), .A3(new_n672), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n297), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n953), .B1(new_n952), .B2(new_n951), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n672), .A2(new_n310), .A3(new_n311), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT125), .B1(new_n942), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT60), .ZN(G1350gat));
  NOR3_X1   g757(.A1(new_n941), .A2(G190gat), .A3(new_n698), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n936), .A2(new_n438), .A3(new_n614), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n960), .A2(G190gat), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n961), .A2(KEYINPUT126), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n961), .A2(KEYINPUT126), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT61), .B1(new_n961), .B2(KEYINPUT126), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(G1351gat));
  INV_X1    g766(.A(new_n918), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n664), .A2(new_n935), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(G197gat), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n970), .A2(new_n971), .A3(new_n551), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n840), .A2(new_n270), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(new_n969), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(G197gat), .B1(new_n975), .B2(new_n713), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n972), .A2(new_n976), .ZN(G1352gat));
  OR3_X1    g776(.A1(new_n974), .A2(G204gat), .A3(new_n635), .ZN(new_n978));
  OR2_X1    g777(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n979));
  OAI21_X1  g778(.A(G204gat), .B1(new_n970), .B2(new_n635), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n981), .A2(KEYINPUT127), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n981), .A2(KEYINPUT127), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n979), .B(new_n980), .C1(new_n982), .C2(new_n983), .ZN(G1353gat));
  NAND3_X1  g783(.A1(new_n975), .A2(new_n211), .A3(new_n672), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n968), .A2(new_n672), .A3(new_n969), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n986), .B2(G211gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(G1354gat));
  OAI21_X1  g788(.A(G218gat), .B1(new_n970), .B2(new_n673), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n975), .A2(new_n212), .A3(new_n830), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1355gat));
endmodule


