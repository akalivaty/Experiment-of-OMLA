//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1229, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n209), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n222), .A2(new_n223), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n211), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n214), .B(new_n219), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  OAI21_X1  g0046(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT65), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n249));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n247), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G226), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(G223), .ZN(new_n258));
  INV_X1    g0058(.A(G77), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n257), .A2(new_n258), .B1(new_n259), .B2(new_n256), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G1698), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n260), .B1(G222), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n249), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n252), .B(new_n255), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G190), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n271), .B1(G200), .B2(new_n269), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n273), .A2(new_n217), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n276));
  INV_X1    g0076(.A(G150), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n209), .A2(G33), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n275), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  XOR2_X1   g0084(.A(new_n284), .B(KEYINPUT66), .Z(new_n285));
  NAND3_X1  g0085(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n286));
  INV_X1    g0086(.A(G50), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n275), .B1(new_n208), .B2(G20), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n288), .B1(new_n289), .B2(new_n287), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT67), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(KEYINPUT9), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT9), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(new_n285), .B2(new_n291), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n272), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n269), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n300), .A2(KEYINPUT68), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(KEYINPUT68), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n292), .B(new_n299), .C1(new_n304), .C2(new_n269), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT12), .B1(new_n286), .B2(G68), .ZN(new_n307));
  OR3_X1    g0107(.A1(new_n286), .A2(KEYINPUT12), .A3(G68), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n289), .A2(G68), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n279), .A2(new_n287), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n282), .A2(new_n259), .B1(new_n209), .B2(G68), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n275), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT11), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n313), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n309), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT73), .ZN(new_n317));
  INV_X1    g0117(.A(G1698), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n256), .A2(G226), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n256), .A2(G232), .A3(G1698), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G33), .A2(G97), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT72), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT72), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n319), .A2(new_n320), .A3(new_n324), .A4(new_n321), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n249), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT13), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n248), .A2(new_n251), .B1(new_n254), .B2(G238), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n327), .B1(new_n326), .B2(new_n328), .ZN(new_n330));
  OAI21_X1  g0130(.A(G169), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n329), .A2(new_n330), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n331), .A2(KEYINPUT14), .B1(new_n332), .B2(G179), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT14), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n334), .B(G169), .C1(new_n329), .C2(new_n330), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT74), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n331), .A2(KEYINPUT14), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n332), .A2(G179), .ZN(new_n338));
  AND4_X1   g0138(.A1(KEYINPUT74), .A2(new_n337), .A3(new_n335), .A4(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n317), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n317), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n332), .A2(G190), .ZN(new_n342));
  OAI21_X1  g0142(.A(G200), .B1(new_n329), .B2(new_n330), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  XOR2_X1   g0145(.A(KEYINPUT8), .B(G58), .Z(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT69), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT69), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n281), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n279), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT15), .B(G87), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n351), .A2(new_n282), .B1(new_n209), .B2(new_n259), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n275), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT70), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g0155(.A(KEYINPUT70), .B(new_n275), .C1(new_n350), .C2(new_n352), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT71), .B1(new_n286), .B2(G77), .ZN(new_n358));
  OR3_X1    g0158(.A1(new_n286), .A2(KEYINPUT71), .A3(G77), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n289), .A2(G77), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n254), .A2(G244), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n252), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n256), .A2(G232), .A3(new_n318), .ZN(new_n364));
  INV_X1    g0164(.A(G238), .ZN(new_n365));
  OAI221_X1 g0165(.A(new_n364), .B1(new_n205), .B2(new_n256), .C1(new_n257), .C2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n363), .B1(new_n249), .B2(new_n366), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n367), .A2(G169), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n303), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n361), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n366), .A2(new_n249), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n371), .A2(G190), .A3(new_n252), .A4(new_n362), .ZN(new_n372));
  INV_X1    g0172(.A(G200), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n372), .B1(new_n367), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n370), .B1(new_n361), .B2(new_n374), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n306), .A2(new_n345), .A3(new_n375), .ZN(new_n376));
  XOR2_X1   g0176(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n377));
  INV_X1    g0177(.A(G58), .ZN(new_n378));
  INV_X1    g0178(.A(G68), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n380), .A2(new_n201), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(G20), .B1(G159), .B2(new_n278), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT76), .ZN(new_n383));
  OR3_X1    g0183(.A1(new_n263), .A2(KEYINPUT76), .A3(KEYINPUT3), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT7), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n385), .A2(G20), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n383), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n385), .B1(new_n256), .B2(G20), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n379), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n382), .B1(new_n389), .B2(KEYINPUT77), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT77), .ZN(new_n391));
  AOI211_X1 g0191(.A(new_n391), .B(new_n379), .C1(new_n387), .C2(new_n388), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n377), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT78), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g0195(.A(KEYINPUT78), .B(new_n377), .C1(new_n390), .C2(new_n392), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n265), .A2(new_n386), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n388), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(G68), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n399), .A2(KEYINPUT16), .A3(new_n382), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n275), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n395), .A2(new_n396), .A3(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n262), .A2(new_n264), .A3(G223), .A4(new_n318), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT79), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT79), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n256), .A2(new_n406), .A3(G223), .A4(new_n318), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G87), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n262), .A2(new_n264), .A3(G226), .A4(G1698), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n405), .A2(new_n407), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT80), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n409), .A2(new_n408), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT80), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n412), .A2(new_n413), .A3(new_n407), .A4(new_n405), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n411), .A2(new_n414), .A3(new_n249), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n254), .A2(G232), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n252), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n415), .A2(new_n270), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n268), .B1(new_n410), .B2(KEYINPUT80), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n417), .B1(new_n420), .B2(new_n414), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n419), .B(KEYINPUT81), .C1(G200), .C2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n286), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n346), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n289), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n424), .B1(new_n425), .B2(new_n346), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT81), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n421), .A2(new_n428), .A3(new_n270), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n403), .A2(new_n422), .A3(new_n427), .A4(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n401), .B1(new_n393), .B2(new_n394), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n426), .B1(new_n433), .B2(new_n396), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n434), .A2(KEYINPUT17), .A3(new_n422), .A4(new_n429), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT82), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n403), .A2(new_n427), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT18), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n415), .A2(new_n304), .A3(new_n418), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n298), .B2(new_n421), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n439), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n440), .B1(new_n439), .B2(new_n442), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n432), .A2(new_n435), .A3(KEYINPUT82), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n438), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n376), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n256), .A2(G264), .A3(G1698), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n265), .A2(G303), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n256), .A2(new_n318), .ZN(new_n453));
  INV_X1    g0253(.A(G257), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n451), .B(new_n452), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n249), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n208), .A2(G45), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  XNOR2_X1  g0258(.A(KEYINPUT5), .B(G41), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n249), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n459), .A2(new_n458), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n460), .A2(G270), .B1(new_n461), .B2(new_n251), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G116), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n423), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n208), .A2(G33), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n286), .A2(new_n466), .A3(new_n217), .A4(new_n273), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n273), .A2(new_n217), .B1(G20), .B2(new_n464), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G283), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n469), .B(new_n209), .C1(G33), .C2(new_n204), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n468), .A2(KEYINPUT20), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT20), .B1(new_n468), .B2(new_n470), .ZN(new_n472));
  OAI221_X1 g0272(.A(new_n465), .B1(new_n464), .B2(new_n467), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n463), .A2(new_n473), .A3(G169), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT21), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n463), .A2(new_n473), .A3(KEYINPUT21), .A4(G169), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n456), .A2(G179), .A3(new_n462), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n473), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n476), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n456), .A2(G190), .A3(new_n462), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n473), .B1(new_n463), .B2(G200), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n256), .A2(G238), .A3(new_n318), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n256), .A2(G244), .A3(G1698), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G116), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n249), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n457), .A2(G250), .ZN(new_n490));
  OAI22_X1  g0290(.A1(new_n249), .A2(new_n490), .B1(new_n250), .B2(new_n457), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G200), .ZN(new_n494));
  INV_X1    g0294(.A(new_n351), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n286), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n256), .A2(new_n209), .A3(G68), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT19), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n209), .B1(new_n321), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(G87), .B2(new_n206), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n498), .B1(new_n282), .B2(new_n204), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n497), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n496), .B1(new_n502), .B2(new_n275), .ZN(new_n503));
  INV_X1    g0303(.A(new_n467), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(KEYINPUT85), .A3(G87), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT85), .ZN(new_n506));
  INV_X1    g0306(.A(G87), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n506), .B1(new_n467), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n491), .B1(new_n488), .B2(new_n249), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G190), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n494), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n460), .A2(G257), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n461), .A2(new_n251), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT4), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT83), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n266), .A2(G244), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n256), .A2(G244), .A3(new_n318), .ZN(new_n520));
  INV_X1    g0320(.A(new_n518), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n256), .A2(G250), .A3(G1698), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n519), .A2(new_n469), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n516), .B1(new_n524), .B2(new_n249), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n303), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n523), .B(new_n469), .C1(new_n520), .C2(new_n521), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n518), .B1(new_n266), .B2(G244), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n249), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n514), .A2(new_n515), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n298), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT6), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n533), .A2(new_n204), .A3(G107), .ZN(new_n534));
  XNOR2_X1  g0334(.A(G97), .B(G107), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n534), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n536), .A2(new_n209), .B1(new_n259), .B2(new_n279), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n205), .B1(new_n387), .B2(new_n388), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n275), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n286), .A2(G97), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n504), .B2(G97), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n526), .A2(new_n532), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n531), .A2(G200), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n539), .A2(new_n541), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n529), .A2(new_n530), .A3(G190), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n489), .A2(new_n304), .A3(new_n492), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n298), .B2(new_n511), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n504), .A2(new_n495), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n503), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT84), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n503), .A2(KEYINPUT84), .A3(new_n550), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n549), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AND4_X1   g0355(.A1(new_n513), .A2(new_n543), .A3(new_n547), .A4(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n256), .A2(G250), .A3(new_n318), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n256), .A2(G257), .A3(G1698), .ZN(new_n558));
  XNOR2_X1  g0358(.A(KEYINPUT88), .B(G294), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n557), .B(new_n558), .C1(new_n263), .C2(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n560), .A2(new_n249), .B1(G264), .B2(new_n460), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(new_n300), .A3(new_n515), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n249), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n460), .A2(G264), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n515), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n298), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n262), .A2(new_n264), .A3(new_n209), .A4(G87), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT86), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT22), .ZN(new_n569));
  OR3_X1    g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n569), .ZN(new_n571));
  NAND2_X1  g0371(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n567), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(KEYINPUT23), .B1(new_n209), .B2(G107), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT87), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT87), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n576), .B(KEYINPUT23), .C1(new_n209), .C2(G107), .ZN(new_n577));
  OR3_X1    g0377(.A1(new_n209), .A2(KEYINPUT23), .A3(G107), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n209), .A2(G33), .A3(G116), .ZN(new_n579));
  AND4_X1   g0379(.A1(new_n575), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n570), .A2(new_n573), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT24), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n572), .B1(new_n567), .B2(new_n571), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n575), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT24), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n586), .A3(new_n573), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n274), .B1(new_n582), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT25), .B1(new_n423), .B2(new_n205), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n423), .A2(KEYINPUT25), .A3(new_n205), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n590), .A2(new_n591), .B1(new_n504), .B2(G107), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n562), .B(new_n566), .C1(new_n588), .C2(new_n593), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n585), .A2(new_n586), .A3(new_n573), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n586), .B1(new_n585), .B2(new_n573), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n275), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n561), .A2(G190), .A3(new_n515), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n565), .A2(G200), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n597), .A2(new_n592), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n484), .A2(new_n556), .A3(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n450), .A2(new_n602), .ZN(G372));
  AND3_X1   g0403(.A1(new_n432), .A2(KEYINPUT82), .A3(new_n435), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT82), .B1(new_n432), .B2(new_n435), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n344), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n340), .A2(new_n370), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n445), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n297), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n610), .A2(new_n305), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n373), .B1(new_n489), .B2(new_n492), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n503), .A2(new_n509), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n512), .A2(new_n614), .B1(new_n549), .B2(new_n551), .ZN(new_n615));
  AND4_X1   g0415(.A1(new_n600), .A2(new_n615), .A3(new_n543), .A4(new_n547), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n566), .A2(new_n562), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n597), .B2(new_n592), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT89), .B1(new_n618), .B2(new_n481), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT89), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n474), .A2(new_n475), .B1(new_n479), .B2(new_n473), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n594), .A2(new_n620), .A3(new_n621), .A4(new_n477), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n616), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT26), .ZN(new_n624));
  INV_X1    g0424(.A(new_n554), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT84), .B1(new_n503), .B2(new_n550), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n627), .A2(new_n549), .B1(new_n512), .B2(new_n614), .ZN(new_n628));
  INV_X1    g0428(.A(new_n543), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n624), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n511), .A2(new_n298), .ZN(new_n631));
  AOI211_X1 g0431(.A(new_n303), .B(new_n491), .C1(new_n488), .C2(new_n249), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n551), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n531), .A2(new_n298), .B1(new_n539), .B2(new_n541), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(new_n513), .A3(new_n633), .A4(new_n526), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n633), .B1(new_n635), .B2(KEYINPUT26), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n623), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n450), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n611), .A2(new_n639), .ZN(G369));
  INV_X1    g0440(.A(G330), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G213), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n473), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n484), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n481), .A2(new_n473), .A3(new_n647), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n641), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n618), .A2(new_n647), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT90), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n653), .B(new_n647), .C1(new_n588), .C2(new_n593), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n594), .A2(new_n654), .A3(new_n600), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n597), .A2(new_n592), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n653), .B1(new_n656), .B2(new_n647), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n652), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n594), .A2(new_n647), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n655), .A2(new_n657), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n647), .B1(new_n621), .B2(new_n477), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n659), .A2(new_n663), .ZN(G399));
  INV_X1    g0464(.A(new_n212), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G41), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G1), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n215), .B2(new_n667), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT28), .ZN(new_n671));
  INV_X1    g0471(.A(new_n647), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n484), .A2(new_n556), .A3(new_n601), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n561), .A2(new_n511), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n478), .ZN(new_n675));
  AOI21_X1  g0475(.A(KEYINPUT30), .B1(new_n675), .B2(new_n525), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n304), .B1(new_n456), .B2(new_n462), .ZN(new_n677));
  AND4_X1   g0477(.A1(new_n565), .A2(new_n531), .A3(new_n677), .A4(new_n493), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n561), .A2(new_n511), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n680), .A2(new_n479), .A3(KEYINPUT30), .A4(new_n525), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OAI211_X1 g0482(.A(KEYINPUT31), .B(new_n647), .C1(new_n679), .C2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n673), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT91), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n678), .B1(new_n676), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n681), .A2(new_n685), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n680), .A2(new_n479), .A3(new_n525), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT30), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n672), .B1(new_n686), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(KEYINPUT31), .ZN(new_n693));
  OAI21_X1  g0493(.A(G330), .B1(new_n684), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n633), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n635), .A2(new_n624), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT92), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n555), .A2(new_n513), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n624), .B1(new_n699), .B2(new_n543), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n629), .A2(new_n615), .A3(KEYINPUT26), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n701), .A3(KEYINPUT92), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n594), .A2(new_n477), .A3(new_n621), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n543), .A2(new_n547), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n703), .A2(new_n704), .A3(new_n600), .A4(new_n615), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n698), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n706), .A2(KEYINPUT29), .A3(new_n672), .ZN(new_n707));
  AOI21_X1  g0507(.A(KEYINPUT29), .B1(new_n638), .B2(new_n672), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n694), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n671), .B1(new_n710), .B2(G1), .ZN(G364));
  NAND2_X1  g0511(.A1(new_n649), .A2(new_n650), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n713), .A2(KEYINPUT93), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(G330), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n209), .A2(G13), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT94), .ZN(new_n717));
  INV_X1    g0517(.A(G45), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(KEYINPUT95), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n208), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n719), .A2(KEYINPUT95), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n666), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n713), .A2(KEYINPUT93), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n714), .A2(new_n715), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n212), .A2(new_n256), .ZN(new_n728));
  INV_X1    g0528(.A(G355), .ZN(new_n729));
  OAI22_X1  g0529(.A1(new_n728), .A2(new_n729), .B1(G116), .B2(new_n212), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n665), .A2(new_n256), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n718), .B2(new_n216), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n242), .A2(new_n718), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n730), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G13), .A2(G33), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n217), .B1(G20), .B2(new_n298), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n724), .B1(new_n735), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n209), .A2(new_n270), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n373), .A2(G179), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G303), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n265), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n743), .A2(new_n373), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n303), .A2(new_n748), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n749), .A2(G322), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n270), .A2(G20), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n303), .A2(new_n373), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g0552(.A(KEYINPUT33), .B(G317), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n747), .B(new_n750), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G179), .A2(G200), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT97), .ZN(new_n756));
  OAI21_X1  g0556(.A(G20), .B1(new_n756), .B2(new_n270), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n751), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n304), .A2(new_n373), .A3(new_n759), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n760), .A2(KEYINPUT96), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(KEYINPUT96), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G311), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n754), .B1(new_n559), .B2(new_n758), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n756), .A2(new_n751), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n759), .A2(new_n744), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n766), .A2(G329), .B1(G283), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT99), .ZN(new_n770));
  INV_X1    g0570(.A(G326), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n304), .A2(G200), .A3(new_n743), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT98), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n770), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n766), .A2(G159), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT32), .Z(new_n776));
  NAND2_X1  g0576(.A1(new_n757), .A2(G97), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n776), .B(new_n777), .C1(new_n259), .C2(new_n763), .ZN(new_n778));
  INV_X1    g0578(.A(new_n772), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n779), .A2(G50), .B1(G68), .B2(new_n752), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n256), .B1(new_n745), .B2(new_n507), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G107), .B2(new_n768), .ZN(new_n782));
  INV_X1    g0582(.A(new_n749), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n780), .B(new_n782), .C1(new_n378), .C2(new_n783), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n765), .A2(new_n774), .B1(new_n778), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n742), .B1(new_n785), .B2(new_n739), .ZN(new_n786));
  INV_X1    g0586(.A(new_n738), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n712), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT100), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n727), .A2(new_n789), .ZN(G396));
  AOI21_X1  g0590(.A(new_n647), .B1(new_n623), .B2(new_n637), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n361), .A2(new_n374), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n672), .B1(new_n357), .B2(new_n360), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n370), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n361), .A2(new_n368), .A3(new_n369), .A4(new_n672), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n791), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n791), .A2(new_n797), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n694), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n725), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n802), .B1(new_n804), .B2(KEYINPUT102), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(KEYINPUT102), .B2(new_n804), .ZN(new_n806));
  INV_X1    g0606(.A(new_n763), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G116), .ZN(new_n808));
  INV_X1    g0608(.A(new_n766), .ZN(new_n809));
  INV_X1    g0609(.A(new_n752), .ZN(new_n810));
  INV_X1    g0610(.A(G283), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n764), .A2(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G303), .B2(new_n779), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n265), .B1(new_n745), .B2(new_n205), .C1(new_n767), .C2(new_n507), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G294), .B2(new_n749), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n808), .A2(new_n777), .A3(new_n813), .A4(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n752), .A2(G150), .B1(new_n749), .B2(G143), .ZN(new_n817));
  INV_X1    g0617(.A(G137), .ZN(new_n818));
  INV_X1    g0618(.A(G159), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n817), .B1(new_n818), .B2(new_n772), .C1(new_n763), .C2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(KEYINPUT34), .ZN(new_n822));
  INV_X1    g0622(.A(new_n745), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n265), .B1(new_n823), .B2(G50), .ZN(new_n824));
  INV_X1    g0624(.A(G132), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n824), .B1(new_n379), .B2(new_n767), .C1(new_n809), .C2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G58), .B2(new_n757), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT34), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n820), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n816), .B1(new_n822), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT101), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n739), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n739), .A2(new_n736), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n725), .B1(new_n259), .B2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n832), .B(new_n834), .C1(new_n737), .C2(new_n797), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n806), .A2(new_n835), .ZN(G384));
  INV_X1    g0636(.A(new_n536), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n837), .A2(KEYINPUT35), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(KEYINPUT35), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n838), .A2(G116), .A3(new_n218), .A4(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT36), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n215), .A2(new_n259), .A3(new_n380), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n287), .B2(G68), .ZN(new_n843));
  OR3_X1    g0643(.A1(new_n843), .A2(new_n208), .A3(G13), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n717), .A2(G1), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n645), .B1(new_n443), .B2(new_n444), .ZN(new_n846));
  INV_X1    g0646(.A(new_n377), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n399), .B2(new_n382), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n427), .B1(new_n401), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n645), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n447), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n849), .B1(new_n442), .B2(new_n850), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n430), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n395), .A2(new_n396), .A3(new_n402), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n857), .A2(new_n426), .B1(new_n442), .B2(new_n850), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(new_n859), .A3(new_n430), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n856), .A2(new_n860), .A3(KEYINPUT104), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT104), .B1(new_n856), .B2(new_n860), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n853), .A2(KEYINPUT38), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT38), .B1(new_n853), .B2(new_n863), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n647), .B(new_n796), .C1(new_n623), .C2(new_n637), .ZN(new_n867));
  INV_X1    g0667(.A(new_n795), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT103), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT103), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n799), .A2(new_n870), .A3(new_n795), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n341), .A2(new_n672), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n340), .A2(new_n344), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n873), .B1(new_n336), .B2(new_n339), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n846), .B1(new_n866), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n853), .A2(new_n863), .A3(KEYINPUT38), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n439), .A2(new_n850), .ZN(new_n882));
  INV_X1    g0682(.A(new_n436), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n882), .B1(new_n883), .B2(new_n445), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n858), .A2(new_n430), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(new_n859), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n881), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n880), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT39), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n851), .B1(new_n606), .B2(new_n445), .ZN(new_n891));
  INV_X1    g0691(.A(new_n862), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n856), .A2(new_n860), .A3(KEYINPUT104), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n881), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(KEYINPUT39), .A3(new_n880), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n340), .A2(new_n647), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n879), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n707), .A2(new_n708), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n376), .A2(new_n448), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n611), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n900), .B(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT31), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n686), .A2(new_n691), .ZN(new_n906));
  OAI211_X1 g0706(.A(KEYINPUT105), .B(new_n905), .C1(new_n906), .C2(new_n672), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT105), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n692), .B2(KEYINPUT31), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n602), .A2(new_n672), .B1(KEYINPUT31), .B2(new_n692), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n796), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n877), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n864), .B2(new_n865), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT40), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n912), .A2(new_n877), .A3(KEYINPUT40), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n915), .A2(new_n916), .B1(new_n888), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n910), .A2(new_n911), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n450), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(G330), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n921), .B2(new_n919), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n845), .B1(new_n904), .B2(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n904), .A2(new_n923), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n841), .B(new_n844), .C1(new_n924), .C2(new_n925), .ZN(G367));
  INV_X1    g0726(.A(new_n723), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT45), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT109), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n542), .A2(new_n647), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n543), .A2(new_n547), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT107), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n629), .A2(new_n647), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n543), .A2(new_n547), .A3(KEYINPUT107), .A4(new_n930), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n929), .B1(new_n663), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n656), .A2(new_n647), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT90), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n601), .A2(new_n939), .A3(new_n654), .A4(new_n662), .ZN(new_n940));
  INV_X1    g0740(.A(new_n660), .ZN(new_n941));
  AND4_X1   g0741(.A1(new_n929), .A2(new_n936), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n928), .B1(new_n937), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT44), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n663), .A2(new_n936), .B1(KEYINPUT110), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n940), .A2(new_n941), .ZN(new_n946));
  INV_X1    g0746(.A(new_n936), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n944), .A2(KEYINPUT110), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n944), .A2(KEYINPUT110), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n945), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT109), .B1(new_n946), .B2(new_n947), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n663), .A2(new_n929), .A3(new_n936), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(new_n953), .A3(KEYINPUT45), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n943), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n659), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n481), .A2(new_n672), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n652), .B(new_n958), .C1(new_n655), .C2(new_n657), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT111), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n940), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n940), .A2(KEYINPUT111), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n715), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n655), .A2(new_n958), .A3(new_n657), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n959), .B2(new_n960), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n967), .A2(new_n651), .A3(new_n963), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n969), .A2(new_n709), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n943), .A2(new_n951), .A3(new_n954), .A4(new_n659), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n957), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT112), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n957), .A2(new_n970), .A3(KEYINPUT112), .A4(new_n971), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n709), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n666), .B(new_n977), .Z(new_n978));
  OAI21_X1  g0778(.A(new_n927), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n936), .A2(new_n966), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT42), .Z(new_n981));
  AOI21_X1  g0781(.A(new_n594), .B1(new_n933), .B2(new_n935), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n672), .B1(new_n982), .B2(new_n629), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n615), .B1(new_n510), .B2(new_n672), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n695), .A2(new_n613), .A3(new_n647), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT43), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n984), .B(new_n989), .C1(new_n990), .C2(new_n987), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n984), .B2(new_n989), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n659), .A2(new_n947), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n992), .B(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n979), .A2(new_n994), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n256), .B1(new_n745), .B2(new_n378), .C1(new_n767), .C2(new_n259), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n818), .A2(new_n809), .B1(new_n810), .B2(new_n819), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n996), .B(new_n997), .C1(G150), .C2(new_n749), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n758), .A2(new_n379), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n807), .B2(G50), .ZN(new_n1000));
  INV_X1    g0800(.A(G143), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n998), .B(new_n1000), .C1(new_n1001), .C2(new_n773), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n758), .A2(new_n205), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n823), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT46), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n745), .B2(new_n464), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1004), .B(new_n1006), .C1(new_n810), .C2(new_n559), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n1003), .B(new_n1007), .C1(new_n807), .C2(G283), .ZN(new_n1008));
  INV_X1    g0808(.A(G317), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n265), .B1(new_n204), .B2(new_n767), .C1(new_n809), .C2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT114), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT113), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n773), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1013), .A2(G311), .B1(G303), .B2(new_n749), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1008), .B(new_n1011), .C1(new_n1012), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1014), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1016), .A2(KEYINPUT113), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1002), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT47), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1020), .A2(new_n739), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n987), .A2(new_n738), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n731), .A2(new_n238), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n741), .B1(new_n665), .B2(new_n495), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n725), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1022), .A2(new_n1023), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n995), .A2(new_n1027), .ZN(G387));
  NAND2_X1  g0828(.A1(new_n807), .A2(G68), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n810), .A2(new_n281), .B1(new_n772), .B2(new_n819), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G150), .B2(new_n766), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n757), .A2(new_n495), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n823), .A2(G77), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1033), .B(new_n256), .C1(new_n204), .C2(new_n767), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G50), .B2(new_n749), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1029), .A2(new_n1031), .A3(new_n1032), .A4(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n256), .B1(new_n768), .B2(G116), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n752), .A2(G311), .B1(new_n749), .B2(G317), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n763), .B2(new_n746), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G322), .B2(new_n1013), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1040), .A2(KEYINPUT48), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(KEYINPUT48), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n758), .A2(new_n811), .B1(new_n559), .B2(new_n745), .ZN(new_n1043));
  OR3_X1    g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT49), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1037), .B1(new_n771), .B2(new_n809), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1036), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n739), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n347), .A2(new_n349), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n287), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT115), .Z(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(KEYINPUT50), .ZN(new_n1053));
  AOI21_X1  g0853(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1053), .A2(new_n668), .A3(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1052), .A2(KEYINPUT50), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n731), .B1(new_n718), .B2(new_n235), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(G107), .B2(new_n212), .C1(new_n668), .C2(new_n728), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n725), .B1(new_n1058), .B2(new_n740), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1049), .B(new_n1059), .C1(new_n658), .C2(new_n787), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n666), .B1(new_n969), .B2(new_n709), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n969), .A2(new_n709), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1060), .B1(new_n927), .B2(new_n969), .C1(new_n1061), .C2(new_n1062), .ZN(G393));
  NAND2_X1  g0863(.A1(new_n974), .A2(new_n975), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n970), .B1(new_n957), .B2(new_n971), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1065), .A2(new_n667), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n957), .A2(new_n723), .A3(new_n971), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n936), .A2(new_n787), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT116), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n807), .A2(G294), .B1(G116), .B2(new_n757), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1009), .A2(new_n772), .B1(new_n783), .B2(new_n764), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT52), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n265), .B1(new_n745), .B2(new_n811), .C1(new_n767), .C2(new_n205), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n810), .A2(new_n746), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(G322), .C2(new_n766), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1071), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n256), .B1(new_n745), .B2(new_n379), .C1(new_n767), .C2(new_n507), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n810), .A2(new_n287), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(G143), .C2(new_n766), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n807), .A2(new_n1050), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n757), .A2(G77), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n277), .A2(new_n772), .B1(new_n783), .B2(new_n819), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT51), .Z(new_n1085));
  OAI21_X1  g0885(.A(new_n1077), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n739), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n740), .B1(new_n204), .B2(new_n212), .C1(new_n732), .C2(new_n245), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1070), .A2(new_n724), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1068), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1067), .A2(new_n1091), .ZN(G390));
  NOR2_X1   g0892(.A1(new_n694), .A2(new_n796), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n913), .A2(new_n641), .B1(new_n877), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n920), .A2(G330), .A3(new_n797), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(new_n875), .A3(new_n876), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n706), .A2(new_n672), .A3(new_n794), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n795), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n1093), .B2(new_n877), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1094), .A2(new_n872), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n376), .A2(G330), .A3(new_n448), .A4(new_n920), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1101), .A2(new_n610), .A3(new_n902), .A4(new_n305), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n913), .A2(new_n641), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n899), .B1(new_n872), .B2(new_n877), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n864), .A2(new_n865), .A3(new_n889), .ZN(new_n1109));
  AOI21_X1  g0909(.A(KEYINPUT39), .B1(new_n880), .B2(new_n887), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n899), .B1(new_n877), .B2(new_n1098), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n888), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1106), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1107), .B1(new_n890), .B2(new_n896), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1113), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1093), .A2(new_n877), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n1115), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1104), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1111), .A2(new_n1113), .A3(new_n1117), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1105), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1121), .A2(new_n1122), .A3(new_n1103), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1120), .A2(new_n666), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1121), .A2(new_n1122), .A3(new_n723), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n833), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n724), .B1(new_n346), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n256), .B1(new_n767), .B2(new_n287), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n823), .A2(G150), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT53), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1128), .B(new_n1130), .C1(G132), .C2(new_n749), .ZN(new_n1131));
  INV_X1    g0931(.A(G128), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n810), .A2(new_n818), .B1(new_n772), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G125), .B2(new_n766), .ZN(new_n1134));
  XOR2_X1   g0934(.A(KEYINPUT54), .B(G143), .Z(new_n1135));
  NAND2_X1  g0935(.A1(new_n807), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n757), .A2(G159), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1131), .A2(new_n1134), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n807), .A2(G97), .ZN(new_n1139));
  INV_X1    g0939(.A(G294), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n809), .A2(new_n1140), .B1(new_n772), .B2(new_n811), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G107), .B2(new_n752), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n265), .B1(new_n745), .B2(new_n507), .C1(new_n767), .C2(new_n379), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G116), .B2(new_n749), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1139), .A2(new_n1082), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1138), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1127), .B1(new_n1146), .B2(new_n739), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n898), .B2(new_n737), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1125), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1124), .A2(new_n1149), .ZN(G378));
  INV_X1    g0950(.A(new_n899), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n846), .B1(new_n866), .B2(new_n878), .C1(new_n897), .C2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n292), .A2(new_n850), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n306), .B(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1154), .B(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n918), .B2(G330), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n888), .A2(new_n917), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n913), .B1(new_n895), .B2(new_n880), .ZN(new_n1159));
  OAI211_X1 g0959(.A(G330), .B(new_n1158), .C1(new_n1159), .C2(KEYINPUT40), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1154), .B(new_n1155), .Z(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1152), .B1(new_n1157), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n918), .A2(G330), .A3(new_n1156), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n900), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1161), .A2(new_n736), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n724), .B1(G50), .B2(new_n1126), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n256), .A2(G41), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1033), .B(new_n1170), .C1(new_n378), .C2(new_n767), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1171), .B(new_n999), .C1(G107), .C2(new_n749), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n809), .A2(new_n811), .B1(new_n772), .B2(new_n464), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G97), .B2(new_n752), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1172), .B(new_n1174), .C1(new_n351), .C2(new_n763), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT58), .ZN(new_n1176));
  INV_X1    g0976(.A(G41), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n261), .B2(new_n263), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1175), .A2(new_n1176), .B1(new_n287), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n766), .A2(G124), .ZN(new_n1180));
  AOI211_X1 g0980(.A(G33), .B(G41), .C1(new_n768), .C2(G159), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n749), .A2(G128), .B1(new_n823), .B2(new_n1135), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n825), .B2(new_n810), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n763), .A2(new_n818), .B1(new_n277), .B2(new_n758), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(G125), .C2(new_n779), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT59), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1180), .B(new_n1181), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1179), .B1(new_n1176), .B2(new_n1175), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1169), .B1(new_n1189), .B2(new_n739), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1167), .A2(new_n723), .B1(new_n1168), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1102), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1163), .A2(new_n1166), .B1(new_n1123), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n666), .B1(new_n1193), .B2(KEYINPUT57), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1123), .A2(new_n1192), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1167), .A2(KEYINPUT57), .A3(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1191), .B1(new_n1194), .B2(new_n1196), .ZN(G375));
  INV_X1    g0997(.A(new_n978), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1104), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n724), .B1(G68), .B2(new_n1126), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n772), .A2(new_n1140), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n265), .B1(new_n259), .B2(new_n767), .C1(new_n783), .C2(new_n811), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(G116), .C2(new_n752), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n766), .A2(G303), .B1(G97), .B2(new_n823), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT117), .Z(new_n1206));
  NAND2_X1  g1006(.A1(new_n807), .A2(G107), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n1032), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n265), .B1(new_n768), .B2(G58), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n819), .B2(new_n745), .C1(new_n809), .C2(new_n1132), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n807), .B2(G150), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n752), .A2(new_n1135), .B1(new_n749), .B2(G137), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n825), .B2(new_n772), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT118), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1211), .B(new_n1215), .C1(new_n287), .C2(new_n758), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1208), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1201), .B1(new_n1218), .B2(new_n739), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n877), .B2(new_n737), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n1100), .B2(new_n927), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1200), .A2(new_n1222), .ZN(G381));
  INV_X1    g1023(.A(G375), .ZN(new_n1224));
  INV_X1    g1024(.A(G378), .ZN(new_n1225));
  OR3_X1    g1025(.A1(G384), .A2(G393), .A3(G396), .ZN(new_n1226));
  NOR4_X1   g1026(.A1(G387), .A2(new_n1226), .A3(G390), .A4(G381), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1227), .ZN(G407));
  NAND2_X1  g1028(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1229));
  OAI211_X1 g1029(.A(G407), .B(G213), .C1(new_n1229), .C2(G343), .ZN(G409));
  INV_X1    g1030(.A(G213), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1231), .A2(G343), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(G2897), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(KEYINPUT60), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1199), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT120), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT120), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1235), .A2(new_n1238), .A3(new_n1199), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1199), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n667), .B1(new_n1240), .B2(KEYINPUT60), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1237), .A2(new_n1239), .A3(new_n1241), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1242), .A2(G384), .A3(new_n1222), .ZN(new_n1243));
  AOI21_X1  g1043(.A(G384), .B1(new_n1242), .B2(new_n1222), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1234), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1222), .ZN(new_n1246));
  INV_X1    g1046(.A(G384), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1242), .A2(G384), .A3(new_n1222), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n1249), .A3(new_n1233), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1245), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(G375), .A2(G378), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1167), .A2(new_n1198), .A3(new_n1195), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1168), .A2(new_n1190), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1124), .A2(new_n1149), .A3(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT119), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1167), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1163), .A2(KEYINPUT119), .A3(new_n1166), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n723), .A3(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1232), .B1(new_n1256), .B2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1251), .B1(new_n1252), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT121), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n667), .B(new_n1065), .C1(new_n974), .C2(new_n975), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1263), .B1(new_n1264), .B2(new_n1090), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1067), .A2(KEYINPUT121), .A3(new_n1091), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1027), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(new_n979), .B2(new_n994), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT122), .B1(new_n1267), .B2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT121), .B1(new_n1067), .B2(new_n1091), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1263), .B(new_n1090), .C1(new_n1064), .C2(new_n1066), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT122), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(G387), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  XOR2_X1   g1075(.A(G393), .B(G396), .Z(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(new_n1269), .B2(G390), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1270), .A2(new_n1275), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT123), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1270), .A2(new_n1275), .A3(new_n1277), .A4(KEYINPUT123), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1269), .B(G390), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1280), .A2(new_n1281), .B1(new_n1276), .B2(new_n1282), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1262), .A2(new_n1283), .A3(KEYINPUT61), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1252), .A2(new_n1261), .A3(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT63), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1252), .A2(new_n1261), .A3(KEYINPUT63), .A4(new_n1285), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1284), .A2(KEYINPUT124), .A3(new_n1288), .A4(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT124), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1245), .A2(new_n1250), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1193), .A2(new_n1198), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1225), .A2(new_n1254), .A3(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1260), .ZN(new_n1296));
  OAI22_X1  g1096(.A1(new_n1295), .A2(new_n1296), .B1(new_n1231), .B2(G343), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1167), .A2(new_n1195), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT57), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1193), .A2(KEYINPUT57), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(new_n666), .A3(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1225), .B1(new_n1302), .B2(new_n1191), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1293), .B1(new_n1297), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1282), .A2(new_n1276), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT61), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1304), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1291), .B1(new_n1292), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1290), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1304), .A2(new_n1308), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT62), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1286), .A2(KEYINPUT125), .A3(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(KEYINPUT125), .B1(new_n1286), .B2(new_n1313), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1252), .A2(new_n1261), .A3(KEYINPUT62), .A4(new_n1285), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT126), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(new_n1317), .B(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1312), .B1(new_n1316), .B2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1311), .B1(new_n1320), .B2(new_n1307), .ZN(G405));
  NAND2_X1  g1121(.A1(new_n1285), .A2(KEYINPUT127), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1283), .B(new_n1322), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1229), .B(new_n1252), .C1(KEYINPUT127), .C2(new_n1285), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1323), .B(new_n1324), .ZN(G402));
endmodule


