//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n981, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(KEYINPUT102), .ZN(new_n202));
  XNOR2_X1  g001(.A(G183gat), .B(G211gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n204));
  XNOR2_X1  g003(.A(G127gat), .B(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G57gat), .B(G64gat), .Z(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT96), .ZN(new_n208));
  XNOR2_X1  g007(.A(G57gat), .B(G64gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT96), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(G71gat), .A2(G78gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT9), .ZN(new_n214));
  NAND2_X1  g013(.A1(G71gat), .A2(G78gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n213), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(new_n215), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n219), .B1(new_n207), .B2(KEYINPUT9), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G231gat), .A2(G233gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT97), .B(KEYINPUT21), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n223), .B1(new_n222), .B2(new_n224), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n206), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NOR3_X1   g028(.A1(new_n226), .A2(new_n227), .A3(new_n206), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n204), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n230), .ZN(new_n232));
  INV_X1    g031(.A(new_n204), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(new_n228), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n203), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G15gat), .B(G22gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT16), .ZN(new_n238));
  AOI21_X1  g037(.A(G1gat), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT93), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n237), .B(new_n240), .C1(new_n238), .C2(G1gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(G8gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT21), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n246), .B1(new_n247), .B2(new_n222), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n248), .B(KEYINPUT98), .Z(new_n249));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n234), .A3(new_n203), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n236), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n249), .ZN(new_n252));
  INV_X1    g051(.A(new_n250), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(new_n253), .B2(new_n235), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G232gat), .A2(G233gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n258), .A2(KEYINPUT41), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT99), .ZN(new_n260));
  XOR2_X1   g059(.A(G134gat), .B(G162gat), .Z(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G99gat), .A2(G106gat), .ZN(new_n263));
  INV_X1    g062(.A(G85gat), .ZN(new_n264));
  INV_X1    g063(.A(G92gat), .ZN(new_n265));
  AOI22_X1  g064(.A1(KEYINPUT8), .A2(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT7), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n267), .B1(new_n264), .B2(new_n265), .ZN(new_n268));
  NAND3_X1  g067(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(G99gat), .B(G106gat), .Z(new_n271));
  OR2_X1    g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT100), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n271), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n273), .B1(new_n272), .B2(new_n274), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT14), .ZN(new_n279));
  INV_X1    g078(.A(G29gat), .ZN(new_n280));
  INV_X1    g079(.A(G36gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT89), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT89), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n284), .A2(new_n279), .A3(new_n280), .A4(new_n281), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT90), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n287), .A2(new_n288), .B1(G29gat), .B2(G36gat), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n283), .A2(new_n285), .A3(KEYINPUT90), .A4(new_n286), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G43gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G50gat), .ZN(new_n293));
  INV_X1    g092(.A(G50gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G43gat), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n293), .A2(new_n295), .A3(KEYINPUT15), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n296), .B1(G29gat), .B2(G36gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT91), .B(G43gat), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n293), .B1(new_n299), .B2(G50gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT15), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n282), .A2(new_n286), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n304), .B(KEYINPUT92), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n297), .A2(new_n306), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n278), .A2(new_n307), .B1(KEYINPUT41), .B2(new_n258), .ZN(new_n308));
  XNOR2_X1  g107(.A(G190gat), .B(G218gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT17), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT94), .B1(new_n307), .B2(new_n311), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n296), .A2(new_n291), .B1(new_n303), .B2(new_n305), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT94), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT17), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n278), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n318), .B1(new_n313), .B2(KEYINPUT17), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n308), .B(new_n310), .C1(new_n317), .C2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT101), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n262), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n319), .B1(new_n312), .B2(new_n315), .ZN(new_n323));
  INV_X1    g122(.A(new_n308), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n309), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n320), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n325), .B(new_n320), .C1(new_n321), .C2(new_n262), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n202), .B1(new_n256), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n255), .A2(new_n329), .A3(KEYINPUT102), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G230gat), .A2(G233gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n217), .A2(KEYINPUT10), .A3(new_n221), .ZN(new_n335));
  NOR3_X1   g134(.A1(new_n276), .A2(new_n335), .A3(new_n277), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n208), .A2(new_n211), .B1(new_n215), .B2(new_n214), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n337), .A2(new_n220), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n272), .A2(new_n274), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n272), .B(new_n274), .C1(new_n337), .C2(new_n220), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT10), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n334), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n341), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n343), .B1(new_n334), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G120gat), .B(G148gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(G176gat), .B(G204gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n345), .A2(new_n348), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n333), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT88), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n246), .A2(new_n313), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n307), .A2(new_n245), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G229gat), .A2(G233gat), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n359), .B(KEYINPUT13), .Z(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n245), .B1(new_n307), .B2(new_n311), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n307), .A2(KEYINPUT94), .A3(new_n311), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n314), .B1(new_n313), .B2(KEYINPUT17), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n365), .A2(new_n359), .A3(new_n357), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT18), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n361), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n316), .A2(new_n362), .B1(new_n307), .B2(new_n245), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT18), .B1(new_n369), .B2(new_n359), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n355), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G113gat), .B(G141gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(KEYINPUT11), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(G169gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT87), .B(G197gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT12), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n371), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n366), .A2(new_n367), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n369), .A2(KEYINPUT18), .A3(new_n359), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n381), .A3(new_n361), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(new_n355), .A3(new_n377), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT84), .ZN(new_n386));
  AND2_X1   g185(.A1(G141gat), .A2(G148gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(G141gat), .A2(G148gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G155gat), .B(G162gat), .ZN(new_n390));
  INV_X1    g189(.A(G155gat), .ZN(new_n391));
  INV_X1    g190(.A(G162gat), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT2), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n389), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(G134gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(G127gat), .ZN(new_n396));
  INV_X1    g195(.A(G127gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G134gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G113gat), .B(G120gat), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n399), .B1(new_n400), .B2(KEYINPUT1), .ZN(new_n401));
  INV_X1    g200(.A(G120gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(G113gat), .ZN(new_n403));
  INV_X1    g202(.A(G113gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(G120gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G127gat), .B(G134gat), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT1), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(G141gat), .ZN(new_n410));
  INV_X1    g209(.A(G148gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT2), .ZN(new_n413));
  NAND2_X1  g212(.A1(G141gat), .A2(G148gat), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  AND2_X1   g214(.A1(G155gat), .A2(G162gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(G155gat), .A2(G162gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n394), .A2(new_n401), .A3(new_n409), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT4), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT79), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n401), .A2(new_n409), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n394), .A2(new_n419), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT4), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT78), .A4(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT78), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(new_n420), .B2(KEYINPUT4), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT79), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n420), .A2(new_n429), .A3(KEYINPUT4), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n422), .A2(new_n426), .A3(new_n428), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n394), .A2(new_n419), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT3), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n401), .A2(new_n409), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT3), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n394), .A2(new_n419), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(G225gat), .A2(G233gat), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n439), .A2(KEYINPUT5), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n431), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n425), .B1(new_n423), .B2(new_n424), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n420), .A2(KEYINPUT4), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n438), .B(new_n437), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT5), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n434), .A2(new_n432), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT76), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT76), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n434), .A2(new_n432), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n438), .B1(new_n450), .B2(new_n420), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n445), .A2(new_n451), .A3(KEYINPUT77), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT77), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT5), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n439), .B1(new_n455), .B2(new_n421), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n454), .B1(new_n456), .B2(new_n437), .ZN(new_n457));
  INV_X1    g256(.A(new_n449), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n448), .B1(new_n434), .B2(new_n432), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n420), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n439), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n453), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n441), .B1(new_n452), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G1gat), .B(G29gat), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT0), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(G57gat), .B(G85gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n463), .A2(KEYINPUT6), .A3(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n468), .B(new_n441), .C1(new_n452), .C2(new_n462), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT81), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n468), .B(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT77), .B1(new_n445), .B2(new_n451), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n457), .A2(new_n453), .A3(new_n461), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n476), .B1(new_n479), .B2(new_n441), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n470), .B1(new_n473), .B2(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(G211gat), .B(G218gat), .Z(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(G197gat), .B(G204gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT71), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n485), .B1(new_n484), .B2(new_n487), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n483), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(G204gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(G197gat), .ZN(new_n493));
  INV_X1    g292(.A(G197gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(G204gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT71), .B1(new_n496), .B2(new_n486), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(new_n482), .A3(new_n488), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n491), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(G226gat), .A2(G233gat), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT25), .ZN(new_n503));
  NAND2_X1  g302(.A1(G169gat), .A2(G176gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT23), .ZN(new_n505));
  INV_X1    g304(.A(G169gat), .ZN(new_n506));
  INV_X1    g305(.A(G176gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT23), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G183gat), .A2(G190gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT24), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT24), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(G183gat), .A3(G190gat), .ZN(new_n515));
  INV_X1    g314(.A(G183gat), .ZN(new_n516));
  INV_X1    g315(.A(G190gat), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n513), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g317(.A(KEYINPUT64), .B(new_n503), .C1(new_n511), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n516), .A2(KEYINPUT65), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT65), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G183gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n522), .A3(new_n517), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n514), .B1(G183gat), .B2(G190gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n512), .A2(KEYINPUT24), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT23), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n527), .A2(G169gat), .A3(G176gat), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n528), .B1(new_n508), .B2(new_n505), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(new_n529), .A3(KEYINPUT25), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n519), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n517), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(new_n524), .B2(new_n525), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT64), .B1(new_n534), .B2(new_n503), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT27), .B(G183gat), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n536), .A2(KEYINPUT28), .A3(new_n517), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT27), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n538), .B1(new_n520), .B2(new_n522), .ZN(new_n539));
  NOR2_X1   g338(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n517), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT28), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n537), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT26), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n504), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n508), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n546), .B1(KEYINPUT26), .B2(new_n508), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n512), .ZN(new_n548));
  OAI22_X1  g347(.A1(new_n531), .A2(new_n535), .B1(new_n543), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT72), .B(KEYINPUT29), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n502), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n503), .B1(new_n511), .B2(new_n518), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT64), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(new_n519), .A3(new_n530), .ZN(new_n555));
  INV_X1    g354(.A(new_n540), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT65), .B(G183gat), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n556), .B1(new_n557), .B2(new_n538), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT28), .B1(new_n558), .B2(new_n517), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n512), .B(new_n547), .C1(new_n559), .C2(new_n537), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n501), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n500), .B1(new_n551), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT37), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n549), .A2(new_n502), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT29), .B1(new_n555), .B2(new_n560), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n564), .B(new_n499), .C1(new_n565), .C2(new_n502), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n499), .B1(new_n551), .B2(new_n561), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n564), .B(new_n500), .C1(new_n565), .C2(new_n502), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(KEYINPUT37), .A3(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G8gat), .B(G36gat), .Z(new_n571));
  XNOR2_X1  g370(.A(G64gat), .B(G92gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT73), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(KEYINPUT38), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n567), .A2(new_n570), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n562), .A2(new_n566), .A3(new_n573), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT75), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n562), .A2(KEYINPUT75), .A3(new_n566), .A4(new_n573), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n386), .B1(new_n481), .B2(new_n581), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n463), .A2(new_n475), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(new_n472), .A3(new_n471), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n583), .A2(KEYINPUT84), .A3(new_n470), .A4(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n567), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n587), .A2(new_n573), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n563), .B1(new_n562), .B2(new_n566), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT38), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n582), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(G228gat), .ZN(new_n592));
  INV_X1    g391(.A(G233gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n550), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n595), .B1(new_n491), .B2(new_n498), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n432), .B1(new_n596), .B2(KEYINPUT3), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n436), .A2(new_n550), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n500), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n594), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT29), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n497), .A2(new_n482), .A3(new_n488), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n482), .B1(new_n497), .B2(new_n488), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n424), .B1(new_n604), .B2(new_n435), .ZN(new_n605));
  INV_X1    g404(.A(new_n598), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n594), .B1(new_n499), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(G22gat), .B1(new_n600), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n550), .B1(new_n602), .B2(new_n603), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n424), .B1(new_n610), .B2(new_n435), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n499), .A2(new_n606), .ZN(new_n612));
  OAI22_X1  g411(.A1(new_n611), .A2(new_n612), .B1(new_n592), .B2(new_n593), .ZN(new_n613));
  INV_X1    g412(.A(G22gat), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT29), .B1(new_n491), .B2(new_n498), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n432), .B1(new_n615), .B2(KEYINPUT3), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(new_n594), .A3(new_n599), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n613), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT80), .B(KEYINPUT31), .Z(new_n619));
  AND3_X1   g418(.A1(new_n609), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n619), .B1(new_n609), .B2(new_n618), .ZN(new_n621));
  XNOR2_X1  g420(.A(G78gat), .B(G106gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(new_n294), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n620), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n619), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n600), .A2(new_n608), .A3(G22gat), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n614), .B1(new_n613), .B2(new_n617), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n609), .A2(new_n618), .A3(new_n619), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n623), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT82), .ZN(new_n633));
  AOI211_X1 g432(.A(KEYINPUT39), .B(new_n438), .C1(new_n431), .C2(new_n437), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n634), .B2(new_n475), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n438), .B(new_n420), .C1(new_n458), .C2(new_n459), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n636), .B1(new_n637), .B2(KEYINPUT83), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT83), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n450), .A2(new_n639), .A3(new_n438), .A4(new_n420), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n431), .A2(new_n437), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n439), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI211_X1 g443(.A(KEYINPUT82), .B(new_n476), .C1(new_n643), .C2(KEYINPUT39), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n635), .A2(new_n644), .A3(new_n645), .A4(KEYINPUT40), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n584), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n438), .B1(new_n431), .B2(new_n437), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n475), .B1(new_n648), .B2(new_n636), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n649), .A2(KEYINPUT82), .B1(new_n641), .B2(new_n643), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT40), .B1(new_n650), .B2(new_n635), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT30), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n579), .A2(new_n653), .A3(new_n580), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n562), .A2(new_n566), .ZN(new_n655));
  INV_X1    g454(.A(new_n574), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n562), .A2(KEYINPUT30), .A3(new_n566), .A4(new_n573), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT74), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n654), .B(new_n657), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n632), .B1(new_n652), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n591), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT85), .ZN(new_n665));
  INV_X1    g464(.A(new_n470), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n463), .A2(new_n469), .ZN(new_n667));
  INV_X1    g466(.A(new_n473), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n662), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n632), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT70), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT67), .B(KEYINPUT34), .Z(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n549), .A2(new_n423), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n555), .A2(new_n434), .A3(new_n560), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(G227gat), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n593), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n676), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  AOI211_X1 g482(.A(new_n681), .B(new_n675), .C1(new_n677), .C2(new_n678), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n677), .A2(new_n681), .A3(new_n678), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT33), .ZN(new_n687));
  XNOR2_X1  g486(.A(G15gat), .B(G43gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT66), .ZN(new_n689));
  XNOR2_X1  g488(.A(G71gat), .B(G99gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n686), .B(KEYINPUT32), .C1(new_n687), .C2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n686), .A2(KEYINPUT32), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n686), .A2(new_n687), .ZN(new_n694));
  INV_X1    g493(.A(new_n691), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n685), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n685), .A2(new_n696), .A3(new_n692), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT68), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n685), .A2(new_n696), .A3(KEYINPUT68), .A4(new_n692), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n697), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n674), .B1(new_n702), .B2(KEYINPUT36), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n701), .ZN(new_n704));
  INV_X1    g503(.A(new_n697), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT36), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n706), .A2(KEYINPUT70), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT69), .ZN(new_n709));
  AND4_X1   g508(.A1(new_n709), .A2(new_n704), .A3(KEYINPUT36), .A4(new_n705), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n702), .B2(KEYINPUT36), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n703), .B(new_n708), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT85), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n591), .A2(new_n663), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n665), .A2(new_n673), .A3(new_n712), .A4(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT86), .ZN(new_n716));
  INV_X1    g515(.A(new_n632), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n702), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT35), .B1(new_n672), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT35), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n717), .A2(new_n720), .A3(new_n671), .A4(new_n481), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n706), .B2(new_n721), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n715), .A2(new_n716), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n716), .B1(new_n715), .B2(new_n722), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n385), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT95), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g526(.A(KEYINPUT95), .B(new_n385), .C1(new_n723), .C2(new_n724), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n354), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n669), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G1gat), .ZN(G1324gat));
  INV_X1    g530(.A(KEYINPUT103), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n662), .ZN(new_n733));
  XNOR2_X1  g532(.A(KEYINPUT16), .B(G8gat), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n735), .A2(KEYINPUT42), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(KEYINPUT42), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n733), .A2(G8gat), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(G1325gat));
  AOI21_X1  g538(.A(G15gat), .B1(new_n729), .B2(new_n702), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n740), .A2(KEYINPUT104), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(KEYINPUT104), .ZN(new_n743));
  INV_X1    g542(.A(new_n712), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n729), .A2(G15gat), .A3(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n741), .A2(new_n742), .A3(new_n743), .A4(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n740), .B2(KEYINPUT104), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n748));
  AOI211_X1 g547(.A(new_n748), .B(G15gat), .C1(new_n729), .C2(new_n702), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT105), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n746), .A2(new_n750), .ZN(G1326gat));
  NAND2_X1  g550(.A1(new_n729), .A2(new_n632), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT106), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n729), .A2(new_n754), .A3(new_n632), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT43), .B(G22gat), .Z(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT107), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n756), .B(new_n758), .ZN(G1327gat));
  NOR2_X1   g558(.A1(new_n255), .A2(new_n352), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(new_n329), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n727), .B2(new_n728), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n764), .A2(new_n280), .A3(new_n669), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n715), .A2(new_n722), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT86), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n715), .A2(new_n716), .A3(new_n722), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n772), .A2(KEYINPUT44), .A3(new_n330), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n329), .B1(new_n715), .B2(new_n722), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n774), .A2(KEYINPUT44), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n384), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(G29gat), .B1(new_n778), .B2(new_n670), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n767), .A2(new_n768), .A3(new_n779), .ZN(G1328gat));
  OAI21_X1  g579(.A(G36gat), .B1(new_n778), .B2(new_n671), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n671), .A2(G36gat), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n764), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n764), .A2(KEYINPUT108), .A3(new_n782), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n785), .A2(KEYINPUT46), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT46), .B1(new_n785), .B2(new_n786), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n781), .B1(new_n787), .B2(new_n788), .ZN(G1329gat));
  AOI21_X1  g588(.A(KEYINPUT95), .B1(new_n772), .B2(new_n385), .ZN(new_n790));
  INV_X1    g589(.A(new_n728), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n762), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n299), .B1(new_n792), .B2(new_n706), .ZN(new_n793));
  INV_X1    g592(.A(new_n299), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n744), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n778), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g596(.A(KEYINPUT109), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n717), .B1(new_n792), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n764), .A2(KEYINPUT109), .ZN(new_n800));
  AOI21_X1  g599(.A(G50gat), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n776), .A2(G50gat), .A3(new_n632), .A4(new_n777), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT48), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n632), .B1(new_n764), .B2(KEYINPUT109), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n792), .A2(new_n798), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n294), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT48), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n808), .A3(new_n802), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n804), .A2(new_n809), .ZN(G1331gat));
  AND3_X1   g609(.A1(new_n333), .A2(new_n384), .A3(new_n352), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n769), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT110), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n669), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n662), .ZN(new_n816));
  NOR2_X1   g615(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n817));
  AND2_X1   g616(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n817), .B2(new_n816), .ZN(G1333gat));
  NAND2_X1  g619(.A1(new_n813), .A2(new_n744), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n706), .A2(G71gat), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n821), .A2(G71gat), .B1(new_n813), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g623(.A1(new_n813), .A2(new_n632), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g625(.A1(new_n774), .A2(new_n384), .A3(new_n256), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT111), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n827), .A2(new_n828), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n829), .A2(KEYINPUT111), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n669), .A2(new_n264), .A3(new_n352), .ZN(new_n835));
  XOR2_X1   g634(.A(new_n835), .B(KEYINPUT112), .Z(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n385), .A2(new_n255), .A3(new_n353), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n776), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n839), .A2(new_n669), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n837), .B1(new_n840), .B2(new_n264), .ZN(G1336gat));
  NOR3_X1   g640(.A1(new_n671), .A2(G92gat), .A3(new_n353), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n834), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n776), .A2(new_n662), .A3(new_n838), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(G92gat), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n827), .B(new_n828), .ZN(new_n848));
  AOI22_X1  g647(.A1(new_n844), .A2(G92gat), .B1(new_n848), .B2(new_n842), .ZN(new_n849));
  OAI22_X1  g648(.A1(new_n843), .A2(new_n847), .B1(new_n849), .B2(new_n846), .ZN(G1337gat));
  INV_X1    g649(.A(G99gat), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n834), .A2(new_n851), .A3(new_n702), .A4(new_n352), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n839), .A2(new_n744), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n851), .ZN(G1338gat));
  NOR3_X1   g653(.A1(new_n717), .A2(new_n353), .A3(G106gat), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(new_n832), .B2(new_n833), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n773), .A2(new_n632), .A3(new_n775), .A4(new_n838), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(G106gat), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT113), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n856), .A2(new_n858), .A3(KEYINPUT113), .A4(new_n859), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n855), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT53), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n862), .A2(new_n863), .A3(new_n866), .ZN(G1339gat));
  INV_X1    g666(.A(KEYINPUT55), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n343), .A2(KEYINPUT54), .ZN(new_n869));
  OR3_X1    g668(.A1(new_n276), .A2(new_n335), .A3(new_n277), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT10), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n344), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n334), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT114), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n336), .A2(new_n342), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(KEYINPUT114), .A3(new_n873), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n869), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n348), .B1(new_n343), .B2(KEYINPUT54), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n868), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n870), .A2(new_n872), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n334), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT114), .B1(new_n877), .B2(new_n873), .ZN(new_n885));
  NOR4_X1   g684(.A1(new_n336), .A2(new_n342), .A3(new_n875), .A4(new_n334), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n880), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(KEYINPUT55), .A3(new_n888), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n881), .A2(new_n350), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n379), .A2(new_n890), .A3(new_n383), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n369), .A2(new_n359), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n358), .A2(new_n360), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n376), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n894), .B(new_n352), .C1(new_n382), .C2(new_n378), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n330), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n890), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n894), .B1(new_n382), .B2(new_n378), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n897), .A2(new_n898), .A3(new_n329), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n256), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n331), .A2(new_n384), .A3(new_n332), .A4(new_n353), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n718), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n670), .A2(new_n662), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n904), .A2(new_n384), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(new_n404), .ZN(G1340gat));
  NOR2_X1   g705(.A1(new_n904), .A2(new_n353), .ZN(new_n907));
  XOR2_X1   g706(.A(KEYINPUT115), .B(G120gat), .Z(new_n908));
  XNOR2_X1  g707(.A(new_n907), .B(new_n908), .ZN(G1341gat));
  NOR2_X1   g708(.A1(new_n904), .A2(new_n256), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(new_n397), .ZN(G1342gat));
  AOI21_X1  g710(.A(new_n670), .B1(new_n900), .B2(new_n901), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n329), .A2(new_n662), .ZN(new_n913));
  AND4_X1   g712(.A1(new_n702), .A2(new_n912), .A3(new_n717), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n395), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n915), .A2(KEYINPUT56), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT116), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n914), .A2(new_n395), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n918), .B1(KEYINPUT56), .B2(new_n915), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT117), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT117), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n917), .A2(new_n922), .A3(new_n919), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1343gat));
  AND3_X1   g723(.A1(new_n887), .A2(KEYINPUT118), .A3(new_n888), .ZN(new_n925));
  AOI21_X1  g724(.A(KEYINPUT118), .B1(new_n887), .B2(new_n888), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n868), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n889), .A2(new_n350), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n379), .A2(new_n927), .A3(new_n383), .A4(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n330), .B1(new_n929), .B2(new_n895), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n256), .B1(new_n930), .B2(new_n899), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n717), .B1(new_n931), .B2(new_n901), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n932), .A2(KEYINPUT57), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n717), .B1(new_n900), .B2(new_n901), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n934), .A2(KEYINPUT57), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n712), .B(new_n903), .C1(new_n933), .C2(new_n935), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n936), .A2(new_n384), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G141gat), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT119), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n912), .A2(new_n632), .A3(new_n712), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n384), .A2(G141gat), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n671), .ZN(new_n942));
  OAI22_X1  g741(.A1(new_n938), .A2(new_n939), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT119), .B1(new_n937), .B2(G141gat), .ZN(new_n944));
  OAI21_X1  g743(.A(KEYINPUT58), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT58), .ZN(new_n946));
  INV_X1    g745(.A(new_n941), .ZN(new_n947));
  XOR2_X1   g746(.A(new_n940), .B(KEYINPUT120), .Z(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n671), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n938), .B(new_n946), .C1(new_n947), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n945), .A2(new_n950), .ZN(G1344gat));
  NAND2_X1  g750(.A1(new_n712), .A2(new_n903), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT121), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n900), .A2(new_n901), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n954), .A2(new_n955), .A3(KEYINPUT57), .A4(new_n632), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n956), .B1(new_n932), .B2(KEYINPUT57), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n955), .B1(new_n934), .B2(KEYINPUT57), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n352), .B(new_n953), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n959), .A2(KEYINPUT123), .ZN(new_n960));
  OAI21_X1  g759(.A(G148gat), .B1(new_n959), .B2(KEYINPUT123), .ZN(new_n961));
  OAI21_X1  g760(.A(KEYINPUT59), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g763(.A(KEYINPUT124), .B(KEYINPUT59), .C1(new_n960), .C2(new_n961), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n411), .A2(KEYINPUT59), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n966), .B1(new_n936), .B2(new_n353), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n948), .A2(new_n411), .A3(new_n671), .A4(new_n352), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(G1345gat));
  OAI21_X1  g769(.A(G155gat), .B1(new_n936), .B2(new_n256), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n255), .A2(new_n391), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n949), .B2(new_n972), .ZN(G1346gat));
  NAND3_X1  g772(.A1(new_n948), .A2(new_n392), .A3(new_n913), .ZN(new_n974));
  OAI21_X1  g773(.A(G162gat), .B1(new_n936), .B2(new_n329), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1347gat));
  NOR2_X1   g775(.A1(new_n671), .A2(new_n669), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n902), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n978), .A2(new_n384), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(new_n506), .ZN(G1348gat));
  NOR2_X1   g779(.A1(new_n978), .A2(new_n353), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n981), .B(new_n507), .ZN(G1349gat));
  NOR2_X1   g781(.A1(new_n978), .A2(new_n256), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(new_n536), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n984), .B1(new_n557), .B2(new_n983), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g785(.A1(new_n902), .A2(new_n330), .A3(new_n977), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(G190gat), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT61), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n989), .B1(G190gat), .B2(new_n987), .ZN(G1351gat));
  XNOR2_X1  g789(.A(KEYINPUT125), .B(G197gat), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n712), .A2(new_n977), .ZN(new_n992));
  INV_X1    g791(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n993), .B1(new_n957), .B2(new_n958), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n991), .B1(new_n994), .B2(new_n384), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n934), .A2(new_n993), .ZN(new_n996));
  OR2_X1    g795(.A1(new_n384), .A2(new_n991), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(G1352gat));
  OAI21_X1  g797(.A(new_n352), .B1(new_n957), .B2(new_n958), .ZN(new_n999));
  OAI21_X1  g798(.A(G204gat), .B1(new_n999), .B2(new_n992), .ZN(new_n1000));
  NOR3_X1   g799(.A1(new_n996), .A2(G204gat), .A3(new_n353), .ZN(new_n1001));
  XNOR2_X1  g800(.A(new_n1001), .B(KEYINPUT62), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1000), .A2(new_n1002), .ZN(G1353gat));
  OR3_X1    g802(.A1(new_n996), .A2(G211gat), .A3(new_n256), .ZN(new_n1004));
  OAI211_X1 g803(.A(new_n255), .B(new_n993), .C1(new_n957), .C2(new_n958), .ZN(new_n1005));
  AND3_X1   g804(.A1(new_n1005), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1006));
  AOI21_X1  g805(.A(KEYINPUT63), .B1(new_n1005), .B2(G211gat), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g807(.A(new_n1008), .B(KEYINPUT126), .ZN(G1354gat));
  OAI21_X1  g808(.A(G218gat), .B1(new_n994), .B2(new_n329), .ZN(new_n1010));
  OR3_X1    g809(.A1(new_n996), .A2(G218gat), .A3(new_n329), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g811(.A(new_n1012), .B(KEYINPUT127), .Z(G1355gat));
endmodule


