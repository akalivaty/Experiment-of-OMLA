//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT68), .ZN(new_n188));
  XOR2_X1   g002(.A(KEYINPUT2), .B(G113), .Z(new_n189));
  XNOR2_X1  g003(.A(G116), .B(G119), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G116), .ZN(new_n193));
  INV_X1    g007(.A(G116), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT2), .B(G113), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n188), .B1(new_n191), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n189), .A2(new_n190), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n196), .A2(new_n197), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(KEYINPUT68), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT30), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT11), .A3(G134), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G137), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n205), .A2(G134), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT11), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI211_X1 g028(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n205), .C2(G134), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n209), .B(new_n210), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n213), .B1(new_n207), .B2(G137), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n212), .A2(new_n211), .A3(new_n213), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n222), .A2(KEYINPUT66), .A3(new_n210), .A4(new_n209), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n210), .B1(new_n212), .B2(new_n208), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  INV_X1    g042(.A(G146), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G143), .ZN(new_n230));
  INV_X1    g044(.A(G143), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G146), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n228), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n227), .A2(new_n229), .A3(G143), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n234), .B1(new_n228), .B2(new_n232), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n226), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT69), .B1(new_n224), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n239));
  AOI211_X1 g053(.A(new_n239), .B(new_n236), .C1(new_n218), .C2(new_n223), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n206), .A2(new_n208), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n243), .B1(new_n220), .B2(new_n221), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n242), .B1(new_n244), .B2(new_n210), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n209), .B1(new_n214), .B2(new_n215), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(KEYINPUT67), .A3(G131), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n224), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n230), .A2(new_n232), .ZN(new_n250));
  XOR2_X1   g064(.A(KEYINPUT0), .B(G128), .Z(new_n251));
  OR2_X1    g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT0), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n250), .B1(new_n253), .B2(new_n227), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n204), .B1(new_n241), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n236), .B1(new_n218), .B2(new_n223), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n254), .B(KEYINPUT64), .C1(new_n250), .C2(new_n251), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(new_n248), .B2(new_n224), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT64), .B1(new_n252), .B2(new_n254), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  AOI211_X1 g077(.A(KEYINPUT30), .B(new_n258), .C1(new_n261), .C2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n203), .B1(new_n257), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT31), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n203), .B(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n241), .A2(new_n268), .A3(new_n256), .ZN(new_n269));
  INV_X1    g083(.A(G237), .ZN(new_n270));
  INV_X1    g084(.A(G953), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(G210), .ZN(new_n272));
  INV_X1    g086(.A(G101), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n275));
  XOR2_X1   g089(.A(new_n274), .B(new_n275), .Z(new_n276));
  NAND4_X1  g090(.A1(new_n265), .A2(new_n266), .A3(new_n269), .A4(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n276), .ZN(new_n278));
  XOR2_X1   g092(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n245), .A2(new_n247), .B1(new_n218), .B2(new_n223), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n281), .A2(new_n262), .A3(new_n260), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n203), .B1(new_n282), .B2(new_n258), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n280), .B1(new_n283), .B2(new_n269), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n203), .A2(new_n267), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT70), .B1(new_n199), .B2(new_n202), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n224), .A2(new_n237), .ZN(new_n288));
  INV_X1    g102(.A(new_n255), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n288), .B1(new_n281), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n287), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n256), .A2(KEYINPUT72), .A3(new_n288), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT28), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n278), .B1(new_n284), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n277), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n289), .B1(new_n248), .B2(new_n224), .ZN(new_n297));
  NOR4_X1   g111(.A1(new_n287), .A2(new_n297), .A3(new_n238), .A4(new_n240), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n249), .A2(new_n263), .A3(new_n259), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(new_n204), .A3(new_n288), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n297), .A2(new_n238), .A3(new_n240), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n300), .B1(new_n301), .B2(new_n204), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n298), .B1(new_n302), .B2(new_n203), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n266), .B1(new_n303), .B2(new_n276), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n187), .B1(new_n296), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT32), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n203), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n288), .A2(new_n239), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n258), .A2(KEYINPUT69), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n256), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT30), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n308), .B1(new_n312), .B2(new_n300), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n278), .B1(new_n313), .B2(new_n298), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n308), .B1(new_n299), .B2(new_n288), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n279), .B1(new_n298), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n290), .A2(new_n291), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(new_n293), .A3(new_n268), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT28), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n316), .A2(new_n320), .A3(new_n276), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n314), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n278), .A2(new_n322), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n268), .B1(new_n241), .B2(new_n256), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n298), .A2(new_n325), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n320), .B(new_n324), .C1(new_n326), .C2(new_n319), .ZN(new_n327));
  INV_X1    g141(.A(G902), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(G472), .B1(new_n323), .B2(new_n329), .ZN(new_n330));
  OAI211_X1 g144(.A(KEYINPUT32), .B(new_n187), .C1(new_n296), .C2(new_n304), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n307), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G140), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT16), .B1(new_n333), .B2(G125), .ZN(new_n334));
  INV_X1    g148(.A(G125), .ZN(new_n335));
  OAI21_X1  g149(.A(G140), .B1(new_n335), .B2(KEYINPUT74), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT74), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(new_n333), .A3(G125), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n334), .B1(new_n339), .B2(KEYINPUT16), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n340), .A2(new_n229), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n229), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT23), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n192), .B2(G128), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n192), .A2(G128), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n227), .A2(KEYINPUT23), .A3(G119), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G110), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n227), .A2(G119), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n346), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT24), .B(G110), .ZN(new_n352));
  OR2_X1    g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n343), .A2(new_n349), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT75), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n354), .B(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G110), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n345), .A2(new_n347), .A3(new_n357), .A4(new_n346), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n358), .A2(KEYINPUT76), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n351), .A2(new_n352), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n358), .A2(KEYINPUT76), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n359), .A2(new_n360), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n363), .A2(new_n341), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n333), .A2(G125), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n335), .A2(G140), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n366), .A3(new_n229), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(KEYINPUT77), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n364), .A2(KEYINPUT78), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT78), .B1(new_n364), .B2(new_n370), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n356), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT22), .B(G137), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n271), .A2(G221), .A3(G234), .ZN(new_n375));
  XOR2_X1   g189(.A(new_n374), .B(new_n375), .Z(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n356), .B(new_n376), .C1(new_n371), .C2(new_n372), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n328), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT25), .ZN(new_n381));
  INV_X1    g195(.A(G217), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(G234), .B2(new_n328), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n384), .A2(KEYINPUT73), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT25), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n378), .A2(new_n386), .A3(new_n328), .A4(new_n379), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(KEYINPUT73), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n381), .A2(new_n385), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n380), .A2(new_n383), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n332), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n339), .A2(G146), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n270), .A2(new_n271), .A3(G214), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n231), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n270), .A2(new_n271), .A3(G143), .A4(G214), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT88), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT18), .ZN(new_n400));
  OAI22_X1  g214(.A1(new_n398), .A2(new_n399), .B1(new_n400), .B2(new_n210), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n400), .A2(new_n210), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n396), .A2(KEYINPUT88), .A3(new_n397), .A4(new_n402), .ZN(new_n403));
  AOI221_X4 g217(.A(KEYINPUT89), .B1(new_n394), .B2(new_n367), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT89), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n401), .A2(new_n403), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n394), .A2(new_n367), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT90), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n396), .A2(new_n210), .A3(new_n397), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n210), .B1(new_n396), .B2(new_n397), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n412), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(KEYINPUT90), .A3(new_n410), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n415), .A3(new_n341), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n333), .B1(new_n337), .B2(G125), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n335), .A2(KEYINPUT74), .A3(G140), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT19), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT19), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n365), .A2(new_n366), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n229), .A3(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(KEYINPUT91), .ZN(new_n423));
  OAI22_X1  g237(.A1(new_n404), .A2(new_n408), .B1(new_n416), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G113), .B(G122), .ZN(new_n425));
  INV_X1    g239(.A(G104), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n425), .B(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT17), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n414), .A2(new_n430), .A3(new_n410), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n412), .A2(KEYINPUT17), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n431), .A2(new_n341), .A3(new_n342), .A4(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n427), .B(new_n433), .C1(new_n404), .C2(new_n408), .ZN(new_n434));
  AOI21_X1  g248(.A(G475), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT20), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n436), .A3(new_n328), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n436), .B1(new_n435), .B2(new_n328), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n437), .B1(new_n438), .B2(KEYINPUT92), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT92), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n435), .A2(new_n440), .A3(new_n436), .A4(new_n328), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n443), .B1(G128), .B2(new_n231), .ZN(new_n444));
  XNOR2_X1  g258(.A(G128), .B(G143), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(new_n207), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n443), .B2(new_n207), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n194), .A2(G122), .ZN(new_n449));
  INV_X1    g263(.A(G122), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G116), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G107), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n452), .A2(new_n453), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n447), .B(new_n448), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT94), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n449), .B2(KEYINPUT14), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n449), .A2(KEYINPUT14), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT14), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n460), .A2(new_n194), .A3(KEYINPUT94), .A4(G122), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n458), .A2(new_n459), .A3(new_n461), .A4(new_n451), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G107), .ZN(new_n463));
  INV_X1    g277(.A(new_n454), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n445), .B(new_n207), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT95), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n454), .B1(new_n462), .B2(G107), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT95), .B1(new_n469), .B2(new_n465), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n456), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  XOR2_X1   g285(.A(KEYINPUT9), .B(G234), .Z(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n473), .A2(new_n382), .A3(G953), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n456), .B(new_n474), .C1(new_n468), .C2(new_n470), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(KEYINPUT96), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT96), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n471), .A2(new_n479), .A3(new_n475), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(new_n328), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G478), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(KEYINPUT15), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n481), .B(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n408), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n406), .A2(new_n405), .A3(new_n407), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n427), .B1(new_n488), .B2(new_n433), .ZN(new_n489));
  INV_X1    g303(.A(new_n434), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n328), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G475), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n442), .A2(new_n485), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(G234), .A2(G237), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(G952), .A3(new_n271), .ZN(new_n495));
  XOR2_X1   g309(.A(new_n495), .B(KEYINPUT97), .Z(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  XOR2_X1   g311(.A(KEYINPUT21), .B(G898), .Z(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n494), .A2(G902), .A3(G953), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n502), .B(KEYINPUT98), .Z(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n493), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(G214), .B1(G237), .B2(G902), .ZN(new_n506));
  XOR2_X1   g320(.A(new_n506), .B(KEYINPUT82), .Z(new_n507));
  NOR2_X1   g321(.A1(new_n233), .A2(new_n235), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n335), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n289), .B2(new_n335), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n271), .A2(G224), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT3), .B1(new_n426), .B2(G107), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT3), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(new_n453), .A3(G104), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n426), .A2(G107), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G101), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n514), .A2(new_n516), .A3(new_n273), .A4(new_n517), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(KEYINPUT4), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT80), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n519), .A2(KEYINPUT4), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n519), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n520), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n203), .A2(new_n523), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT5), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(new_n192), .A3(G116), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT83), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n529), .B(G113), .C1(new_n527), .C2(new_n196), .ZN(new_n530));
  INV_X1    g344(.A(new_n517), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n426), .A2(G107), .ZN(new_n532));
  OAI21_X1  g346(.A(G101), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n520), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n530), .A2(new_n200), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n526), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G110), .B(G122), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n526), .A2(new_n538), .A3(new_n536), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(KEYINPUT6), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT84), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT6), .ZN(new_n544));
  AND4_X1   g358(.A1(new_n543), .A2(new_n537), .A3(new_n544), .A4(new_n539), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n538), .B1(new_n526), .B2(new_n536), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n543), .B1(new_n546), .B2(new_n544), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n513), .B(new_n542), .C1(new_n545), .C2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(G210), .B1(G237), .B2(G902), .ZN(new_n549));
  XOR2_X1   g363(.A(new_n549), .B(KEYINPUT87), .Z(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n512), .A2(KEYINPUT7), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n511), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(new_n538), .B(KEYINPUT8), .Z(new_n554));
  NAND2_X1  g368(.A1(new_n530), .A2(new_n200), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(KEYINPUT85), .B2(new_n534), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n534), .A2(KEYINPUT85), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n530), .A2(new_n557), .A3(new_n200), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n554), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(KEYINPUT86), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT86), .ZN(new_n561));
  AOI211_X1 g375(.A(new_n561), .B(new_n554), .C1(new_n556), .C2(new_n558), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n541), .B(new_n553), .C1(new_n560), .C2(new_n562), .ZN(new_n563));
  AND4_X1   g377(.A1(new_n328), .A2(new_n548), .A3(new_n551), .A4(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n548), .A2(new_n328), .A3(new_n563), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n550), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n507), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G221), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n472), .B2(new_n328), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n508), .A2(new_n534), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT81), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n235), .B(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(new_n233), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n571), .B1(new_n574), .B2(new_n534), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n575), .A2(KEYINPUT12), .A3(new_n249), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT12), .B1(new_n575), .B2(new_n249), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT10), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n574), .B2(new_n534), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n523), .A2(new_n255), .A3(new_n524), .A4(new_n525), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n509), .A2(new_n535), .A3(KEYINPUT10), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n580), .A2(new_n281), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n271), .A2(G227), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(G140), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT79), .B(G110), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n578), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n249), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n588), .B1(new_n592), .B2(new_n583), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(G469), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n328), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(new_n328), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n583), .B1(new_n576), .B2(new_n577), .ZN(new_n598));
  INV_X1    g412(.A(new_n589), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n598), .A2(new_n587), .B1(new_n599), .B2(new_n592), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n597), .B1(new_n600), .B2(G469), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n570), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n505), .A2(new_n568), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n393), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n567), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n565), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n566), .A2(KEYINPUT100), .A3(new_n550), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n507), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n442), .A2(new_n492), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n481), .A2(new_n482), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n478), .A2(new_n614), .A3(new_n480), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n476), .A2(KEYINPUT33), .A3(new_n477), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n328), .A2(G478), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n613), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n612), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n611), .A2(new_n621), .A3(new_n622), .A4(new_n503), .ZN(new_n623));
  INV_X1    g437(.A(new_n507), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n564), .B1(new_n606), .B2(new_n567), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n503), .B(new_n624), .C1(new_n625), .C2(new_n609), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n612), .A2(new_n620), .ZN(new_n627));
  OAI21_X1  g441(.A(KEYINPUT101), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n265), .A2(new_n269), .A3(new_n276), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT31), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n631), .A2(new_n277), .A3(new_n295), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n328), .ZN(new_n633));
  NAND2_X1  g447(.A1(KEYINPUT99), .A2(G472), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n389), .A2(new_n390), .ZN(new_n636));
  INV_X1    g450(.A(new_n602), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n629), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  INV_X1    g457(.A(new_n485), .ZN(new_n644));
  INV_X1    g458(.A(new_n438), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n645), .A2(new_n437), .B1(G475), .B2(new_n491), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n611), .A2(new_n503), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n639), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT35), .B(G107), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  NOR2_X1   g465(.A1(new_n377), .A2(KEYINPUT36), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n373), .B(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n328), .A3(new_n384), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n389), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n603), .A2(new_n635), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT37), .B(G110), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G12));
  AND3_X1   g472(.A1(new_n332), .A2(new_n602), .A3(new_n655), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n496), .B(KEYINPUT102), .Z(new_n660));
  INV_X1    g474(.A(G900), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n660), .B1(new_n661), .B2(new_n501), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n659), .A2(new_n611), .A3(new_n647), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G128), .ZN(G30));
  NAND2_X1  g479(.A1(new_n565), .A2(new_n567), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n666), .B(KEYINPUT38), .Z(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT104), .B(KEYINPUT39), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n662), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n602), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(KEYINPUT40), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n442), .A2(new_n492), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n672), .A2(new_n485), .A3(new_n673), .ZN(new_n674));
  AOI211_X1 g488(.A(new_n507), .B(new_n655), .C1(new_n671), .C2(KEYINPUT40), .ZN(new_n675));
  INV_X1    g489(.A(new_n331), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT32), .B1(new_n632), .B2(new_n187), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n630), .B(G472), .C1(new_n276), .C2(new_n326), .ZN(new_n679));
  NAND2_X1  g493(.A1(G472), .A2(G902), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n679), .A2(KEYINPUT103), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(KEYINPUT103), .B1(new_n679), .B2(new_n680), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n668), .A2(new_n674), .A3(new_n675), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G143), .ZN(G45));
  AND2_X1   g500(.A1(new_n389), .A2(new_n654), .ZN(new_n687));
  INV_X1    g501(.A(G472), .ZN(new_n688));
  INV_X1    g502(.A(new_n329), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n314), .A2(new_n321), .A3(new_n322), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n676), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n687), .B1(new_n692), .B2(new_n307), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n612), .A2(new_n620), .A3(new_n663), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n693), .A2(new_n602), .A3(new_n611), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  OAI21_X1  g511(.A(new_n328), .B1(new_n590), .B2(new_n593), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n595), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n570), .ZN(new_n702));
  OAI221_X1 g516(.A(new_n328), .B1(new_n699), .B2(new_n595), .C1(new_n590), .C2(new_n593), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n332), .A2(new_n391), .A3(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n629), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NOR2_X1   g523(.A1(new_n705), .A2(new_n648), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n194), .ZN(G18));
  NAND3_X1  g525(.A1(new_n332), .A2(new_n505), .A3(new_n655), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n608), .A2(new_n610), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(new_n714), .A3(new_n624), .A4(new_n704), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n624), .B(new_n704), .C1(new_n625), .C2(new_n609), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT106), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n712), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n192), .ZN(G21));
  NAND2_X1  g533(.A1(new_n311), .A2(new_n287), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n319), .B1(new_n720), .B2(new_n269), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n278), .B1(new_n721), .B2(new_n294), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n631), .A2(KEYINPUT107), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n277), .ZN(new_n724));
  AOI21_X1  g538(.A(KEYINPUT107), .B1(new_n631), .B2(new_n722), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n187), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n633), .A2(G472), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n391), .A3(new_n704), .A4(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n485), .B1(new_n442), .B2(new_n492), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n713), .A2(new_n503), .A3(new_n624), .A4(new_n729), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  AND3_X1   g546(.A1(new_n726), .A2(new_n655), .A3(new_n727), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n714), .B1(new_n611), .B2(new_n704), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n716), .A2(KEYINPUT106), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n733), .B(new_n695), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  OR2_X1    g551(.A1(new_n307), .A2(KEYINPUT108), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n307), .A2(KEYINPUT108), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n692), .A3(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT42), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n565), .A2(new_n624), .A3(new_n567), .ZN(new_n742));
  NOR4_X1   g556(.A1(new_n694), .A2(new_n637), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n740), .A2(new_n743), .A3(new_n391), .ZN(new_n744));
  INV_X1    g558(.A(new_n742), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n695), .A2(new_n602), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n741), .B1(new_n746), .B2(new_n392), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT109), .B(G131), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G33));
  NOR2_X1   g564(.A1(new_n742), .A2(new_n662), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n638), .A2(new_n332), .A3(new_n647), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G134), .ZN(G36));
  NAND2_X1  g567(.A1(new_n673), .A2(new_n620), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT43), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  AOI211_X1 g572(.A(new_n635), .B(new_n687), .C1(new_n756), .C2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n742), .B1(new_n759), .B2(KEYINPUT44), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n600), .A2(KEYINPUT45), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n600), .A2(KEYINPUT110), .A3(KEYINPUT45), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n595), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n600), .A2(KEYINPUT45), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n597), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n767), .A2(KEYINPUT46), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n596), .B1(new_n767), .B2(KEYINPUT46), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n702), .A3(new_n670), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n760), .B(new_n772), .C1(KEYINPUT44), .C2(new_n759), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G137), .ZN(G39));
  OAI21_X1  g588(.A(new_n702), .B1(new_n768), .B2(new_n769), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT47), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n391), .A2(new_n694), .A3(new_n742), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n777), .A2(new_n307), .A3(new_n692), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  INV_X1    g594(.A(new_n660), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n781), .B1(new_n756), .B2(new_n758), .ZN(new_n782));
  INV_X1    g596(.A(new_n704), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n742), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n733), .ZN(new_n786));
  INV_X1    g600(.A(new_n684), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n783), .A2(new_n636), .A3(new_n742), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n497), .A3(new_n673), .A4(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n790));
  OR3_X1    g604(.A1(new_n789), .A2(new_n790), .A3(new_n620), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n790), .B1(new_n789), .B2(new_n620), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n786), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n726), .A2(new_n727), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n782), .A2(new_n391), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n704), .A2(new_n507), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT115), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n796), .A2(KEYINPUT50), .A3(new_n667), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n782), .A2(new_n391), .A3(new_n667), .A4(new_n795), .ZN(new_n801));
  INV_X1    g615(.A(new_n798), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n793), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT118), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n701), .A2(new_n703), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n702), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n745), .B(new_n796), .C1(new_n777), .C2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT118), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n793), .A2(new_n804), .A3(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n806), .A2(KEYINPUT51), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n799), .A2(new_n803), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n814), .B1(new_n799), .B2(new_n803), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n810), .B(new_n793), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n740), .A2(new_n391), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n785), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT48), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n796), .B1(new_n735), .B2(new_n734), .ZN(new_n823));
  AND4_X1   g637(.A1(G952), .A2(new_n822), .A3(new_n271), .A4(new_n823), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n813), .A2(new_n819), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n332), .A2(new_n485), .A3(new_n646), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n627), .B2(new_n794), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n602), .A3(new_n655), .A4(new_n751), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n748), .A2(new_n828), .A3(new_n752), .ZN(new_n829));
  MUX2_X1   g643(.A(new_n644), .B(new_n620), .S(new_n612), .Z(new_n830));
  NAND4_X1  g644(.A1(new_n640), .A2(new_n503), .A3(new_n568), .A4(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n604), .A3(new_n656), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n710), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n693), .B(new_n505), .C1(new_n734), .C2(new_n735), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n707), .A2(new_n834), .A3(new_n835), .A4(new_n731), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(KEYINPUT112), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT112), .ZN(new_n838));
  OAI22_X1  g652(.A1(new_n705), .A2(new_n648), .B1(new_n728), .B2(new_n730), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n718), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n838), .B1(new_n840), .B2(new_n707), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n829), .B(new_n833), .C1(new_n837), .C2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT113), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n637), .B1(new_n678), .B2(new_n683), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n729), .B(new_n624), .C1(new_n625), .C2(new_n609), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n844), .A2(new_n687), .A3(new_n663), .A4(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n664), .A2(new_n736), .A3(new_n847), .A4(new_n696), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n694), .B1(new_n715), .B2(new_n717), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n332), .A2(new_n611), .A3(new_n602), .A4(new_n655), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n851), .A2(new_n733), .B1(new_n852), .B2(new_n695), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(KEYINPUT52), .A3(new_n664), .A4(new_n847), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT114), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n850), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n836), .A2(KEYINPUT112), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n840), .A2(new_n838), .A3(new_n707), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n832), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT113), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(new_n863), .A3(new_n829), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n843), .A2(new_n859), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT53), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n843), .A2(new_n864), .A3(new_n867), .A4(new_n855), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(KEYINPUT54), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n865), .A2(new_n867), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n832), .A2(new_n867), .ZN(new_n872));
  INV_X1    g686(.A(new_n836), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n855), .A2(new_n872), .A3(new_n829), .A4(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n825), .A2(new_n869), .A3(new_n875), .ZN(new_n876));
  AND4_X1   g690(.A1(new_n497), .A2(new_n787), .A3(new_n621), .A4(new_n788), .ZN(new_n877));
  OAI22_X1  g691(.A1(new_n876), .A2(new_n877), .B1(G952), .B2(G953), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n391), .A2(new_n624), .A3(new_n702), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(KEYINPUT111), .ZN(new_n880));
  AOI211_X1 g694(.A(new_n668), .B(new_n880), .C1(KEYINPUT49), .C2(new_n808), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n755), .B1(KEYINPUT49), .B2(new_n808), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(KEYINPUT111), .B2(new_n879), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n881), .A2(new_n787), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n878), .A2(new_n884), .ZN(G75));
  OAI21_X1  g699(.A(new_n542), .B1(new_n545), .B2(new_n547), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n513), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT55), .Z(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n888), .B1(KEYINPUT119), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n874), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n865), .B2(new_n867), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n893), .A2(new_n328), .A3(new_n551), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n891), .B1(new_n894), .B2(KEYINPUT56), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n870), .A2(new_n874), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(G902), .A3(new_n550), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n889), .A3(new_n890), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n271), .A2(G952), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n895), .A2(new_n898), .A3(new_n900), .ZN(G51));
  XNOR2_X1  g715(.A(new_n597), .B(KEYINPUT120), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT57), .Z(new_n903));
  AOI21_X1  g717(.A(new_n871), .B1(new_n870), .B2(new_n874), .ZN(new_n904));
  AOI211_X1 g718(.A(KEYINPUT54), .B(new_n892), .C1(new_n865), .C2(new_n867), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n594), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n893), .A2(new_n328), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n766), .A3(new_n765), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n899), .B1(new_n907), .B2(new_n909), .ZN(G54));
  NAND4_X1  g724(.A1(new_n896), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n911), .A2(new_n434), .A3(new_n429), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n429), .A2(new_n434), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n908), .A2(KEYINPUT58), .A3(G475), .A4(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n912), .A2(new_n900), .A3(new_n914), .ZN(G60));
  NAND2_X1  g729(.A1(G478), .A2(G902), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT59), .Z(new_n917));
  NOR2_X1   g731(.A1(new_n618), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n904), .B2(new_n905), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n917), .B1(new_n869), .B2(new_n875), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n919), .B(new_n900), .C1(new_n920), .C2(new_n617), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(G63));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n896), .A2(new_n653), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n378), .A2(new_n379), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n893), .B2(new_n924), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n926), .A2(new_n900), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT61), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n926), .A2(new_n928), .A3(KEYINPUT61), .A4(new_n900), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(G66));
  INV_X1    g747(.A(G224), .ZN(new_n934));
  OAI21_X1  g748(.A(G953), .B1(new_n499), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n862), .B2(G953), .ZN(new_n936));
  MUX2_X1   g750(.A(new_n935), .B(new_n936), .S(KEYINPUT121), .Z(new_n937));
  OAI21_X1  g751(.A(new_n886), .B1(G898), .B2(new_n271), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G69));
  NAND2_X1  g753(.A1(new_n419), .A2(new_n421), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n302), .B(new_n940), .Z(new_n941));
  NAND2_X1  g755(.A1(G900), .A2(G953), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n773), .A2(new_n779), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n748), .A2(new_n752), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n664), .A2(new_n736), .A3(new_n696), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n945), .A2(KEYINPUT122), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(KEYINPUT122), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n772), .A2(new_n846), .A3(new_n820), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n943), .A2(new_n944), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n941), .B(new_n942), .C1(new_n950), .C2(G953), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT123), .ZN(new_n953));
  AOI211_X1 g767(.A(new_n742), .B(new_n392), .C1(new_n830), .C2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n671), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n954), .B(new_n955), .C1(new_n953), .C2(new_n830), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n946), .A2(new_n685), .A3(new_n947), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT62), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n943), .B(new_n956), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n941), .B1(new_n961), .B2(new_n271), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n952), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(G227), .ZN(new_n964));
  OAI21_X1  g778(.A(G953), .B1(new_n964), .B2(new_n661), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n963), .B(new_n965), .ZN(G72));
  XNOR2_X1  g780(.A(new_n680), .B(KEYINPUT63), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n862), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n968), .B1(new_n961), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n303), .B(KEYINPUT124), .Z(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(new_n278), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n314), .B(KEYINPUT126), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n967), .B1(new_n974), .B2(new_n630), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n866), .A2(new_n868), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n968), .B1(new_n950), .B2(new_n969), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n971), .A2(new_n278), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT125), .Z(new_n979));
  AOI21_X1  g793(.A(new_n899), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n973), .A2(new_n976), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(KEYINPUT127), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n973), .A2(new_n980), .A3(new_n983), .A4(new_n976), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(G57));
endmodule


