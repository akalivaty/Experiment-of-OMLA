//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974;
  INV_X1    g000(.A(KEYINPUT99), .ZN(new_n202));
  NOR2_X1   g001(.A1(G71gat), .A2(G78gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT9), .ZN(new_n204));
  INV_X1    g003(.A(G71gat), .ZN(new_n205));
  INV_X1    g004(.A(G78gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G57gat), .ZN(new_n208));
  AND2_X1   g007(.A1(new_n208), .A2(G64gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n209), .B(KEYINPUT94), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n208), .A2(G64gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(new_n203), .B(KEYINPUT93), .Z(new_n213));
  OAI21_X1  g012(.A(KEYINPUT9), .B1(new_n209), .B2(new_n211), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n213), .B(new_n214), .C1(new_n205), .C2(new_n206), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT21), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n219));
  XOR2_X1   g018(.A(new_n218), .B(new_n219), .Z(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G15gat), .B(G22gat), .ZN(new_n222));
  INV_X1    g021(.A(G1gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT16), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G1gat), .B2(new_n222), .ZN(new_n226));
  INV_X1    g025(.A(G8gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(new_n216), .B2(new_n217), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(G183gat), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n230), .A2(KEYINPUT95), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(KEYINPUT95), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n233), .A2(G231gat), .A3(G233gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(G231gat), .A2(G233gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(new_n231), .B2(new_n232), .ZN(new_n236));
  XNOR2_X1  g035(.A(G127gat), .B(G155gat), .ZN(new_n237));
  INV_X1    g036(.A(G211gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n234), .A2(new_n236), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n240), .B1(new_n234), .B2(new_n236), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n221), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n243), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(new_n220), .A3(new_n241), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G85gat), .A2(G92gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT7), .ZN(new_n250));
  NAND2_X1  g049(.A1(G99gat), .A2(G106gat), .ZN(new_n251));
  INV_X1    g050(.A(G85gat), .ZN(new_n252));
  INV_X1    g051(.A(G92gat), .ZN(new_n253));
  AOI22_X1  g052(.A1(KEYINPUT8), .A2(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G99gat), .B(G106gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT96), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT96), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n250), .A2(new_n259), .A3(new_n256), .A4(new_n254), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  OR3_X1    g062(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n263), .B1(new_n264), .B2(KEYINPUT90), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n265), .B1(KEYINPUT90), .B2(new_n264), .ZN(new_n266));
  INV_X1    g065(.A(G29gat), .ZN(new_n267));
  INV_X1    g066(.A(G36gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G43gat), .B(G50gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT15), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(KEYINPUT91), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT17), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n264), .A2(new_n262), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n275), .B1(new_n267), .B2(new_n268), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n276), .A2(KEYINPUT15), .A3(new_n270), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n273), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n274), .B1(new_n273), .B2(new_n277), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n261), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT97), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n273), .A2(new_n277), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n258), .A2(new_n260), .ZN(new_n283));
  AND2_X1   g082(.A1(G232gat), .A2(G233gat), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n282), .A2(new_n283), .B1(KEYINPUT41), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT97), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n286), .B(new_n261), .C1(new_n278), .C2(new_n279), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n281), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G134gat), .B(G162gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n289), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n281), .A2(new_n291), .A3(new_n285), .A4(new_n287), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  XOR2_X1   g092(.A(G190gat), .B(G218gat), .Z(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT98), .ZN(new_n295));
  OR2_X1    g094(.A1(new_n284), .A2(KEYINPUT41), .ZN(new_n296));
  XOR2_X1   g095(.A(new_n295), .B(new_n296), .Z(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n290), .A2(new_n297), .A3(new_n292), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n202), .B1(new_n248), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n247), .A2(new_n301), .A3(KEYINPUT99), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G230gat), .ZN(new_n306));
  INV_X1    g105(.A(G233gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n283), .A2(new_n216), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n216), .A2(new_n257), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT10), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n283), .A2(KEYINPUT10), .A3(new_n212), .A4(new_n215), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n309), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n310), .A2(new_n311), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n316), .B1(new_n308), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G176gat), .B(G204gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(KEYINPUT100), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(G120gat), .ZN(new_n322));
  INV_X1    g121(.A(G148gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n319), .B(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n305), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT18), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n228), .B1(new_n278), .B2(new_n279), .ZN(new_n329));
  INV_X1    g128(.A(new_n228), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n282), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G229gat), .A2(G233gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n328), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n282), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n228), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT92), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n338), .A3(new_n331), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n333), .B(KEYINPUT13), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n282), .A2(KEYINPUT92), .A3(new_n330), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n329), .A2(KEYINPUT18), .A3(new_n333), .A4(new_n331), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n335), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(G169gat), .B(G197gat), .Z(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(KEYINPUT89), .ZN(new_n347));
  XNOR2_X1  g146(.A(G113gat), .B(G141gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  XOR2_X1   g148(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT12), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n345), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n335), .A2(new_n343), .A3(new_n352), .A4(new_n344), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT85), .ZN(new_n358));
  XOR2_X1   g157(.A(G78gat), .B(G106gat), .Z(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT31), .ZN(new_n360));
  XOR2_X1   g159(.A(new_n360), .B(G50gat), .Z(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n323), .A2(G141gat), .ZN(new_n363));
  INV_X1    g162(.A(G141gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G148gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT74), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G141gat), .B(G148gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT74), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT75), .B(KEYINPUT2), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n368), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G155gat), .ZN(new_n374));
  INV_X1    g173(.A(G162gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT76), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n363), .A2(new_n365), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n380), .B1(new_n363), .B2(new_n365), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n377), .B1(new_n376), .B2(KEYINPUT2), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n373), .A2(new_n379), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(G211gat), .A2(G218gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT22), .ZN(new_n387));
  NAND2_X1  g186(.A1(G211gat), .A2(G218gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G197gat), .B(G204gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT81), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(KEYINPUT22), .ZN(new_n393));
  INV_X1    g192(.A(new_n388), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(new_n386), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n389), .A2(new_n397), .A3(new_n390), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n392), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n385), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n393), .A2(new_n395), .B1(new_n389), .B2(new_n390), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n373), .A2(new_n379), .ZN(new_n406));
  INV_X1    g205(.A(new_n382), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n369), .A2(new_n380), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(new_n408), .A3(new_n384), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n406), .A2(new_n402), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n405), .B1(new_n410), .B2(new_n400), .ZN(new_n411));
  INV_X1    g210(.A(G228gat), .ZN(new_n412));
  OAI22_X1  g211(.A1(new_n403), .A2(new_n411), .B1(new_n412), .B2(new_n307), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n307), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT3), .B1(new_n405), .B2(new_n400), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT29), .B1(new_n385), .B2(new_n402), .ZN(new_n416));
  OAI221_X1 g215(.A(new_n414), .B1(new_n415), .B2(new_n385), .C1(new_n416), .C2(new_n405), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n362), .B1(new_n418), .B2(G22gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT82), .B(G22gat), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n413), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT84), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT84), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n413), .A2(new_n417), .A3(new_n424), .A4(new_n421), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n419), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT83), .ZN(new_n427));
  INV_X1    g226(.A(new_n422), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n421), .B1(new_n413), .B2(new_n417), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n362), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g230(.A(KEYINPUT83), .B(new_n362), .C1(new_n428), .C2(new_n429), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AND2_X1   g232(.A1(KEYINPUT67), .A2(G113gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(KEYINPUT67), .A2(G113gat), .ZN(new_n435));
  OAI21_X1  g234(.A(G120gat), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(G120gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G113gat), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT1), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G127gat), .B(G134gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(G127gat), .A2(G134gat), .ZN(new_n442));
  AND2_X1   g241(.A1(KEYINPUT66), .A2(G127gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(KEYINPUT66), .A2(G127gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n442), .B1(new_n445), .B2(G134gat), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT1), .ZN(new_n447));
  INV_X1    g246(.A(new_n438), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n437), .A2(G113gat), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n441), .A2(new_n451), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n363), .A2(new_n365), .A3(KEYINPUT74), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT74), .B1(new_n363), .B2(new_n365), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n453), .A2(new_n454), .A3(new_n371), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n409), .B1(new_n455), .B2(new_n378), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT77), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT3), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT77), .B1(new_n385), .B2(new_n402), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n385), .A2(new_n402), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n452), .B(new_n458), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n439), .A2(new_n440), .B1(new_n446), .B2(new_n450), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT4), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n462), .A2(new_n406), .A3(new_n463), .A4(new_n409), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT80), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT4), .B1(new_n456), .B2(new_n452), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT80), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n385), .A2(new_n467), .A3(new_n463), .A4(new_n462), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(G225gat), .A2(G233gat), .ZN(new_n470));
  XOR2_X1   g269(.A(new_n470), .B(KEYINPUT78), .Z(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(KEYINPUT5), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n461), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n471), .B1(new_n466), .B2(new_n464), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n461), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT79), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT5), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n456), .B(new_n452), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n477), .B1(new_n478), .B2(new_n471), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n475), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n476), .B1(new_n475), .B2(new_n479), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n473), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT0), .B(G57gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(G85gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(G1gat), .B(G29gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n484), .B(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT6), .ZN(new_n488));
  INV_X1    g287(.A(new_n486), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n489), .B(new_n473), .C1(new_n480), .C2(new_n481), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n482), .A2(KEYINPUT6), .A3(new_n486), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(G64gat), .B(G92gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(KEYINPUT73), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(G8gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(new_n268), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT71), .ZN(new_n498));
  AND2_X1   g297(.A1(G226gat), .A2(G233gat), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(G183gat), .A2(G190gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g303(.A1(G169gat), .A2(G176gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT23), .ZN(new_n506));
  INV_X1    g305(.A(G169gat), .ZN(new_n507));
  INV_X1    g306(.A(G176gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT25), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n503), .A2(KEYINPUT64), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT64), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n516), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n502), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n518), .A2(new_n511), .A3(KEYINPUT25), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT26), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT26), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(G169gat), .B2(G176gat), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n521), .B(new_n501), .C1(new_n523), .C2(new_n505), .ZN(new_n524));
  INV_X1    g323(.A(G190gat), .ZN(new_n525));
  AND2_X1   g324(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT28), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g329(.A(KEYINPUT28), .B(new_n525), .C1(new_n526), .C2(new_n527), .ZN(new_n531));
  AOI211_X1 g330(.A(KEYINPUT65), .B(new_n524), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT65), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n530), .A2(new_n531), .ZN(new_n534));
  INV_X1    g333(.A(new_n524), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n499), .B(new_n520), .C1(new_n532), .C2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT27), .B(G183gat), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT28), .B1(new_n538), .B2(new_n525), .ZN(new_n539));
  INV_X1    g338(.A(new_n531), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n535), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n519), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT25), .B1(new_n504), .B2(new_n511), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n499), .A2(KEYINPUT29), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n537), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n498), .B1(new_n547), .B2(new_n405), .ZN(new_n548));
  AOI211_X1 g347(.A(KEYINPUT71), .B(new_n404), .C1(new_n537), .C2(new_n546), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n520), .A2(new_n499), .A3(new_n541), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n541), .A2(KEYINPUT65), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n534), .A2(new_n533), .A3(new_n535), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n552), .A2(new_n553), .B1(new_n514), .B2(new_n519), .ZN(new_n554));
  INV_X1    g353(.A(new_n545), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n404), .B(new_n551), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT70), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n520), .B1(new_n532), .B2(new_n536), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(new_n545), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT70), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n559), .A2(new_n560), .A3(new_n404), .A4(new_n551), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n550), .A2(new_n562), .A3(KEYINPUT72), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT72), .B1(new_n550), .B2(new_n562), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n497), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT30), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n562), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n566), .B1(new_n567), .B2(new_n497), .ZN(new_n568));
  INV_X1    g367(.A(new_n567), .ZN(new_n569));
  INV_X1    g368(.A(new_n497), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(KEYINPUT30), .A3(new_n570), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n565), .A2(new_n568), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n433), .B1(new_n493), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT34), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT68), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n574), .A2(KEYINPUT68), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n558), .A2(new_n452), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n462), .B(new_n520), .C1(new_n532), .C2(new_n536), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(G227gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n581), .A2(new_n307), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n575), .B(new_n577), .C1(new_n580), .C2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n582), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n578), .A2(new_n584), .A3(new_n579), .A4(new_n576), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G15gat), .B(G43gat), .Z(new_n587));
  XNOR2_X1  g386(.A(G71gat), .B(G99gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n584), .B1(new_n578), .B2(new_n579), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n589), .B1(new_n590), .B2(KEYINPUT33), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT32), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  AOI221_X4 g393(.A(new_n592), .B1(KEYINPUT33), .B2(new_n589), .C1(new_n580), .C2(new_n582), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n586), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT69), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n552), .A2(new_n553), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n462), .B1(new_n598), .B2(new_n520), .ZN(new_n599));
  INV_X1    g398(.A(new_n579), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n582), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT32), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n602), .A2(new_n604), .A3(new_n589), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n591), .A2(new_n593), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n583), .A2(new_n585), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n596), .A2(new_n597), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n605), .A2(new_n606), .A3(new_n607), .A4(KEYINPUT69), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n596), .A2(KEYINPUT36), .A3(new_n608), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n358), .B1(new_n573), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n565), .A2(new_n568), .A3(new_n571), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n478), .A2(new_n471), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT87), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n461), .A2(new_n469), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n471), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(KEYINPUT39), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n619), .A2(new_n622), .A3(new_n471), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n623), .A2(KEYINPUT86), .A3(new_n489), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT86), .B1(new_n623), .B2(new_n489), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT40), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n621), .B(KEYINPUT40), .C1(new_n624), .C2(new_n625), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n616), .A2(new_n628), .A3(new_n487), .A4(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n567), .A2(KEYINPUT37), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT38), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n547), .A2(new_n404), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n559), .A2(new_n405), .A3(new_n551), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n633), .A2(new_n634), .A3(KEYINPUT37), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n631), .A2(new_n632), .A3(new_n497), .A4(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n570), .B1(new_n569), .B2(KEYINPUT38), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n491), .A2(new_n636), .A3(new_n637), .A4(new_n492), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT37), .B1(new_n563), .B2(new_n564), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n632), .B1(new_n639), .B2(new_n631), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n630), .B(new_n433), .C1(new_n638), .C2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n612), .A2(new_n613), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n616), .B1(new_n492), .B2(new_n491), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n642), .B(KEYINPUT85), .C1(new_n643), .C2(new_n433), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n615), .A2(new_n641), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n433), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT35), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n596), .A2(new_n608), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n609), .A2(new_n611), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n493), .A2(new_n572), .A3(new_n433), .A4(new_n650), .ZN(new_n651));
  AOI22_X1  g450(.A1(new_n649), .A2(new_n643), .B1(new_n651), .B2(new_n647), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n357), .B1(new_n645), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n327), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n493), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT101), .B(G1gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(G1324gat));
  NOR2_X1   g456(.A1(new_n654), .A2(new_n572), .ZN(new_n658));
  NAND2_X1  g457(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n659));
  OR2_X1    g458(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n663), .B(new_n664), .C1(new_n227), .C2(new_n658), .ZN(G1325gat));
  INV_X1    g464(.A(G15gat), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n654), .A2(new_n666), .A3(new_n642), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n327), .A2(new_n650), .A3(new_n653), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n667), .B1(new_n666), .B2(new_n668), .ZN(G1326gat));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n433), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT43), .B(G22gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1327gat));
  NAND4_X1  g471(.A1(new_n653), .A2(new_n248), .A3(new_n302), .A4(new_n326), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n673), .A2(G29gat), .A3(new_n493), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(KEYINPUT45), .Z(new_n675));
  AND2_X1   g474(.A1(new_n491), .A2(new_n492), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n645), .A2(new_n652), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n302), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(new_n679), .A3(KEYINPUT44), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT104), .B1(new_n643), .B2(new_n433), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n682), .B(new_n646), .C1(new_n676), .C2(new_n616), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n681), .A2(new_n641), .A3(new_n683), .A4(new_n642), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n301), .B1(new_n684), .B2(new_n652), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n301), .B1(new_n645), .B2(new_n652), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT103), .B1(new_n688), .B2(new_n686), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n680), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n247), .B(KEYINPUT102), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n357), .A2(new_n325), .ZN(new_n692));
  AND4_X1   g491(.A1(new_n676), .A2(new_n690), .A3(new_n691), .A4(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n675), .B1(new_n267), .B2(new_n693), .ZN(G1328gat));
  AOI21_X1  g493(.A(new_n673), .B1(KEYINPUT105), .B2(KEYINPUT46), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n695), .A2(new_n268), .A3(new_n616), .ZN(new_n696));
  NOR2_X1   g495(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(new_n698));
  AND4_X1   g497(.A1(new_n616), .A2(new_n690), .A3(new_n691), .A4(new_n692), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n268), .B2(new_n699), .ZN(G1329gat));
  NAND4_X1  g499(.A1(new_n690), .A2(new_n614), .A3(new_n691), .A4(new_n692), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(G43gat), .ZN(new_n702));
  INV_X1    g501(.A(new_n650), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n673), .A2(G43gat), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT47), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708));
  AOI211_X1 g507(.A(KEYINPUT106), .B(new_n708), .C1(new_n702), .C2(new_n704), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n707), .A2(new_n709), .ZN(G1330gat));
  NAND4_X1  g509(.A1(new_n690), .A2(new_n646), .A3(new_n691), .A4(new_n692), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT107), .B1(new_n711), .B2(G50gat), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n673), .A2(G50gat), .A3(new_n433), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n713), .B1(new_n711), .B2(G50gat), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT48), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI221_X4 g515(.A(new_n713), .B1(KEYINPUT107), .B2(KEYINPUT48), .C1(new_n711), .C2(G50gat), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(G1331gat));
  NAND2_X1  g517(.A1(new_n684), .A2(new_n652), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n305), .A2(new_n357), .A3(new_n325), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT108), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n493), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(new_n208), .ZN(G1332gat));
  NOR2_X1   g522(.A1(new_n721), .A2(new_n572), .ZN(new_n724));
  NOR2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  AND2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n724), .B2(new_n725), .ZN(G1333gat));
  XOR2_X1   g527(.A(new_n720), .B(KEYINPUT108), .Z(new_n729));
  AOI21_X1  g528(.A(G71gat), .B1(new_n729), .B2(new_n650), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n721), .A2(new_n205), .A3(new_n642), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT50), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n729), .A2(G71gat), .A3(new_n614), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n205), .B1(new_n721), .B2(new_n703), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n732), .A2(new_n736), .ZN(G1334gat));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n433), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(new_n206), .ZN(G1335gat));
  NAND4_X1  g538(.A1(new_n244), .A2(new_n246), .A3(new_n354), .A4(new_n355), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n719), .A2(new_n302), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT51), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(KEYINPUT109), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n742), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(KEYINPUT109), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(new_n676), .A3(new_n325), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n740), .A2(new_n326), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n690), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n493), .A2(new_n252), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n748), .A2(new_n252), .B1(new_n750), .B2(new_n751), .ZN(G1336gat));
  NAND3_X1  g551(.A1(new_n690), .A2(new_n616), .A3(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G92gat), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n747), .A2(new_n325), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n572), .A2(G92gat), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n754), .B(new_n755), .C1(new_n756), .C2(new_n758), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n753), .A2(KEYINPUT110), .A3(G92gat), .ZN(new_n760));
  AOI211_X1 g559(.A(KEYINPUT111), .B(new_n743), .C1(new_n685), .C2(new_n741), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT51), .B1(new_n742), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n764), .A2(KEYINPUT112), .A3(new_n325), .A4(new_n757), .ZN(new_n765));
  AOI211_X1 g564(.A(new_n301), .B(new_n740), .C1(new_n684), .C2(new_n652), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n743), .B1(new_n766), .B2(KEYINPUT111), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n742), .A2(new_n762), .A3(KEYINPUT51), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n767), .A2(new_n325), .A3(new_n768), .A4(new_n757), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n765), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT110), .B1(new_n753), .B2(G92gat), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n760), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n759), .B1(new_n774), .B2(new_n755), .ZN(G1337gat));
  NAND2_X1  g574(.A1(new_n750), .A2(new_n614), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G99gat), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n756), .A2(G99gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n703), .ZN(G1338gat));
  NOR3_X1   g578(.A1(new_n326), .A2(G106gat), .A3(new_n433), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n747), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n750), .A2(new_n646), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G106gat), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI22_X1  g586(.A1(new_n784), .A2(G106gat), .B1(new_n764), .B2(new_n780), .ZN(new_n788));
  OAI22_X1  g587(.A1(new_n783), .A2(new_n787), .B1(new_n788), .B2(new_n786), .ZN(G1339gat));
  XNOR2_X1  g588(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n316), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n324), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT10), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n317), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(new_n308), .A3(new_n313), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(KEYINPUT54), .A3(new_n315), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n791), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n319), .A2(new_n324), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n791), .A2(new_n796), .A3(KEYINPUT55), .A4(new_n792), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT115), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT115), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n803), .A2(new_n356), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n332), .A2(new_n334), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n339), .A2(new_n342), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n340), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n332), .A2(KEYINPUT116), .A3(new_n334), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n810), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n351), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(new_n355), .A3(new_n325), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n302), .B1(new_n807), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n803), .A2(new_n806), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n355), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n818), .A2(new_n301), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n691), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n303), .A2(new_n357), .A3(new_n304), .A4(new_n326), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n646), .A2(new_n648), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n493), .A2(new_n616), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n826), .A2(KEYINPUT118), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n434), .A2(new_n435), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(KEYINPUT118), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n827), .A2(new_n828), .A3(new_n356), .A4(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n823), .A2(new_n825), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n650), .A3(new_n433), .ZN(new_n832));
  OAI21_X1  g631(.A(G113gat), .B1(new_n832), .B2(new_n357), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n830), .B1(new_n835), .B2(new_n836), .ZN(G1340gat));
  NAND4_X1  g636(.A1(new_n827), .A2(new_n437), .A3(new_n325), .A4(new_n829), .ZN(new_n838));
  OAI21_X1  g637(.A(G120gat), .B1(new_n832), .B2(new_n326), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(new_n839), .A3(KEYINPUT119), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1341gat));
  NOR2_X1   g643(.A1(new_n826), .A2(new_n248), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n445), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n832), .A2(new_n691), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n445), .ZN(G1342gat));
  OAI21_X1  g647(.A(G134gat), .B1(new_n832), .B2(new_n301), .ZN(new_n849));
  INV_X1    g648(.A(G134gat), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n831), .A2(new_n850), .A3(new_n824), .A4(new_n302), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT56), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n826), .A2(G134gat), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n854), .A3(new_n302), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n849), .A2(new_n852), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT120), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n849), .A2(new_n852), .A3(new_n855), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(G1343gat));
  NAND2_X1  g659(.A1(new_n823), .A2(new_n646), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n816), .A2(KEYINPUT121), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n356), .A2(new_n802), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n815), .A2(new_n866), .A3(new_n355), .A4(new_n325), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n820), .B1(new_n301), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n822), .B1(new_n869), .B2(new_n247), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(KEYINPUT57), .A3(new_n646), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n863), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n825), .A2(new_n642), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n356), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(G141gat), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n823), .A2(new_n646), .A3(new_n874), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n878), .A2(G141gat), .A3(new_n357), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n873), .B1(new_n863), .B2(new_n871), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n364), .B1(new_n882), .B2(new_n356), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT58), .B1(new_n883), .B2(new_n879), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(new_n884), .ZN(G1344gat));
  INV_X1    g684(.A(new_n878), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n323), .A3(new_n325), .ZN(new_n887));
  AOI211_X1 g686(.A(KEYINPUT59), .B(new_n323), .C1(new_n882), .C2(new_n325), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n861), .A2(KEYINPUT57), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n868), .A2(new_n301), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n302), .A2(new_n355), .A3(new_n802), .A4(new_n815), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n247), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n822), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n862), .B(new_n646), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n890), .A2(new_n895), .A3(new_n325), .A4(new_n874), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n889), .B1(new_n896), .B2(G148gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n887), .B1(new_n888), .B2(new_n897), .ZN(G1345gat));
  NOR2_X1   g697(.A1(new_n878), .A2(new_n248), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT122), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n691), .A2(new_n374), .ZN(new_n901));
  AOI22_X1  g700(.A1(new_n900), .A2(new_n374), .B1(new_n882), .B2(new_n901), .ZN(G1346gat));
  AOI21_X1  g701(.A(G162gat), .B1(new_n886), .B2(new_n302), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n301), .A2(new_n375), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n903), .B1(new_n882), .B2(new_n904), .ZN(G1347gat));
  AOI21_X1  g704(.A(KEYINPUT123), .B1(new_n823), .B2(new_n493), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907));
  AOI211_X1 g706(.A(new_n907), .B(new_n676), .C1(new_n821), .C2(new_n822), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n616), .B(new_n824), .C1(new_n906), .C2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n507), .A3(new_n356), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n493), .A2(new_n616), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(new_n703), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n646), .B1(new_n913), .B2(KEYINPUT124), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n913), .A2(KEYINPUT124), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n823), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(G169gat), .B1(new_n916), .B2(new_n357), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n911), .A2(new_n917), .ZN(G1348gat));
  NOR3_X1   g717(.A1(new_n916), .A2(new_n508), .A3(new_n326), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n910), .A2(new_n325), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n920), .B2(new_n508), .ZN(G1349gat));
  OAI21_X1  g720(.A(G183gat), .B1(new_n916), .B2(new_n691), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n247), .A2(new_n538), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n909), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT60), .ZN(G1350gat));
  NOR3_X1   g724(.A1(new_n909), .A2(G190gat), .A3(new_n301), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n823), .A2(new_n302), .A3(new_n914), .A4(new_n915), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n927), .A2(new_n928), .A3(G190gat), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n928), .B1(new_n927), .B2(G190gat), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT125), .B1(new_n926), .B2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n931), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n929), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n676), .B1(new_n821), .B2(new_n822), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT123), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n938), .A2(new_n525), .A3(new_n616), .A4(new_n824), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n935), .B(new_n936), .C1(new_n939), .C2(new_n301), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n933), .A2(new_n940), .ZN(G1351gat));
  AND2_X1   g740(.A1(new_n890), .A2(new_n895), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n614), .A2(new_n912), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(G197gat), .B1(new_n944), .B2(new_n357), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n614), .A2(new_n572), .A3(new_n433), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n938), .A2(KEYINPUT126), .A3(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(G197gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n946), .B1(new_n906), .B2(new_n908), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n947), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n945), .B1(new_n357), .B2(new_n952), .ZN(G1352gat));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n942), .A2(new_n954), .A3(new_n325), .A4(new_n943), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n890), .A2(new_n895), .A3(new_n325), .A4(new_n943), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(KEYINPUT127), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n955), .A2(G204gat), .A3(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n949), .ZN(new_n959));
  INV_X1    g758(.A(G204gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(new_n960), .A3(new_n325), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(KEYINPUT62), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n959), .A2(new_n963), .A3(new_n960), .A4(new_n325), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n958), .A2(new_n962), .A3(new_n964), .ZN(G1353gat));
  NAND4_X1  g764(.A1(new_n947), .A2(new_n951), .A3(new_n238), .A4(new_n247), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n890), .A2(new_n895), .A3(new_n247), .A4(new_n943), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n967), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n968));
  AOI21_X1  g767(.A(KEYINPUT63), .B1(new_n967), .B2(G211gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(G1354gat));
  NAND3_X1  g769(.A1(new_n947), .A2(new_n951), .A3(new_n302), .ZN(new_n971));
  INV_X1    g770(.A(G218gat), .ZN(new_n972));
  INV_X1    g771(.A(new_n944), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n301), .A2(new_n972), .ZN(new_n974));
  AOI22_X1  g773(.A1(new_n971), .A2(new_n972), .B1(new_n973), .B2(new_n974), .ZN(G1355gat));
endmodule


