

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  NOR2_X1 U323 ( .A1(n360), .A2(n546), .ZN(n362) );
  OR2_X1 U324 ( .A1(n481), .A2(n553), .ZN(n482) );
  XNOR2_X1 U325 ( .A(n556), .B(KEYINPUT79), .ZN(n535) );
  AND2_X1 U326 ( .A1(G227GAT), .A2(G233GAT), .ZN(n291) );
  XOR2_X1 U327 ( .A(n331), .B(KEYINPUT9), .Z(n292) );
  INV_X1 U328 ( .A(KEYINPUT111), .ZN(n361) );
  XNOR2_X1 U329 ( .A(n362), .B(n361), .ZN(n369) );
  XNOR2_X1 U330 ( .A(n434), .B(n291), .ZN(n435) );
  XNOR2_X1 U331 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U332 ( .A(n444), .B(n443), .Z(n518) );
  XNOR2_X1 U333 ( .A(n487), .B(n486), .ZN(n497) );
  NOR2_X1 U334 ( .A1(n513), .A2(n497), .ZN(n489) );
  XNOR2_X1 U335 ( .A(n446), .B(G190GAT), .ZN(n447) );
  XNOR2_X1 U336 ( .A(n448), .B(n447), .ZN(G1351GAT) );
  INV_X1 U337 ( .A(KEYINPUT68), .ZN(n295) );
  XOR2_X1 U338 ( .A(G92GAT), .B(G218GAT), .Z(n294) );
  XNOR2_X1 U339 ( .A(G36GAT), .B(G190GAT), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n382) );
  XNOR2_X1 U341 ( .A(n295), .B(n382), .ZN(n297) );
  XOR2_X1 U342 ( .A(G50GAT), .B(G162GAT), .Z(n422) );
  XNOR2_X1 U343 ( .A(G134GAT), .B(n422), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n302) );
  XOR2_X1 U345 ( .A(KEYINPUT75), .B(G85GAT), .Z(n299) );
  XNOR2_X1 U346 ( .A(G99GAT), .B(G106GAT), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n331) );
  NAND2_X1 U348 ( .A1(G232GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n292), .B(n300), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n310) );
  XOR2_X1 U351 ( .A(KEYINPUT71), .B(KEYINPUT8), .Z(n304) );
  XNOR2_X1 U352 ( .A(G43GAT), .B(G29GAT), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U354 ( .A(KEYINPUT7), .B(n305), .Z(n355) );
  XOR2_X1 U355 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n307) );
  XNOR2_X1 U356 ( .A(KEYINPUT11), .B(KEYINPUT78), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U358 ( .A(n355), .B(n308), .Z(n309) );
  XNOR2_X1 U359 ( .A(n310), .B(n309), .ZN(n556) );
  XOR2_X1 U360 ( .A(KEYINPUT67), .B(KEYINPUT45), .Z(n326) );
  XNOR2_X1 U361 ( .A(G71GAT), .B(G78GAT), .ZN(n311) );
  XNOR2_X1 U362 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n327) );
  XNOR2_X1 U363 ( .A(n311), .B(n327), .ZN(n324) );
  XOR2_X1 U364 ( .A(G8GAT), .B(G183GAT), .Z(n376) );
  XOR2_X1 U365 ( .A(G22GAT), .B(G155GAT), .Z(n415) );
  XOR2_X1 U366 ( .A(n376), .B(n415), .Z(n313) );
  NAND2_X1 U367 ( .A1(G231GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U369 ( .A(KEYINPUT12), .B(KEYINPUT80), .Z(n315) );
  XNOR2_X1 U370 ( .A(KEYINPUT81), .B(KEYINPUT15), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U372 ( .A(n317), .B(n316), .Z(n322) );
  XOR2_X1 U373 ( .A(G15GAT), .B(G127GAT), .Z(n429) );
  XOR2_X1 U374 ( .A(KEYINPUT14), .B(G64GAT), .Z(n319) );
  XNOR2_X1 U375 ( .A(G1GAT), .B(G211GAT), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n429), .B(n320), .ZN(n321) );
  XNOR2_X1 U378 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U379 ( .A(n324), .B(n323), .Z(n553) );
  INV_X1 U380 ( .A(n553), .ZN(n580) );
  XNOR2_X1 U381 ( .A(KEYINPUT36), .B(n535), .ZN(n481) );
  NOR2_X1 U382 ( .A1(n580), .A2(n481), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n342) );
  XNOR2_X1 U384 ( .A(G204GAT), .B(G92GAT), .ZN(n328) );
  XOR2_X1 U385 ( .A(n328), .B(n327), .Z(n341) );
  XOR2_X1 U386 ( .A(G176GAT), .B(G64GAT), .Z(n373) );
  XOR2_X1 U387 ( .A(G148GAT), .B(G78GAT), .Z(n421) );
  XOR2_X1 U388 ( .A(n373), .B(n421), .Z(n330) );
  NAND2_X1 U389 ( .A1(G230GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U390 ( .A(n330), .B(n329), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n331), .B(KEYINPUT32), .ZN(n332) );
  XNOR2_X1 U392 ( .A(n332), .B(KEYINPUT31), .ZN(n333) );
  XOR2_X1 U393 ( .A(n334), .B(n333), .Z(n339) );
  XOR2_X1 U394 ( .A(G120GAT), .B(G71GAT), .Z(n428) );
  XOR2_X1 U395 ( .A(KEYINPUT76), .B(KEYINPUT33), .Z(n336) );
  XNOR2_X1 U396 ( .A(KEYINPUT77), .B(KEYINPUT74), .ZN(n335) );
  XNOR2_X1 U397 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U398 ( .A(n428), .B(n337), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U400 ( .A(n341), .B(n340), .Z(n575) );
  AND2_X1 U401 ( .A1(n342), .A2(n575), .ZN(n343) );
  XOR2_X1 U402 ( .A(n343), .B(KEYINPUT110), .Z(n360) );
  XOR2_X1 U403 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n345) );
  XNOR2_X1 U404 ( .A(G141GAT), .B(G8GAT), .ZN(n344) );
  XNOR2_X1 U405 ( .A(n345), .B(n344), .ZN(n359) );
  XOR2_X1 U406 ( .A(G22GAT), .B(G197GAT), .Z(n347) );
  XNOR2_X1 U407 ( .A(G36GAT), .B(G50GAT), .ZN(n346) );
  XNOR2_X1 U408 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U409 ( .A(n348), .B(G15GAT), .Z(n350) );
  XOR2_X1 U410 ( .A(G113GAT), .B(G1GAT), .Z(n399) );
  XNOR2_X1 U411 ( .A(G169GAT), .B(n399), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U413 ( .A(KEYINPUT70), .B(KEYINPUT30), .Z(n352) );
  NAND2_X1 U414 ( .A1(G229GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U415 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U416 ( .A(n354), .B(n353), .Z(n357) );
  XNOR2_X1 U417 ( .A(n355), .B(KEYINPUT29), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U419 ( .A(n359), .B(n358), .Z(n546) );
  XNOR2_X1 U420 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n575), .B(n363), .ZN(n548) );
  NAND2_X1 U422 ( .A1(n546), .A2(n548), .ZN(n364) );
  XNOR2_X1 U423 ( .A(KEYINPUT46), .B(n364), .ZN(n365) );
  NAND2_X1 U424 ( .A1(n365), .A2(n580), .ZN(n366) );
  NOR2_X1 U425 ( .A1(n556), .A2(n366), .ZN(n367) );
  XOR2_X1 U426 ( .A(KEYINPUT47), .B(n367), .Z(n368) );
  NOR2_X1 U427 ( .A1(n369), .A2(n368), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n370), .B(KEYINPUT48), .ZN(n543) );
  XOR2_X1 U429 ( .A(G204GAT), .B(G211GAT), .Z(n372) );
  XNOR2_X1 U430 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n412) );
  XOR2_X1 U432 ( .A(n412), .B(n373), .Z(n375) );
  NAND2_X1 U433 ( .A1(G226GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n377) );
  XOR2_X1 U435 ( .A(n377), .B(n376), .Z(n379) );
  XNOR2_X1 U436 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n378) );
  XNOR2_X1 U437 ( .A(n379), .B(n378), .ZN(n384) );
  XOR2_X1 U438 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n381) );
  XNOR2_X1 U439 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n381), .B(n380), .ZN(n442) );
  XOR2_X1 U441 ( .A(n442), .B(n382), .Z(n383) );
  XOR2_X1 U442 ( .A(n384), .B(n383), .Z(n473) );
  INV_X1 U443 ( .A(n473), .ZN(n515) );
  NOR2_X1 U444 ( .A1(n543), .A2(n515), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n385), .B(KEYINPUT54), .ZN(n408) );
  XOR2_X1 U446 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n387) );
  XNOR2_X1 U447 ( .A(KEYINPUT88), .B(KEYINPUT6), .ZN(n386) );
  XNOR2_X1 U448 ( .A(n387), .B(n386), .ZN(n407) );
  XOR2_X1 U449 ( .A(G148GAT), .B(G162GAT), .Z(n389) );
  XNOR2_X1 U450 ( .A(G127GAT), .B(G120GAT), .ZN(n388) );
  XNOR2_X1 U451 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U452 ( .A(KEYINPUT89), .B(KEYINPUT4), .Z(n391) );
  XNOR2_X1 U453 ( .A(G155GAT), .B(KEYINPUT90), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U455 ( .A(n393), .B(n392), .Z(n405) );
  XNOR2_X1 U456 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n394), .B(KEYINPUT82), .ZN(n441) );
  XOR2_X1 U458 ( .A(n441), .B(G57GAT), .Z(n396) );
  NAND2_X1 U459 ( .A1(G225GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U460 ( .A(n396), .B(n395), .ZN(n403) );
  XOR2_X1 U461 ( .A(KEYINPUT2), .B(KEYINPUT86), .Z(n398) );
  XNOR2_X1 U462 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n397) );
  XNOR2_X1 U463 ( .A(n398), .B(n397), .ZN(n419) );
  XOR2_X1 U464 ( .A(G85GAT), .B(n419), .Z(n401) );
  XNOR2_X1 U465 ( .A(G29GAT), .B(n399), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U468 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U469 ( .A(n407), .B(n406), .Z(n470) );
  INV_X1 U470 ( .A(n470), .ZN(n513) );
  NAND2_X1 U471 ( .A1(n408), .A2(n513), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n409), .B(KEYINPUT65), .ZN(n571) );
  XOR2_X1 U473 ( .A(KEYINPUT85), .B(KEYINPUT87), .Z(n411) );
  XNOR2_X1 U474 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n410) );
  XNOR2_X1 U475 ( .A(n411), .B(n410), .ZN(n426) );
  XOR2_X1 U476 ( .A(n412), .B(KEYINPUT23), .Z(n414) );
  NAND2_X1 U477 ( .A1(G228GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U478 ( .A(n414), .B(n413), .ZN(n416) );
  XOR2_X1 U479 ( .A(n416), .B(n415), .Z(n418) );
  XNOR2_X1 U480 ( .A(G218GAT), .B(G106GAT), .ZN(n417) );
  XNOR2_X1 U481 ( .A(n418), .B(n417), .ZN(n420) );
  XOR2_X1 U482 ( .A(n420), .B(n419), .Z(n424) );
  XNOR2_X1 U483 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U485 ( .A(n426), .B(n425), .ZN(n462) );
  BUF_X1 U486 ( .A(n462), .Z(n453) );
  NAND2_X1 U487 ( .A1(n571), .A2(n453), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n427), .B(KEYINPUT55), .ZN(n445) );
  XOR2_X1 U489 ( .A(G190GAT), .B(G99GAT), .Z(n431) );
  XNOR2_X1 U490 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n431), .B(n430), .ZN(n436) );
  XOR2_X1 U492 ( .A(G176GAT), .B(G183GAT), .Z(n433) );
  XNOR2_X1 U493 ( .A(KEYINPUT20), .B(KEYINPUT83), .ZN(n432) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U495 ( .A(KEYINPUT84), .B(KEYINPUT66), .Z(n438) );
  XNOR2_X1 U496 ( .A(G43GAT), .B(G113GAT), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U498 ( .A(n440), .B(n439), .Z(n444) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n443) );
  INV_X1 U500 ( .A(n518), .ZN(n527) );
  NAND2_X1 U501 ( .A1(n445), .A2(n527), .ZN(n559) );
  NOR2_X1 U502 ( .A1(n535), .A2(n559), .ZN(n448) );
  XNOR2_X1 U503 ( .A(KEYINPUT121), .B(KEYINPUT58), .ZN(n446) );
  NOR2_X1 U504 ( .A1(n462), .A2(n527), .ZN(n450) );
  INV_X1 U505 ( .A(KEYINPUT26), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n541) );
  XOR2_X1 U507 ( .A(KEYINPUT27), .B(n473), .Z(n460) );
  NOR2_X1 U508 ( .A1(n541), .A2(n460), .ZN(n451) );
  XNOR2_X1 U509 ( .A(n451), .B(KEYINPUT94), .ZN(n458) );
  NOR2_X1 U510 ( .A1(n518), .A2(n515), .ZN(n452) );
  XNOR2_X1 U511 ( .A(n452), .B(KEYINPUT95), .ZN(n454) );
  NAND2_X1 U512 ( .A1(n454), .A2(n453), .ZN(n456) );
  XOR2_X1 U513 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n455) );
  XOR2_X1 U514 ( .A(n456), .B(n455), .Z(n457) );
  NOR2_X1 U515 ( .A1(n458), .A2(n457), .ZN(n459) );
  NOR2_X1 U516 ( .A1(n470), .A2(n459), .ZN(n464) );
  NOR2_X1 U517 ( .A1(n460), .A2(n513), .ZN(n461) );
  XOR2_X1 U518 ( .A(KEYINPUT93), .B(n461), .Z(n542) );
  XOR2_X1 U519 ( .A(KEYINPUT28), .B(n462), .Z(n478) );
  INV_X1 U520 ( .A(n478), .ZN(n522) );
  NAND2_X1 U521 ( .A1(n542), .A2(n522), .ZN(n525) );
  NOR2_X1 U522 ( .A1(n527), .A2(n525), .ZN(n463) );
  NOR2_X1 U523 ( .A1(n464), .A2(n463), .ZN(n465) );
  XOR2_X1 U524 ( .A(KEYINPUT97), .B(n465), .Z(n483) );
  NAND2_X1 U525 ( .A1(n553), .A2(n535), .ZN(n466) );
  XNOR2_X1 U526 ( .A(KEYINPUT16), .B(n466), .ZN(n467) );
  NOR2_X1 U527 ( .A1(n483), .A2(n467), .ZN(n499) );
  INV_X1 U528 ( .A(n546), .ZN(n572) );
  INV_X1 U529 ( .A(n575), .ZN(n468) );
  NOR2_X1 U530 ( .A1(n572), .A2(n468), .ZN(n485) );
  NAND2_X1 U531 ( .A1(n499), .A2(n485), .ZN(n469) );
  XOR2_X1 U532 ( .A(KEYINPUT98), .B(n469), .Z(n479) );
  NAND2_X1 U533 ( .A1(n479), .A2(n470), .ZN(n471) );
  XNOR2_X1 U534 ( .A(n471), .B(KEYINPUT34), .ZN(n472) );
  XNOR2_X1 U535 ( .A(G1GAT), .B(n472), .ZN(G1324GAT) );
  XOR2_X1 U536 ( .A(G8GAT), .B(KEYINPUT99), .Z(n475) );
  NAND2_X1 U537 ( .A1(n473), .A2(n479), .ZN(n474) );
  XNOR2_X1 U538 ( .A(n475), .B(n474), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(G15GAT), .B(KEYINPUT35), .Z(n477) );
  NAND2_X1 U540 ( .A1(n527), .A2(n479), .ZN(n476) );
  XNOR2_X1 U541 ( .A(n477), .B(n476), .ZN(G1326GAT) );
  NAND2_X1 U542 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U543 ( .A(n480), .B(G22GAT), .ZN(G1327GAT) );
  OR2_X2 U544 ( .A1(n483), .A2(n482), .ZN(n484) );
  XNOR2_X1 U545 ( .A(KEYINPUT37), .B(n484), .ZN(n512) );
  NAND2_X1 U546 ( .A1(n512), .A2(n485), .ZN(n487) );
  XNOR2_X1 U547 ( .A(KEYINPUT38), .B(KEYINPUT100), .ZN(n486) );
  XNOR2_X1 U548 ( .A(KEYINPUT101), .B(KEYINPUT39), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U550 ( .A(G29GAT), .B(n490), .Z(G1328GAT) );
  INV_X1 U551 ( .A(KEYINPUT102), .ZN(n492) );
  NOR2_X1 U552 ( .A1(n515), .A2(n497), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U554 ( .A(G36GAT), .B(n493), .ZN(G1329GAT) );
  NOR2_X1 U555 ( .A1(n518), .A2(n497), .ZN(n495) );
  XNOR2_X1 U556 ( .A(KEYINPUT103), .B(KEYINPUT40), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U558 ( .A(G43GAT), .B(n496), .ZN(G1330GAT) );
  NOR2_X1 U559 ( .A1(n522), .A2(n497), .ZN(n498) );
  XOR2_X1 U560 ( .A(G50GAT), .B(n498), .Z(G1331GAT) );
  INV_X1 U561 ( .A(n548), .ZN(n564) );
  NOR2_X1 U562 ( .A1(n546), .A2(n564), .ZN(n511) );
  NAND2_X1 U563 ( .A1(n499), .A2(n511), .ZN(n507) );
  NOR2_X1 U564 ( .A1(n513), .A2(n507), .ZN(n501) );
  XNOR2_X1 U565 ( .A(KEYINPUT42), .B(KEYINPUT104), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U567 ( .A(G57GAT), .B(n502), .Z(G1332GAT) );
  NOR2_X1 U568 ( .A1(n515), .A2(n507), .ZN(n504) );
  XNOR2_X1 U569 ( .A(G64GAT), .B(KEYINPUT105), .ZN(n503) );
  XNOR2_X1 U570 ( .A(n504), .B(n503), .ZN(G1333GAT) );
  NOR2_X1 U571 ( .A1(n518), .A2(n507), .ZN(n505) );
  XOR2_X1 U572 ( .A(KEYINPUT106), .B(n505), .Z(n506) );
  XNOR2_X1 U573 ( .A(G71GAT), .B(n506), .ZN(G1334GAT) );
  NOR2_X1 U574 ( .A1(n522), .A2(n507), .ZN(n509) );
  XNOR2_X1 U575 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U577 ( .A(G78GAT), .B(n510), .Z(G1335GAT) );
  NAND2_X1 U578 ( .A1(n512), .A2(n511), .ZN(n521) );
  NOR2_X1 U579 ( .A1(n513), .A2(n521), .ZN(n514) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n514), .Z(G1336GAT) );
  NOR2_X1 U581 ( .A1(n515), .A2(n521), .ZN(n516) );
  XOR2_X1 U582 ( .A(KEYINPUT108), .B(n516), .Z(n517) );
  XNOR2_X1 U583 ( .A(G92GAT), .B(n517), .ZN(G1337GAT) );
  NOR2_X1 U584 ( .A1(n518), .A2(n521), .ZN(n520) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(G1338GAT) );
  NOR2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U588 ( .A(KEYINPUT44), .B(n523), .Z(n524) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  NOR2_X1 U590 ( .A1(n543), .A2(n525), .ZN(n526) );
  NAND2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n536) );
  NOR2_X1 U592 ( .A1(n572), .A2(n536), .ZN(n528) );
  XOR2_X1 U593 ( .A(KEYINPUT112), .B(n528), .Z(n529) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n529), .ZN(G1340GAT) );
  NOR2_X1 U595 ( .A1(n564), .A2(n536), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  NOR2_X1 U598 ( .A1(n580), .A2(n536), .ZN(n533) );
  XNOR2_X1 U599 ( .A(KEYINPUT113), .B(KEYINPUT50), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  NOR2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n540) );
  XOR2_X1 U603 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n538) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT114), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  INV_X1 U607 ( .A(n541), .ZN(n570) );
  NAND2_X1 U608 ( .A1(n542), .A2(n570), .ZN(n544) );
  NOR2_X1 U609 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n545), .B(KEYINPUT116), .ZN(n557) );
  NAND2_X1 U611 ( .A1(n557), .A2(n546), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n547), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n550) );
  NAND2_X1 U614 ( .A1(n548), .A2(n557), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(n552) );
  XOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT53), .Z(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U618 ( .A1(n557), .A2(n553), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(KEYINPUT118), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G155GAT), .B(n555), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U622 ( .A(n558), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U623 ( .A1(n572), .A2(n559), .ZN(n561) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(KEYINPUT119), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n561), .B(n560), .ZN(G1348GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n563) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n566) );
  NOR2_X1 U629 ( .A1(n564), .A2(n559), .ZN(n565) );
  XOR2_X1 U630 ( .A(n566), .B(n565), .Z(G1349GAT) );
  NOR2_X1 U631 ( .A1(n580), .A2(n559), .ZN(n567) );
  XOR2_X1 U632 ( .A(G183GAT), .B(n567), .Z(G1350GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n585) );
  NOR2_X1 U637 ( .A1(n572), .A2(n585), .ZN(n573) );
  XOR2_X1 U638 ( .A(n574), .B(n573), .Z(G1352GAT) );
  NOR2_X1 U639 ( .A1(n585), .A2(n575), .ZN(n579) );
  XOR2_X1 U640 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n577) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n585), .ZN(n582) );
  XNOR2_X1 U645 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(G1354GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n587) );
  NOR2_X1 U650 ( .A1(n481), .A2(n585), .ZN(n586) );
  XOR2_X1 U651 ( .A(n587), .B(n586), .Z(G1355GAT) );
endmodule

