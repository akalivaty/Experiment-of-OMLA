//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n618, new_n619, new_n620, new_n621, new_n622, new_n624,
    new_n625, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910;
  INV_X1    g000(.A(KEYINPUT3), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(KEYINPUT22), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n202), .B1(new_n209), .B2(KEYINPUT29), .ZN(new_n210));
  INV_X1    g009(.A(G155gat), .ZN(new_n211));
  INV_X1    g010(.A(G162gat), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT2), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n211), .A2(new_n212), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT78), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n219), .A2(new_n220), .B1(G155gat), .B2(G162gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n217), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n218), .ZN(new_n223));
  INV_X1    g022(.A(new_n214), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(new_n215), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n213), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n228), .A2(KEYINPUT82), .B1(G228gat), .B2(G233gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT31), .B(G50gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n209), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n222), .A2(new_n226), .A3(new_n202), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT79), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n222), .A2(new_n226), .A3(KEYINPUT79), .A4(new_n202), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT29), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n228), .B1(new_n232), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G78gat), .B(G106gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n239), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n228), .B(new_n241), .C1(new_n232), .C2(new_n237), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n231), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(new_n231), .A3(new_n242), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n230), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT83), .B(G22gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n244), .A2(new_n230), .A3(new_n245), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n248), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n244), .A2(new_n230), .A3(new_n245), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n251), .B1(new_n252), .B2(new_n246), .ZN(new_n253));
  XOR2_X1   g052(.A(G15gat), .B(G43gat), .Z(new_n254));
  XNOR2_X1  g053(.A(G71gat), .B(G99gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258));
  NOR3_X1   g057(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262));
  OAI22_X1  g061(.A1(new_n259), .A2(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NOR4_X1   g062(.A1(KEYINPUT70), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n258), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT71), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n267), .B(new_n258), .C1(new_n263), .C2(new_n264), .ZN(new_n268));
  INV_X1    g067(.A(G183gat), .ZN(new_n269));
  NOR3_X1   g068(.A1(new_n269), .A2(KEYINPUT69), .A3(KEYINPUT27), .ZN(new_n270));
  NOR3_X1   g069(.A1(new_n270), .A2(KEYINPUT28), .A3(G190gat), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT27), .B1(new_n269), .B2(KEYINPUT69), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT27), .B(G183gat), .ZN(new_n273));
  INV_X1    g072(.A(G190gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n271), .A2(new_n272), .B1(new_n275), .B2(KEYINPUT28), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n266), .A2(new_n268), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT67), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n280), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(G183gat), .A2(G190gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT24), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n258), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n279), .A2(new_n281), .A3(new_n283), .A4(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(new_n282), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n290), .A2(KEYINPUT68), .A3(new_n279), .A4(new_n281), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n262), .A2(KEYINPUT23), .ZN(new_n292));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(G169gat), .B2(G176gat), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n292), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n288), .A2(new_n291), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT25), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT66), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT65), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n289), .A2(KEYINPUT65), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n283), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT64), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n278), .B(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n299), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT25), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n296), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n278), .B(KEYINPUT64), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n282), .B1(new_n285), .B2(new_n300), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n309), .A2(KEYINPUT66), .A3(new_n302), .A4(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n306), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n277), .A2(new_n298), .A3(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(G127gat), .B(G134gat), .Z(new_n314));
  INV_X1    g113(.A(G120gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G113gat), .ZN(new_n316));
  INV_X1    g115(.A(G113gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G120gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n318), .A3(KEYINPUT72), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT72), .B1(new_n316), .B2(new_n318), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n314), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n314), .A2(KEYINPUT1), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n318), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n317), .A2(KEYINPUT73), .A3(G120gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n316), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n323), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G227gat), .ZN(new_n331));
  INV_X1    g130(.A(G233gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n323), .A2(new_n329), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n277), .A2(new_n298), .A3(new_n312), .A4(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n330), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT33), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n257), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT34), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n330), .A2(new_n335), .ZN(new_n340));
  INV_X1    g139(.A(new_n333), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI211_X1 g141(.A(KEYINPUT34), .B(new_n333), .C1(new_n330), .C2(new_n335), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n338), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n336), .A2(KEYINPUT32), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n338), .B1(new_n342), .B2(new_n343), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n345), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n348), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n346), .B1(new_n350), .B2(new_n344), .ZN(new_n351));
  AND4_X1   g150(.A1(new_n250), .A2(new_n253), .A3(new_n349), .A4(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT35), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT4), .B1(new_n334), .B2(new_n227), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n222), .A2(new_n226), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT4), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n355), .A2(new_n356), .A3(new_n323), .A4(new_n329), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n354), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  OAI211_X1 g158(.A(KEYINPUT80), .B(KEYINPUT4), .C1(new_n334), .C2(new_n227), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n235), .A2(new_n236), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n227), .A2(KEYINPUT3), .B1(new_n323), .B2(new_n329), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT81), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n365), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(new_n362), .B2(new_n363), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n369), .A2(new_n359), .A3(new_n370), .A4(new_n360), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n334), .B(new_n355), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT5), .B1(new_n373), .B2(new_n365), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT0), .ZN(new_n378));
  XNOR2_X1  g177(.A(G57gat), .B(G85gat), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  INV_X1    g179(.A(KEYINPUT5), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n354), .A2(new_n357), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n369), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n376), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT6), .ZN(new_n385));
  INV_X1    g184(.A(new_n380), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n374), .B1(new_n367), .B2(new_n371), .ZN(new_n387));
  INV_X1    g186(.A(new_n383), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  OAI211_X1 g189(.A(KEYINPUT6), .B(new_n386), .C1(new_n387), .C2(new_n388), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n313), .A2(G226gat), .A3(G233gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(G226gat), .A2(G233gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT74), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT29), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n395), .B1(new_n313), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT75), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n393), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI211_X1 g198(.A(KEYINPUT75), .B(new_n395), .C1(new_n313), .C2(new_n396), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n209), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT76), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(G64gat), .B(G92gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  OAI211_X1 g205(.A(KEYINPUT76), .B(new_n209), .C1(new_n399), .C2(new_n400), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n313), .A2(new_n395), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT77), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n313), .A2(new_n396), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n394), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT77), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n313), .A2(new_n412), .A3(new_n395), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n409), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n232), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n403), .A2(new_n406), .A3(new_n407), .A4(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT30), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n401), .A2(new_n402), .B1(new_n414), .B2(new_n232), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n419), .A2(KEYINPUT30), .A3(new_n406), .A4(new_n407), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n407), .A3(new_n415), .ZN(new_n421));
  INV_X1    g220(.A(new_n406), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n418), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n352), .A2(new_n353), .A3(new_n392), .A4(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n392), .A2(new_n420), .A3(new_n423), .A4(new_n418), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n250), .A2(new_n253), .A3(new_n349), .A4(new_n351), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT35), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n250), .A2(new_n253), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT37), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n403), .A2(new_n433), .A3(new_n407), .A4(new_n415), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT85), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n419), .A2(KEYINPUT85), .A3(new_n433), .A4(new_n407), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n433), .B1(new_n414), .B2(new_n209), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n232), .B1(new_n399), .B2(new_n400), .ZN(new_n440));
  AOI211_X1 g239(.A(KEYINPUT38), .B(new_n406), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n390), .A2(new_n391), .A3(new_n416), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT38), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n406), .B1(new_n421), .B2(KEYINPUT37), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n446), .B1(new_n438), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n432), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n364), .A2(new_n382), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n368), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT39), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n452), .B1(new_n373), .B2(new_n365), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n450), .A2(new_n452), .A3(new_n368), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n380), .A3(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(KEYINPUT40), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n457), .A2(new_n389), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n424), .A2(KEYINPUT84), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT84), .B1(new_n424), .B2(new_n458), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n449), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n427), .A2(new_n431), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT36), .ZN(new_n464));
  INV_X1    g263(.A(new_n349), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n347), .B1(new_n345), .B2(new_n348), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n349), .A2(new_n351), .A3(KEYINPUT36), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n430), .B1(new_n462), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G113gat), .B(G141gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(G169gat), .B(G197gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(KEYINPUT12), .ZN(new_n477));
  NAND2_X1  g276(.A1(G29gat), .A2(G36gat), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT88), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  OR3_X1    g279(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G43gat), .B(G50gat), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n485), .A2(KEYINPUT87), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT15), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n487), .B1(new_n485), .B2(KEYINPUT87), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT89), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n484), .A2(new_n486), .A3(KEYINPUT89), .A4(new_n488), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n485), .A2(KEYINPUT15), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n484), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n486), .A2(new_n488), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT17), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G15gat), .B(G22gat), .ZN(new_n501));
  INV_X1    g300(.A(G1gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(KEYINPUT16), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT90), .ZN(new_n504));
  OAI221_X1 g303(.A(new_n503), .B1(new_n504), .B2(G8gat), .C1(new_n502), .C2(new_n501), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(G8gat), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n505), .B(new_n506), .Z(new_n507));
  AOI22_X1  g306(.A1(new_n491), .A2(new_n492), .B1(new_n496), .B2(new_n495), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT17), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n500), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n507), .A2(new_n508), .ZN(new_n511));
  NAND2_X1  g310(.A1(G229gat), .A2(G233gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT18), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n477), .B1(new_n515), .B2(KEYINPUT91), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n507), .B(new_n508), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n512), .B(KEYINPUT13), .Z(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT18), .A4(new_n512), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n515), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n513), .A2(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT91), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n524), .B1(new_n513), .B2(new_n514), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n523), .B(new_n520), .C1(new_n525), .C2(new_n477), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n471), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT92), .ZN(new_n529));
  OR2_X1    g328(.A1(G57gat), .A2(G64gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(G57gat), .A2(G64gat), .ZN(new_n531));
  AND2_X1   g330(.A1(G71gat), .A2(G78gat), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n530), .B(new_n531), .C1(new_n532), .C2(KEYINPUT9), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT93), .ZN(new_n534));
  NOR2_X1   g333(.A1(G71gat), .A2(G78gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n536), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT21), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G231gat), .A2(G233gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G127gat), .B(G155gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT20), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n544), .B(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n507), .B1(new_n541), .B2(new_n540), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT95), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n547), .B(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G183gat), .B(G211gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n550), .B(new_n553), .Z(new_n554));
  AND2_X1   g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(KEYINPUT41), .ZN(new_n556));
  XNOR2_X1  g355(.A(G134gat), .B(G162gat), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n556), .B(new_n557), .Z(new_n558));
  NAND2_X1  g357(.A1(G85gat), .A2(G92gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT7), .ZN(new_n560));
  NAND2_X1  g359(.A1(G99gat), .A2(G106gat), .ZN(new_n561));
  INV_X1    g360(.A(G85gat), .ZN(new_n562));
  INV_X1    g361(.A(G92gat), .ZN(new_n563));
  AOI22_X1  g362(.A1(KEYINPUT8), .A2(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G99gat), .B(G106gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n498), .A2(new_n567), .B1(KEYINPUT41), .B2(new_n555), .ZN(new_n568));
  INV_X1    g367(.A(new_n567), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n500), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n509), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n568), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G190gat), .B(G218gat), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n568), .B(new_n573), .C1(new_n570), .C2(new_n571), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n558), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n577), .B(KEYINPUT97), .Z(new_n578));
  NAND3_X1  g377(.A1(new_n575), .A2(new_n558), .A3(new_n576), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT96), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n554), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n539), .A2(new_n567), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT98), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT10), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G230gat), .A2(G233gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n540), .A2(new_n569), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT98), .B1(new_n539), .B2(new_n567), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT10), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n583), .ZN(new_n593));
  INV_X1    g392(.A(new_n588), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G120gat), .B(G148gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(G176gat), .B(G204gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n596), .B(new_n597), .Z(new_n598));
  NAND3_X1  g397(.A1(new_n592), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n599), .A2(KEYINPUT99), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(KEYINPUT99), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n592), .A2(new_n595), .ZN(new_n603));
  INV_X1    g402(.A(new_n598), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n582), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n529), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n392), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n424), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n612), .A2(G8gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT16), .B(G8gat), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(KEYINPUT42), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n616), .B1(KEYINPUT42), .B2(new_n615), .ZN(G1325gat));
  INV_X1    g416(.A(G15gat), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n465), .A2(new_n466), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n608), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n469), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n608), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n620), .B1(new_n622), .B2(new_n618), .ZN(G1326gat));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n431), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT43), .B(G22gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(G1327gat));
  NAND2_X1  g425(.A1(new_n578), .A2(new_n580), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n438), .A2(new_n447), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT38), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n443), .B1(new_n438), .B2(new_n441), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n431), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n424), .A2(new_n458), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT84), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n424), .A2(KEYINPUT84), .A3(new_n458), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n470), .B1(new_n631), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n426), .A2(new_n429), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n627), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n463), .A2(KEYINPUT100), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n427), .A2(new_n641), .A3(new_n431), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(new_n469), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n430), .B1(new_n462), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT101), .B(KEYINPUT44), .Z(new_n645));
  NOR2_X1   g444(.A1(new_n581), .A2(new_n645), .ZN(new_n646));
  AOI22_X1  g445(.A1(KEYINPUT44), .A2(new_n639), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n527), .ZN(new_n648));
  NOR4_X1   g447(.A1(new_n647), .A2(new_n648), .A3(new_n554), .A4(new_n606), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n649), .A2(new_n609), .ZN(new_n650));
  INV_X1    g449(.A(G29gat), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT45), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n550), .B(new_n553), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n600), .A2(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n655));
  AND4_X1   g454(.A1(new_n529), .A2(new_n654), .A3(new_n627), .A4(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n656), .A2(new_n651), .A3(new_n609), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n652), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(new_n653), .B2(new_n657), .ZN(G1328gat));
  AND2_X1   g458(.A1(new_n649), .A2(new_n424), .ZN(new_n660));
  INV_X1    g459(.A(G36gat), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n656), .A2(new_n661), .A3(new_n424), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n662), .B1(KEYINPUT46), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n664), .B1(KEYINPUT46), .B2(new_n663), .ZN(G1329gat));
  AOI21_X1  g464(.A(G43gat), .B1(new_n656), .B2(new_n619), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n649), .A2(G43gat), .A3(new_n621), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n668), .B(new_n670), .ZN(G1330gat));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n431), .ZN(new_n672));
  INV_X1    g471(.A(G50gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n432), .A2(new_n673), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n649), .A2(new_n675), .B1(KEYINPUT103), .B2(KEYINPUT48), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(KEYINPUT103), .A2(KEYINPUT48), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1331gat));
  INV_X1    g478(.A(new_n644), .ZN(new_n680));
  NOR4_X1   g479(.A1(new_n680), .A2(new_n527), .A3(new_n582), .A4(new_n655), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n609), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT104), .B(G57gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1332gat));
  AOI21_X1  g483(.A(new_n425), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT105), .Z(new_n687));
  NOR2_X1   g486(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1333gat));
  NAND2_X1  g488(.A1(new_n681), .A2(new_n621), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n465), .A2(new_n466), .A3(G71gat), .ZN(new_n691));
  AOI22_X1  g490(.A1(new_n690), .A2(G71gat), .B1(new_n681), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g492(.A1(new_n681), .A2(new_n431), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT106), .B(G78gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1335gat));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n654), .A2(new_n648), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT107), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n606), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n697), .B1(new_n647), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n700), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n703), .B1(new_n471), .B2(new_n627), .ZN(new_n704));
  INV_X1    g503(.A(new_n646), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n640), .A2(new_n469), .A3(new_n642), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n631), .A2(new_n636), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n705), .B1(new_n708), .B2(new_n430), .ZN(new_n709));
  OAI211_X1 g508(.A(KEYINPUT108), .B(new_n702), .C1(new_n704), .C2(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n701), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n609), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT109), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n562), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n713), .B2(new_n712), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n644), .A2(KEYINPUT51), .A3(new_n627), .A4(new_n699), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(KEYINPUT110), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n644), .A2(new_n627), .A3(new_n699), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT51), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n718), .B(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n609), .A2(new_n562), .A3(new_n606), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n715), .B1(new_n722), .B2(new_n723), .ZN(G1336gat));
  INV_X1    g523(.A(KEYINPUT52), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n647), .A2(new_n425), .A3(new_n700), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n425), .A2(G92gat), .A3(new_n655), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  OAI221_X1 g527(.A(new_n725), .B1(new_n563), .B2(new_n726), .C1(new_n722), .C2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n701), .A2(new_n424), .A3(new_n710), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G92gat), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT112), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(new_n721), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n731), .A2(KEYINPUT111), .B1(new_n727), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n730), .A2(new_n736), .A3(G92gat), .ZN(new_n737));
  AOI211_X1 g536(.A(KEYINPUT113), .B(new_n725), .C1(new_n735), .C2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT113), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n731), .A2(KEYINPUT111), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n734), .A2(new_n727), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n740), .A2(new_n737), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n739), .B1(new_n742), .B2(KEYINPUT52), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n729), .B1(new_n738), .B2(new_n743), .ZN(G1337gat));
  AND2_X1   g543(.A1(new_n711), .A2(new_n621), .ZN(new_n745));
  INV_X1    g544(.A(G99gat), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n619), .A2(new_n746), .A3(new_n606), .ZN(new_n747));
  OAI22_X1  g546(.A1(new_n745), .A2(new_n746), .B1(new_n722), .B2(new_n747), .ZN(G1338gat));
  INV_X1    g547(.A(KEYINPUT53), .ZN(new_n749));
  INV_X1    g548(.A(G106gat), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n647), .A2(new_n432), .A3(new_n700), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n432), .A2(G106gat), .A3(new_n655), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  OAI221_X1 g552(.A(new_n749), .B1(new_n750), .B2(new_n751), .C1(new_n722), .C2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n711), .A2(new_n431), .ZN(new_n755));
  AOI22_X1  g554(.A1(new_n755), .A2(G106gat), .B1(new_n734), .B2(new_n752), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n756), .B2(new_n749), .ZN(G1339gat));
  NAND2_X1  g556(.A1(new_n591), .A2(new_n589), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n590), .A2(KEYINPUT10), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n594), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(KEYINPUT54), .A3(new_n592), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT114), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n760), .A2(new_n763), .A3(KEYINPUT54), .A4(new_n592), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n604), .B1(new_n592), .B2(KEYINPUT54), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT115), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n768), .B(new_n604), .C1(new_n592), .C2(KEYINPUT54), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT116), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n762), .A2(new_n764), .B1(new_n767), .B2(new_n769), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n774), .A2(new_n775), .A3(KEYINPUT55), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n523), .A2(new_n477), .A3(new_n520), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n517), .A2(new_n518), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n512), .B1(new_n510), .B2(new_n511), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n476), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n782), .B1(new_n578), .B2(new_n580), .ZN(new_n783));
  AOI22_X1  g582(.A1(new_n774), .A2(KEYINPUT55), .B1(new_n601), .B2(new_n600), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n777), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n527), .B(new_n784), .C1(new_n773), .C2(new_n776), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n606), .A2(new_n781), .A3(new_n778), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n627), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n654), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n607), .A2(new_n648), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n428), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n424), .A2(new_n392), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(new_n648), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(new_n317), .ZN(G1340gat));
  NOR2_X1   g594(.A1(new_n793), .A2(new_n655), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(new_n315), .ZN(G1341gat));
  NOR2_X1   g596(.A1(new_n793), .A2(new_n654), .ZN(new_n798));
  XOR2_X1   g597(.A(new_n798), .B(G127gat), .Z(G1342gat));
  NOR2_X1   g598(.A1(new_n581), .A2(new_n424), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n392), .A2(G134gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n791), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n802), .B(KEYINPUT56), .Z(new_n803));
  OAI21_X1  g602(.A(G134gat), .B1(new_n793), .B2(new_n581), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(G1343gat));
  AOI21_X1  g604(.A(new_n432), .B1(new_n789), .B2(new_n790), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n469), .A2(new_n792), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n648), .A2(G141gat), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(KEYINPUT119), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n527), .B1(KEYINPUT55), .B2(new_n774), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n602), .B1(new_n771), .B2(new_n772), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n606), .A2(new_n816), .A3(new_n781), .A4(new_n778), .ZN(new_n817));
  OAI21_X1  g616(.A(KEYINPUT117), .B1(new_n655), .B2(new_n782), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT118), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n771), .A2(new_n772), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n784), .A2(new_n527), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n822), .A2(new_n823), .A3(new_n818), .A4(new_n817), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n820), .A2(new_n581), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n777), .A2(new_n783), .A3(new_n784), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n554), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n582), .A2(new_n527), .A3(new_n606), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n431), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT57), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n808), .B1(new_n806), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(new_n832), .A3(new_n527), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(G141gat), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT58), .B1(new_n812), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT58), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n811), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(G141gat), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n833), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n830), .A2(new_n832), .A3(KEYINPUT120), .A4(new_n527), .ZN(new_n841));
  AOI211_X1 g640(.A(KEYINPUT121), .B(new_n837), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n833), .A2(new_n839), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(G141gat), .A3(new_n841), .ZN(new_n845));
  INV_X1    g644(.A(new_n837), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n835), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT122), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n835), .B(KEYINPUT122), .C1(new_n842), .C2(new_n847), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(G1344gat));
  OR3_X1    g651(.A1(new_n807), .A2(KEYINPUT123), .A3(new_n831), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT123), .B1(new_n807), .B2(new_n831), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n829), .A2(new_n831), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n853), .B(new_n854), .C1(KEYINPUT124), .C2(new_n855), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n855), .A2(KEYINPUT124), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n858), .A2(new_n469), .A3(new_n606), .A4(new_n792), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n830), .A2(new_n832), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n606), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT59), .B1(new_n862), .B2(G148gat), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n655), .A2(G148gat), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n809), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n860), .A2(new_n865), .ZN(G1345gat));
  AOI21_X1  g665(.A(new_n211), .B1(new_n861), .B2(new_n554), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n654), .A2(G155gat), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n809), .B2(new_n868), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT125), .Z(G1346gat));
  NOR3_X1   g669(.A1(new_n621), .A2(G162gat), .A3(new_n392), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n806), .A2(new_n800), .A3(new_n871), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n861), .A2(new_n627), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n212), .ZN(G1347gat));
  NOR2_X1   g673(.A1(new_n425), .A2(new_n609), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n791), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n527), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n606), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(G176gat), .ZN(G1349gat));
  NOR2_X1   g680(.A1(new_n876), .A2(new_n654), .ZN(new_n882));
  MUX2_X1   g681(.A(G183gat), .B(new_n273), .S(new_n882), .Z(new_n883));
  INV_X1    g682(.A(KEYINPUT126), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT60), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT127), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n883), .B(new_n886), .ZN(G1350gat));
  OAI22_X1  g686(.A1(new_n876), .A2(new_n581), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n888), .B(new_n889), .ZN(G1351gat));
  NAND4_X1  g689(.A1(new_n469), .A2(new_n392), .A3(new_n424), .A4(new_n431), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n891), .B1(new_n789), .B2(new_n790), .ZN(new_n892));
  AOI21_X1  g691(.A(G197gat), .B1(new_n892), .B2(new_n527), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n875), .A2(new_n469), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n858), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n527), .A2(G197gat), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n893), .B1(new_n896), .B2(new_n897), .ZN(G1352gat));
  OAI21_X1  g697(.A(G204gat), .B1(new_n895), .B2(new_n655), .ZN(new_n899));
  INV_X1    g698(.A(G204gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n892), .A2(new_n900), .A3(new_n606), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n901), .B(KEYINPUT62), .Z(new_n902));
  NAND2_X1  g701(.A1(new_n899), .A2(new_n902), .ZN(G1353gat));
  NAND3_X1  g702(.A1(new_n892), .A2(new_n204), .A3(new_n554), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n554), .B(new_n894), .C1(new_n856), .C2(new_n857), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n905), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT63), .B1(new_n905), .B2(G211gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(G1354gat));
  OAI21_X1  g707(.A(G218gat), .B1(new_n895), .B2(new_n581), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n205), .A3(new_n627), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1355gat));
endmodule


