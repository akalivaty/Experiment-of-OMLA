

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765;

  NOR2_X1 U370 ( .A1(G953), .A2(G237), .ZN(n518) );
  XNOR2_X1 U371 ( .A(G146), .B(G125), .ZN(n491) );
  AND2_X4 U372 ( .A1(n620), .A2(n621), .ZN(n726) );
  NOR2_X2 U373 ( .A1(n549), .A2(n591), .ZN(n550) );
  XNOR2_X2 U374 ( .A(n748), .B(G146), .ZN(n504) );
  XNOR2_X2 U375 ( .A(n471), .B(n350), .ZN(n583) );
  XNOR2_X2 U376 ( .A(n567), .B(KEYINPUT45), .ZN(n731) );
  NAND2_X1 U377 ( .A1(n373), .A2(n372), .ZN(n371) );
  XNOR2_X1 U378 ( .A(KEYINPUT3), .B(KEYINPUT71), .ZN(n453) );
  INV_X1 U379 ( .A(G472), .ZN(n484) );
  AND2_X1 U380 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X2 U381 ( .A1(n374), .A2(n371), .ZN(n567) );
  NOR2_X1 U382 ( .A1(n598), .A2(n364), .ZN(n363) );
  NOR2_X1 U383 ( .A1(n562), .A2(n555), .ZN(n512) );
  XNOR2_X1 U384 ( .A(n439), .B(n382), .ZN(n693) );
  BUF_X1 U385 ( .A(n589), .Z(n542) );
  XNOR2_X1 U386 ( .A(n494), .B(n493), .ZN(n728) );
  NOR2_X1 U387 ( .A1(n632), .A2(G902), .ZN(n485) );
  XNOR2_X1 U388 ( .A(n488), .B(n487), .ZN(n494) );
  XNOR2_X1 U389 ( .A(n428), .B(n504), .ZN(n632) );
  XNOR2_X1 U390 ( .A(n424), .B(n423), .ZN(n531) );
  XNOR2_X1 U391 ( .A(n385), .B(n492), .ZN(n493) );
  XNOR2_X1 U392 ( .A(n452), .B(n451), .ZN(n479) );
  XNOR2_X1 U393 ( .A(n475), .B(G134), .ZN(n535) );
  XNOR2_X1 U394 ( .A(n462), .B(G128), .ZN(n475) );
  XNOR2_X1 U395 ( .A(n453), .B(G113), .ZN(n452) );
  XNOR2_X1 U396 ( .A(n347), .B(n468), .ZN(n739) );
  XOR2_X1 U397 ( .A(G104), .B(G107), .Z(n347) );
  XNOR2_X1 U398 ( .A(G137), .B(G140), .ZN(n502) );
  XNOR2_X2 U399 ( .A(n541), .B(KEYINPUT22), .ZN(n544) );
  XNOR2_X1 U400 ( .A(n369), .B(KEYINPUT73), .ZN(n395) );
  NAND2_X1 U401 ( .A1(n363), .A2(n362), .ZN(n369) );
  NOR2_X1 U402 ( .A1(G237), .A2(G902), .ZN(n469) );
  XNOR2_X1 U403 ( .A(G119), .B(G116), .ZN(n451) );
  NOR2_X1 U404 ( .A1(n683), .A2(n542), .ZN(n410) );
  NAND2_X1 U405 ( .A1(n409), .A2(KEYINPUT65), .ZN(n408) );
  INV_X1 U406 ( .A(n410), .ZN(n409) );
  XNOR2_X1 U407 ( .A(n507), .B(n506), .ZN(n508) );
  NOR2_X1 U408 ( .A1(G902), .A2(n719), .ZN(n509) );
  INV_X1 U409 ( .A(G469), .ZN(n506) );
  INV_X1 U410 ( .A(n666), .ZN(n455) );
  XOR2_X1 U411 ( .A(n739), .B(n478), .Z(n505) );
  XNOR2_X1 U412 ( .A(n587), .B(n416), .ZN(n415) );
  INV_X1 U413 ( .A(KEYINPUT83), .ZN(n416) );
  XNOR2_X1 U414 ( .A(n547), .B(n546), .ZN(n378) );
  INV_X1 U415 ( .A(KEYINPUT86), .ZN(n546) );
  NOR2_X1 U416 ( .A1(n653), .A2(n763), .ZN(n547) );
  XNOR2_X1 U417 ( .A(n614), .B(n613), .ZN(n615) );
  XOR2_X1 U418 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n467) );
  XNOR2_X1 U419 ( .A(KEYINPUT4), .B(KEYINPUT79), .ZN(n466) );
  XNOR2_X1 U420 ( .A(n465), .B(n464), .ZN(n402) );
  XNOR2_X1 U421 ( .A(n475), .B(n491), .ZN(n465) );
  AND2_X1 U422 ( .A1(n589), .A2(n421), .ZN(n590) );
  NOR2_X1 U423 ( .A1(n679), .A2(n422), .ZN(n421) );
  INV_X1 U424 ( .A(n588), .ZN(n422) );
  NAND2_X1 U425 ( .A1(n472), .A2(G214), .ZN(n694) );
  XNOR2_X1 U426 ( .A(n473), .B(KEYINPUT19), .ZN(n370) );
  NAND2_X1 U427 ( .A1(n583), .A2(n694), .ZN(n473) );
  INV_X1 U428 ( .A(KEYINPUT6), .ZN(n414) );
  XNOR2_X1 U429 ( .A(n427), .B(n483), .ZN(n428) );
  XNOR2_X1 U430 ( .A(n479), .B(n477), .ZN(n427) );
  XNOR2_X1 U431 ( .A(n479), .B(n401), .ZN(n738) );
  XNOR2_X1 U432 ( .A(KEYINPUT16), .B(G122), .ZN(n401) );
  XNOR2_X1 U433 ( .A(G131), .B(G104), .ZN(n521) );
  NAND2_X1 U434 ( .A1(G234), .A2(G237), .ZN(n460) );
  XNOR2_X1 U435 ( .A(n610), .B(n384), .ZN(n616) );
  INV_X1 U436 ( .A(KEYINPUT39), .ZN(n384) );
  INV_X1 U437 ( .A(n586), .ZN(n440) );
  NAND2_X1 U438 ( .A1(n448), .A2(n441), .ZN(n436) );
  NAND2_X1 U439 ( .A1(n439), .A2(KEYINPUT107), .ZN(n438) );
  NAND2_X1 U440 ( .A1(n407), .A2(n408), .ZN(n405) );
  NAND2_X1 U441 ( .A1(n408), .A2(n543), .ZN(n406) );
  INV_X1 U442 ( .A(KEYINPUT1), .ZN(n510) );
  NAND2_X1 U443 ( .A1(n430), .A2(n429), .ZN(n621) );
  INV_X1 U444 ( .A(KEYINPUT2), .ZN(n429) );
  XNOR2_X1 U445 ( .A(n420), .B(n504), .ZN(n719) );
  XNOR2_X1 U446 ( .A(n425), .B(n396), .ZN(n420) );
  XNOR2_X1 U447 ( .A(n503), .B(n397), .ZN(n396) );
  XOR2_X1 U448 ( .A(KEYINPUT91), .B(n628), .Z(n730) );
  NAND2_X1 U449 ( .A1(n377), .A2(n376), .ZN(n375) );
  NOR2_X1 U450 ( .A1(n762), .A2(KEYINPUT44), .ZN(n376) );
  NAND2_X1 U451 ( .A1(n378), .A2(KEYINPUT44), .ZN(n373) );
  XNOR2_X1 U452 ( .A(n499), .B(n498), .ZN(n577) );
  XNOR2_X1 U453 ( .A(n497), .B(n496), .ZN(n498) );
  NOR2_X1 U454 ( .A1(n728), .A2(G902), .ZN(n499) );
  INV_X1 U455 ( .A(KEYINPUT25), .ZN(n496) );
  XOR2_X1 U456 ( .A(G137), .B(KEYINPUT75), .Z(n481) );
  INV_X1 U457 ( .A(KEYINPUT48), .ZN(n388) );
  INV_X1 U458 ( .A(G143), .ZN(n462) );
  XNOR2_X1 U459 ( .A(G113), .B(G143), .ZN(n515) );
  XNOR2_X1 U460 ( .A(n418), .B(n520), .ZN(n522) );
  XNOR2_X1 U461 ( .A(n519), .B(n419), .ZN(n418) );
  INV_X1 U462 ( .A(KEYINPUT11), .ZN(n419) );
  XNOR2_X1 U463 ( .A(KEYINPUT15), .B(G902), .ZN(n617) );
  XNOR2_X1 U464 ( .A(n535), .B(n476), .ZN(n748) );
  XNOR2_X1 U465 ( .A(G131), .B(KEYINPUT4), .ZN(n476) );
  XNOR2_X1 U466 ( .A(n502), .B(KEYINPUT94), .ZN(n747) );
  INV_X1 U467 ( .A(KEYINPUT38), .ZN(n382) );
  NOR2_X1 U468 ( .A1(n445), .A2(KEYINPUT30), .ZN(n444) );
  INV_X1 U469 ( .A(n584), .ZN(n446) );
  XNOR2_X1 U470 ( .A(n458), .B(n457), .ZN(n558) );
  XNOR2_X1 U471 ( .A(n525), .B(G475), .ZN(n457) );
  OR2_X1 U472 ( .A1(n641), .A2(G902), .ZN(n458) );
  NOR2_X2 U473 ( .A1(n577), .A2(n572), .ZN(n684) );
  XNOR2_X1 U474 ( .A(G119), .B(G110), .ZN(n486) );
  XNOR2_X1 U475 ( .A(n514), .B(n351), .ZN(n385) );
  XNOR2_X1 U476 ( .A(G128), .B(KEYINPUT23), .ZN(n489) );
  XOR2_X1 U477 ( .A(KEYINPUT24), .B(KEYINPUT72), .Z(n490) );
  INV_X1 U478 ( .A(KEYINPUT8), .ZN(n423) );
  NAND2_X1 U479 ( .A1(n751), .A2(G234), .ZN(n424) );
  XNOR2_X1 U480 ( .A(G122), .B(KEYINPUT9), .ZN(n527) );
  XOR2_X1 U481 ( .A(KEYINPUT101), .B(KEYINPUT7), .Z(n528) );
  XNOR2_X1 U482 ( .A(G116), .B(G107), .ZN(n526) );
  XNOR2_X1 U483 ( .A(n747), .B(n398), .ZN(n397) );
  INV_X1 U484 ( .A(KEYINPUT78), .ZN(n398) );
  XNOR2_X1 U485 ( .A(n400), .B(n399), .ZN(n625) );
  XNOR2_X1 U486 ( .A(n402), .B(n349), .ZN(n399) );
  XNOR2_X1 U487 ( .A(n738), .B(n505), .ZN(n400) );
  NAND2_X1 U488 ( .A1(n380), .A2(n379), .ZN(n674) );
  INV_X1 U489 ( .A(n673), .ZN(n379) );
  XNOR2_X1 U490 ( .A(n590), .B(n412), .ZN(n593) );
  INV_X1 U491 ( .A(KEYINPUT28), .ZN(n412) );
  AND2_X1 U492 ( .A1(n348), .A2(n474), .ZN(n450) );
  XNOR2_X1 U493 ( .A(n558), .B(n383), .ZN(n560) );
  INV_X1 U494 ( .A(KEYINPUT100), .ZN(n383) );
  XOR2_X1 U495 ( .A(n632), .B(KEYINPUT62), .Z(n633) );
  XNOR2_X1 U496 ( .A(n641), .B(n640), .ZN(n642) );
  AND2_X1 U497 ( .A1(n616), .A2(n658), .ZN(n612) );
  XNOR2_X1 U498 ( .A(n601), .B(KEYINPUT111), .ZN(n759) );
  NOR2_X1 U499 ( .A1(n599), .A2(n448), .ZN(n413) );
  XNOR2_X1 U500 ( .A(n545), .B(KEYINPUT32), .ZN(n763) );
  NAND2_X1 U501 ( .A1(n562), .A2(n411), .ZN(n454) );
  INV_X1 U502 ( .A(n661), .ZN(n658) );
  NAND2_X1 U503 ( .A1(n440), .A2(n436), .ZN(n435) );
  NAND2_X1 U504 ( .A1(n356), .A2(n407), .ZN(n403) );
  XNOR2_X1 U505 ( .A(n719), .B(n459), .ZN(n720) );
  INV_X1 U506 ( .A(n679), .ZN(n411) );
  XNOR2_X1 U507 ( .A(n460), .B(KEYINPUT14), .ZN(n348) );
  XOR2_X1 U508 ( .A(n467), .B(n466), .Z(n349) );
  XOR2_X1 U509 ( .A(n470), .B(KEYINPUT92), .Z(n350) );
  XNOR2_X1 U510 ( .A(KEYINPUT67), .B(G101), .ZN(n477) );
  XOR2_X1 U511 ( .A(KEYINPUT95), .B(KEYINPUT84), .Z(n351) );
  AND2_X1 U512 ( .A1(n410), .A2(n543), .ZN(n352) );
  AND2_X1 U513 ( .A1(n566), .A2(n761), .ZN(n353) );
  NOR2_X1 U514 ( .A1(n667), .A2(n455), .ZN(n354) );
  OR2_X1 U515 ( .A1(n694), .A2(n447), .ZN(n355) );
  AND2_X1 U516 ( .A1(n352), .A2(n411), .ZN(n356) );
  OR2_X1 U517 ( .A1(n578), .A2(n454), .ZN(n357) );
  AND2_X1 U518 ( .A1(n446), .A2(n355), .ZN(n358) );
  AND2_X1 U519 ( .A1(n406), .A2(n411), .ZN(n359) );
  XOR2_X1 U520 ( .A(KEYINPUT88), .B(KEYINPUT0), .Z(n360) );
  INV_X1 U521 ( .A(KEYINPUT30), .ZN(n447) );
  INV_X1 U522 ( .A(KEYINPUT107), .ZN(n441) );
  INV_X1 U523 ( .A(KEYINPUT65), .ZN(n543) );
  XOR2_X1 U524 ( .A(KEYINPUT125), .B(n753), .Z(n361) );
  NAND2_X1 U525 ( .A1(n365), .A2(n366), .ZN(n362) );
  NAND2_X1 U526 ( .A1(n368), .A2(n367), .ZN(n364) );
  NOR2_X1 U527 ( .A1(n657), .A2(KEYINPUT82), .ZN(n365) );
  INV_X1 U528 ( .A(n594), .ZN(n366) );
  NAND2_X1 U529 ( .A1(n657), .A2(KEYINPUT82), .ZN(n367) );
  NAND2_X1 U530 ( .A1(n594), .A2(KEYINPUT82), .ZN(n368) );
  NAND2_X1 U531 ( .A1(n370), .A2(n450), .ZN(n449) );
  NAND2_X1 U532 ( .A1(n603), .A2(n370), .ZN(n595) );
  NAND2_X1 U533 ( .A1(n762), .A2(KEYINPUT44), .ZN(n372) );
  NAND2_X1 U534 ( .A1(n375), .A2(n353), .ZN(n374) );
  INV_X1 U535 ( .A(n378), .ZN(n377) );
  XNOR2_X2 U536 ( .A(n539), .B(KEYINPUT35), .ZN(n762) );
  INV_X1 U537 ( .A(n381), .ZN(n380) );
  NOR2_X2 U538 ( .A1(n731), .A2(n381), .ZN(n669) );
  XNOR2_X1 U539 ( .A(n381), .B(KEYINPUT77), .ZN(n432) );
  XNOR2_X1 U540 ( .A(n381), .B(n361), .ZN(n750) );
  NAND2_X2 U541 ( .A1(n456), .A2(n354), .ZN(n381) );
  XNOR2_X1 U542 ( .A(n391), .B(n615), .ZN(n390) );
  XNOR2_X1 U543 ( .A(n389), .B(n388), .ZN(n456) );
  NOR2_X1 U544 ( .A1(n544), .A2(n357), .ZN(n545) );
  INV_X1 U545 ( .A(n693), .ZN(n609) );
  NAND2_X1 U546 ( .A1(n693), .A2(n694), .ZN(n697) );
  NOR2_X2 U547 ( .A1(n593), .A2(n592), .ZN(n603) );
  NAND2_X1 U548 ( .A1(n576), .A2(n411), .ZN(n599) );
  NOR2_X1 U549 ( .A1(n442), .A2(n386), .ZN(n585) );
  NAND2_X1 U550 ( .A1(n443), .A2(n358), .ZN(n386) );
  NAND2_X1 U551 ( .A1(n585), .A2(n387), .ZN(n608) );
  NAND2_X1 U552 ( .A1(n551), .A2(n387), .ZN(n552) );
  XNOR2_X1 U553 ( .A(n550), .B(KEYINPUT96), .ZN(n387) );
  NAND2_X1 U554 ( .A1(n392), .A2(n390), .ZN(n389) );
  NAND2_X1 U555 ( .A1(n758), .A2(n764), .ZN(n391) );
  XNOR2_X1 U556 ( .A(n393), .B(n602), .ZN(n392) );
  NAND2_X1 U557 ( .A1(n395), .A2(n394), .ZN(n393) );
  INV_X1 U558 ( .A(n759), .ZN(n394) );
  NAND2_X1 U559 ( .A1(n404), .A2(n403), .ZN(n653) );
  NAND2_X1 U560 ( .A1(n405), .A2(n359), .ZN(n404) );
  INV_X1 U561 ( .A(n544), .ZN(n407) );
  NOR2_X1 U562 ( .A1(n544), .A2(n683), .ZN(n563) );
  NAND2_X1 U563 ( .A1(n726), .A2(G475), .ZN(n643) );
  XNOR2_X1 U564 ( .A(n413), .B(KEYINPUT36), .ZN(n600) );
  NAND2_X1 U565 ( .A1(n658), .A2(n573), .ZN(n574) );
  XNOR2_X1 U566 ( .A(n553), .B(n414), .ZN(n573) );
  NAND2_X1 U567 ( .A1(n726), .A2(G210), .ZN(n627) );
  NAND2_X1 U568 ( .A1(n426), .A2(n415), .ZN(n594) );
  INV_X1 U569 ( .A(n596), .ZN(n698) );
  XNOR2_X1 U570 ( .A(n523), .B(n524), .ZN(n641) );
  BUF_X1 U571 ( .A(n731), .Z(n417) );
  NAND2_X1 U572 ( .A1(n664), .A2(n661), .ZN(n596) );
  INV_X1 U573 ( .A(n731), .ZN(n431) );
  NOR2_X1 U574 ( .A1(n608), .A2(n438), .ZN(n437) );
  AND2_X2 U575 ( .A1(n434), .A2(n433), .ZN(n657) );
  XNOR2_X2 U576 ( .A(n591), .B(n511), .ZN(n683) );
  INV_X1 U577 ( .A(n505), .ZN(n425) );
  NAND2_X1 U578 ( .A1(n595), .A2(KEYINPUT47), .ZN(n426) );
  NAND2_X1 U579 ( .A1(n432), .A2(n431), .ZN(n430) );
  NAND2_X1 U580 ( .A1(n608), .A2(n441), .ZN(n433) );
  NOR2_X1 U581 ( .A1(n437), .A2(n435), .ZN(n434) );
  INV_X1 U582 ( .A(n448), .ZN(n439) );
  NAND2_X1 U583 ( .A1(n589), .A2(n444), .ZN(n443) );
  XNOR2_X2 U584 ( .A(n553), .B(KEYINPUT104), .ZN(n589) );
  NOR2_X1 U585 ( .A1(n589), .A2(n447), .ZN(n442) );
  INV_X1 U586 ( .A(n694), .ZN(n445) );
  INV_X1 U587 ( .A(n583), .ZN(n448) );
  XNOR2_X2 U588 ( .A(n449), .B(n360), .ZN(n556) );
  OR2_X1 U589 ( .A1(n560), .A2(n559), .ZN(n661) );
  NAND2_X1 U590 ( .A1(n560), .A2(n559), .ZN(n664) );
  XOR2_X1 U591 ( .A(n718), .B(n717), .Z(n459) );
  INV_X1 U592 ( .A(KEYINPUT46), .ZN(n613) );
  INV_X1 U593 ( .A(n477), .ZN(n478) );
  XNOR2_X1 U594 ( .A(n510), .B(KEYINPUT66), .ZN(n511) );
  INV_X1 U595 ( .A(n577), .ZN(n679) );
  XNOR2_X1 U596 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U597 ( .A(n721), .B(n720), .ZN(n722) );
  INV_X2 U598 ( .A(G953), .ZN(n463) );
  NOR2_X1 U599 ( .A1(G898), .A2(n463), .ZN(n743) );
  NAND2_X1 U600 ( .A1(n743), .A2(G902), .ZN(n461) );
  NAND2_X1 U601 ( .A1(G952), .A2(n463), .ZN(n569) );
  NAND2_X1 U602 ( .A1(n461), .A2(n569), .ZN(n474) );
  XNOR2_X2 U603 ( .A(n463), .B(KEYINPUT64), .ZN(n751) );
  NAND2_X1 U604 ( .A1(G224), .A2(n751), .ZN(n464) );
  XNOR2_X1 U605 ( .A(KEYINPUT76), .B(G110), .ZN(n468) );
  NAND2_X1 U606 ( .A1(n625), .A2(n617), .ZN(n471) );
  XOR2_X1 U607 ( .A(KEYINPUT74), .B(n469), .Z(n472) );
  NAND2_X1 U608 ( .A1(n472), .A2(G210), .ZN(n470) );
  XNOR2_X1 U609 ( .A(n556), .B(KEYINPUT93), .ZN(n548) );
  NAND2_X1 U610 ( .A1(n518), .A2(G210), .ZN(n480) );
  XNOR2_X1 U611 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U612 ( .A(n482), .B(KEYINPUT5), .Z(n483) );
  XNOR2_X2 U613 ( .A(n485), .B(n484), .ZN(n553) );
  INV_X1 U614 ( .A(n573), .ZN(n562) );
  NAND2_X1 U615 ( .A1(n531), .A2(G221), .ZN(n488) );
  XOR2_X1 U616 ( .A(n486), .B(n502), .Z(n487) );
  XNOR2_X1 U617 ( .A(n490), .B(n489), .ZN(n492) );
  XNOR2_X1 U618 ( .A(KEYINPUT10), .B(n491), .ZN(n514) );
  NAND2_X1 U619 ( .A1(G234), .A2(n617), .ZN(n495) );
  XNOR2_X1 U620 ( .A(KEYINPUT20), .B(n495), .ZN(n500) );
  NAND2_X1 U621 ( .A1(n500), .A2(G217), .ZN(n497) );
  NAND2_X1 U622 ( .A1(n500), .A2(G221), .ZN(n501) );
  XOR2_X1 U623 ( .A(n501), .B(KEYINPUT21), .Z(n678) );
  INV_X1 U624 ( .A(n678), .ZN(n572) );
  NAND2_X1 U625 ( .A1(G227), .A2(n751), .ZN(n503) );
  XNOR2_X1 U626 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n507) );
  XNOR2_X2 U627 ( .A(n509), .B(n508), .ZN(n591) );
  NAND2_X1 U628 ( .A1(n684), .A2(n683), .ZN(n555) );
  XNOR2_X1 U629 ( .A(KEYINPUT33), .B(n512), .ZN(n710) );
  NOR2_X1 U630 ( .A1(n548), .A2(n710), .ZN(n513) );
  XNOR2_X1 U631 ( .A(n513), .B(KEYINPUT34), .ZN(n538) );
  XNOR2_X1 U632 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n525) );
  XOR2_X1 U633 ( .A(G140), .B(G122), .Z(n516) );
  XNOR2_X1 U634 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U635 ( .A(n514), .B(n517), .ZN(n524) );
  XOR2_X1 U636 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n520) );
  NAND2_X1 U637 ( .A1(G214), .A2(n518), .ZN(n519) );
  XNOR2_X1 U638 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U639 ( .A(n526), .B(KEYINPUT102), .ZN(n530) );
  XNOR2_X1 U640 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U641 ( .A(n530), .B(n529), .Z(n533) );
  NAND2_X1 U642 ( .A1(G217), .A2(n531), .ZN(n532) );
  XNOR2_X1 U643 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U644 ( .A(n535), .B(n534), .ZN(n724) );
  NOR2_X1 U645 ( .A1(G902), .A2(n724), .ZN(n536) );
  XOR2_X1 U646 ( .A(G478), .B(n536), .Z(n559) );
  NAND2_X1 U647 ( .A1(n558), .A2(n559), .ZN(n586) );
  XOR2_X1 U648 ( .A(n586), .B(KEYINPUT80), .Z(n537) );
  NAND2_X1 U649 ( .A1(n538), .A2(n537), .ZN(n539) );
  OR2_X1 U650 ( .A1(n558), .A2(n559), .ZN(n696) );
  NOR2_X1 U651 ( .A1(n696), .A2(n572), .ZN(n540) );
  NAND2_X1 U652 ( .A1(n556), .A2(n540), .ZN(n541) );
  INV_X1 U653 ( .A(n683), .ZN(n578) );
  INV_X1 U654 ( .A(n548), .ZN(n551) );
  INV_X1 U655 ( .A(n684), .ZN(n549) );
  XNOR2_X1 U656 ( .A(n552), .B(KEYINPUT97), .ZN(n554) );
  INV_X1 U657 ( .A(n553), .ZN(n682) );
  NAND2_X1 U658 ( .A1(n554), .A2(n682), .ZN(n649) );
  NOR2_X1 U659 ( .A1(n682), .A2(n555), .ZN(n690) );
  NAND2_X1 U660 ( .A1(n690), .A2(n556), .ZN(n557) );
  XOR2_X1 U661 ( .A(KEYINPUT31), .B(n557), .Z(n663) );
  NAND2_X1 U662 ( .A1(n649), .A2(n663), .ZN(n561) );
  NAND2_X1 U663 ( .A1(n561), .A2(n596), .ZN(n566) );
  NAND2_X1 U664 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U665 ( .A1(n411), .A2(n564), .ZN(n565) );
  XNOR2_X1 U666 ( .A(n565), .B(KEYINPUT103), .ZN(n761) );
  NOR2_X1 U667 ( .A1(n751), .A2(G900), .ZN(n568) );
  NAND2_X1 U668 ( .A1(G902), .A2(n568), .ZN(n570) );
  NAND2_X1 U669 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U670 ( .A1(n348), .A2(n571), .ZN(n584) );
  NOR2_X1 U671 ( .A1(n572), .A2(n584), .ZN(n588) );
  NAND2_X1 U672 ( .A1(n588), .A2(n694), .ZN(n575) );
  NOR2_X1 U673 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U674 ( .A(n599), .B(KEYINPUT105), .ZN(n579) );
  NAND2_X1 U675 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U676 ( .A(n580), .B(KEYINPUT43), .ZN(n581) );
  XOR2_X1 U677 ( .A(KEYINPUT106), .B(n581), .Z(n582) );
  NOR2_X1 U678 ( .A1(n439), .A2(n582), .ZN(n667) );
  INV_X1 U679 ( .A(KEYINPUT68), .ZN(n602) );
  NAND2_X1 U680 ( .A1(n698), .A2(KEYINPUT47), .ZN(n587) );
  XNOR2_X1 U681 ( .A(n591), .B(KEYINPUT108), .ZN(n592) );
  INV_X1 U682 ( .A(n595), .ZN(n659) );
  NAND2_X1 U683 ( .A1(n659), .A2(n596), .ZN(n597) );
  NOR2_X1 U684 ( .A1(KEYINPUT47), .A2(n597), .ZN(n598) );
  NAND2_X1 U685 ( .A1(n600), .A2(n683), .ZN(n601) );
  INV_X1 U686 ( .A(n603), .ZN(n605) );
  NOR2_X1 U687 ( .A1(n697), .A2(n696), .ZN(n604) );
  XNOR2_X1 U688 ( .A(n604), .B(KEYINPUT41), .ZN(n709) );
  NOR2_X1 U689 ( .A1(n605), .A2(n709), .ZN(n607) );
  XOR2_X1 U690 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n606) );
  XNOR2_X1 U691 ( .A(n607), .B(n606), .ZN(n758) );
  NOR2_X1 U692 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U693 ( .A(KEYINPUT109), .B(KEYINPUT40), .ZN(n611) );
  XNOR2_X1 U694 ( .A(n612), .B(n611), .ZN(n764) );
  INV_X1 U695 ( .A(KEYINPUT85), .ZN(n614) );
  INV_X1 U696 ( .A(n664), .ZN(n654) );
  NAND2_X1 U697 ( .A1(n616), .A2(n654), .ZN(n666) );
  NAND2_X1 U698 ( .A1(n669), .A2(KEYINPUT2), .ZN(n619) );
  INV_X1 U699 ( .A(n617), .ZN(n618) );
  XOR2_X1 U700 ( .A(KEYINPUT54), .B(KEYINPUT118), .Z(n623) );
  XNOR2_X1 U701 ( .A(KEYINPUT87), .B(KEYINPUT55), .ZN(n622) );
  XNOR2_X1 U702 ( .A(n623), .B(n622), .ZN(n624) );
  XOR2_X1 U703 ( .A(n625), .B(n624), .Z(n626) );
  XNOR2_X1 U704 ( .A(n627), .B(n626), .ZN(n629) );
  NOR2_X1 U705 ( .A1(n751), .A2(G952), .ZN(n628) );
  INV_X1 U706 ( .A(n730), .ZN(n644) );
  NAND2_X1 U707 ( .A1(n629), .A2(n644), .ZN(n631) );
  INV_X1 U708 ( .A(KEYINPUT56), .ZN(n630) );
  XNOR2_X1 U709 ( .A(n631), .B(n630), .ZN(G51) );
  NAND2_X1 U710 ( .A1(n726), .A2(G472), .ZN(n634) );
  XNOR2_X1 U711 ( .A(n634), .B(n633), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n635), .A2(n644), .ZN(n639) );
  XOR2_X1 U713 ( .A(KEYINPUT112), .B(KEYINPUT90), .Z(n637) );
  INV_X1 U714 ( .A(KEYINPUT63), .ZN(n636) );
  XNOR2_X1 U715 ( .A(n639), .B(n638), .ZN(G57) );
  XOR2_X1 U716 ( .A(KEYINPUT59), .B(KEYINPUT89), .Z(n640) );
  XNOR2_X1 U717 ( .A(n643), .B(n642), .ZN(n645) );
  NAND2_X1 U718 ( .A1(n645), .A2(n644), .ZN(n647) );
  INV_X1 U719 ( .A(KEYINPUT60), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n647), .B(n646), .ZN(G60) );
  NOR2_X1 U721 ( .A1(n661), .A2(n649), .ZN(n648) );
  XOR2_X1 U722 ( .A(G104), .B(n648), .Z(G6) );
  NOR2_X1 U723 ( .A1(n664), .A2(n649), .ZN(n651) );
  XNOR2_X1 U724 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U726 ( .A(G107), .B(n652), .ZN(G9) );
  XOR2_X1 U727 ( .A(n653), .B(G110), .Z(G12) );
  XOR2_X1 U728 ( .A(G128), .B(KEYINPUT29), .Z(n656) );
  NAND2_X1 U729 ( .A1(n659), .A2(n654), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n656), .B(n655), .ZN(G30) );
  XOR2_X1 U731 ( .A(n657), .B(G143), .Z(G45) );
  NAND2_X1 U732 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n660), .B(G146), .ZN(G48) );
  NOR2_X1 U734 ( .A1(n661), .A2(n663), .ZN(n662) );
  XOR2_X1 U735 ( .A(G113), .B(n662), .Z(G15) );
  NOR2_X1 U736 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U737 ( .A(G116), .B(n665), .Z(G18) );
  XNOR2_X1 U738 ( .A(G134), .B(n666), .ZN(G36) );
  XNOR2_X1 U739 ( .A(G140), .B(n667), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n668), .B(KEYINPUT113), .ZN(G42) );
  NAND2_X1 U741 ( .A1(KEYINPUT81), .A2(KEYINPUT2), .ZN(n672) );
  NOR2_X1 U742 ( .A1(KEYINPUT2), .A2(KEYINPUT81), .ZN(n673) );
  INV_X1 U743 ( .A(n669), .ZN(n670) );
  NAND2_X1 U744 ( .A1(n673), .A2(n670), .ZN(n671) );
  NAND2_X1 U745 ( .A1(n672), .A2(n671), .ZN(n676) );
  NOR2_X1 U746 ( .A1(n417), .A2(n674), .ZN(n675) );
  NOR2_X1 U747 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U748 ( .A1(G953), .A2(n677), .ZN(n715) );
  NAND2_X1 U749 ( .A1(G952), .A2(n348), .ZN(n708) );
  NOR2_X1 U750 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U751 ( .A(n680), .B(KEYINPUT49), .ZN(n681) );
  NAND2_X1 U752 ( .A1(n682), .A2(n681), .ZN(n687) );
  NOR2_X1 U753 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U754 ( .A(n685), .B(KEYINPUT50), .ZN(n686) );
  NOR2_X1 U755 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U756 ( .A(n688), .B(KEYINPUT114), .ZN(n689) );
  NOR2_X1 U757 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U758 ( .A(KEYINPUT51), .B(n691), .Z(n692) );
  NOR2_X1 U759 ( .A1(n709), .A2(n692), .ZN(n704) );
  NOR2_X1 U760 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n701) );
  NOR2_X1 U762 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U763 ( .A(KEYINPUT115), .B(n699), .Z(n700) );
  NOR2_X1 U764 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U765 ( .A1(n702), .A2(n710), .ZN(n703) );
  NOR2_X1 U766 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U767 ( .A(KEYINPUT52), .B(n705), .ZN(n706) );
  XNOR2_X1 U768 ( .A(KEYINPUT116), .B(n706), .ZN(n707) );
  NOR2_X1 U769 ( .A1(n708), .A2(n707), .ZN(n712) );
  NOR2_X1 U770 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U771 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U772 ( .A(KEYINPUT117), .B(n713), .Z(n714) );
  NAND2_X1 U773 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U774 ( .A(KEYINPUT53), .B(n716), .Z(G75) );
  NAND2_X1 U775 ( .A1(n726), .A2(G469), .ZN(n721) );
  XOR2_X1 U776 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n718) );
  XNOR2_X1 U777 ( .A(KEYINPUT120), .B(KEYINPUT119), .ZN(n717) );
  NOR2_X1 U778 ( .A1(n730), .A2(n722), .ZN(G54) );
  NAND2_X1 U779 ( .A1(G478), .A2(n726), .ZN(n723) );
  XNOR2_X1 U780 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U781 ( .A1(n730), .A2(n725), .ZN(G63) );
  NAND2_X1 U782 ( .A1(G217), .A2(n726), .ZN(n727) );
  XNOR2_X1 U783 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U784 ( .A1(n730), .A2(n729), .ZN(G66) );
  NOR2_X1 U785 ( .A1(G953), .A2(n417), .ZN(n737) );
  XOR2_X1 U786 ( .A(KEYINPUT61), .B(KEYINPUT121), .Z(n733) );
  NAND2_X1 U787 ( .A1(G224), .A2(G953), .ZN(n732) );
  XNOR2_X1 U788 ( .A(n733), .B(n732), .ZN(n734) );
  NAND2_X1 U789 ( .A1(G898), .A2(n734), .ZN(n735) );
  XOR2_X1 U790 ( .A(KEYINPUT122), .B(n735), .Z(n736) );
  NOR2_X1 U791 ( .A1(n737), .A2(n736), .ZN(n746) );
  XOR2_X1 U792 ( .A(KEYINPUT123), .B(n738), .Z(n741) );
  XNOR2_X1 U793 ( .A(G101), .B(n739), .ZN(n740) );
  XNOR2_X1 U794 ( .A(n741), .B(n740), .ZN(n742) );
  NOR2_X1 U795 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U796 ( .A(KEYINPUT124), .B(n744), .Z(n745) );
  XNOR2_X1 U797 ( .A(n746), .B(n745), .ZN(G69) );
  XNOR2_X1 U798 ( .A(n747), .B(n514), .ZN(n749) );
  XNOR2_X1 U799 ( .A(n749), .B(n748), .ZN(n753) );
  NAND2_X1 U800 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U801 ( .A(n752), .B(KEYINPUT126), .ZN(n757) );
  XNOR2_X1 U802 ( .A(G227), .B(n753), .ZN(n754) );
  NAND2_X1 U803 ( .A1(n754), .A2(G900), .ZN(n755) );
  NAND2_X1 U804 ( .A1(G953), .A2(n755), .ZN(n756) );
  NAND2_X1 U805 ( .A1(n757), .A2(n756), .ZN(G72) );
  XNOR2_X1 U806 ( .A(n758), .B(G137), .ZN(G39) );
  XNOR2_X1 U807 ( .A(n759), .B(G125), .ZN(n760) );
  XNOR2_X1 U808 ( .A(n760), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U809 ( .A(G101), .B(n761), .ZN(G3) );
  XOR2_X1 U810 ( .A(G122), .B(n762), .Z(G24) );
  XOR2_X1 U811 ( .A(G119), .B(n763), .Z(G21) );
  XOR2_X1 U812 ( .A(G131), .B(n764), .Z(n765) );
  XNOR2_X1 U813 ( .A(KEYINPUT127), .B(n765), .ZN(G33) );
endmodule

