

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U546 ( .A1(n518), .A2(n514), .ZN(n886) );
  AND2_X1 U547 ( .A1(G160), .A2(G40), .ZN(n511) );
  BUF_X1 U548 ( .A(n692), .Z(n736) );
  NOR2_X1 U549 ( .A1(G651), .A2(n640), .ZN(n648) );
  NOR2_X2 U550 ( .A1(G2104), .A2(n518), .ZN(n887) );
  INV_X1 U551 ( .A(G2104), .ZN(n514) );
  NOR2_X4 U552 ( .A1(G2105), .A2(n514), .ZN(n890) );
  NAND2_X1 U553 ( .A1(G101), .A2(n890), .ZN(n513) );
  INV_X1 U554 ( .A(KEYINPUT23), .ZN(n512) );
  XNOR2_X1 U555 ( .A(n513), .B(n512), .ZN(n516) );
  INV_X1 U556 ( .A(G2105), .ZN(n518) );
  NAND2_X1 U557 ( .A1(n886), .A2(G113), .ZN(n515) );
  NAND2_X1 U558 ( .A1(n516), .A2(n515), .ZN(n522) );
  NOR2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n517) );
  XOR2_X2 U560 ( .A(KEYINPUT17), .B(n517), .Z(n891) );
  NAND2_X1 U561 ( .A1(G137), .A2(n891), .ZN(n520) );
  NAND2_X1 U562 ( .A1(G125), .A2(n887), .ZN(n519) );
  NAND2_X1 U563 ( .A1(n520), .A2(n519), .ZN(n521) );
  NOR2_X1 U564 ( .A1(n522), .A2(n521), .ZN(G160) );
  INV_X1 U565 ( .A(G651), .ZN(n531) );
  NOR2_X1 U566 ( .A1(G543), .A2(n531), .ZN(n524) );
  XNOR2_X1 U567 ( .A(KEYINPUT69), .B(KEYINPUT1), .ZN(n523) );
  XNOR2_X1 U568 ( .A(n524), .B(n523), .ZN(n647) );
  NAND2_X1 U569 ( .A1(G63), .A2(n647), .ZN(n527) );
  XOR2_X1 U570 ( .A(G543), .B(KEYINPUT0), .Z(n525) );
  XNOR2_X1 U571 ( .A(KEYINPUT68), .B(n525), .ZN(n640) );
  NAND2_X1 U572 ( .A1(G51), .A2(n648), .ZN(n526) );
  NAND2_X1 U573 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U574 ( .A(KEYINPUT6), .B(n528), .ZN(n537) );
  NOR2_X1 U575 ( .A1(G651), .A2(G543), .ZN(n529) );
  XOR2_X1 U576 ( .A(KEYINPUT67), .B(n529), .Z(n643) );
  NAND2_X1 U577 ( .A1(n643), .A2(G89), .ZN(n530) );
  XNOR2_X1 U578 ( .A(n530), .B(KEYINPUT4), .ZN(n533) );
  NOR2_X1 U579 ( .A1(n531), .A2(n640), .ZN(n644) );
  NAND2_X1 U580 ( .A1(G76), .A2(n644), .ZN(n532) );
  NAND2_X1 U581 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U582 ( .A(KEYINPUT5), .B(n534), .ZN(n535) );
  XNOR2_X1 U583 ( .A(KEYINPUT75), .B(n535), .ZN(n536) );
  NOR2_X1 U584 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U585 ( .A(KEYINPUT7), .B(n538), .Z(G168) );
  XOR2_X1 U586 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U587 ( .A1(G65), .A2(n647), .ZN(n540) );
  NAND2_X1 U588 ( .A1(G91), .A2(n643), .ZN(n539) );
  NAND2_X1 U589 ( .A1(n540), .A2(n539), .ZN(n544) );
  NAND2_X1 U590 ( .A1(G78), .A2(n644), .ZN(n542) );
  NAND2_X1 U591 ( .A1(G53), .A2(n648), .ZN(n541) );
  NAND2_X1 U592 ( .A1(n542), .A2(n541), .ZN(n543) );
  OR2_X1 U593 ( .A1(n544), .A2(n543), .ZN(G299) );
  NAND2_X1 U594 ( .A1(G138), .A2(n891), .ZN(n549) );
  NAND2_X1 U595 ( .A1(G114), .A2(n886), .ZN(n546) );
  NAND2_X1 U596 ( .A1(G126), .A2(n887), .ZN(n545) );
  NAND2_X1 U597 ( .A1(n546), .A2(n545), .ZN(n548) );
  AND2_X1 U598 ( .A1(G102), .A2(n890), .ZN(n547) );
  NOR2_X1 U599 ( .A1(n548), .A2(n547), .ZN(n683) );
  AND2_X1 U600 ( .A1(n549), .A2(n683), .ZN(G164) );
  XOR2_X1 U601 ( .A(G2430), .B(G2451), .Z(n551) );
  XNOR2_X1 U602 ( .A(KEYINPUT107), .B(G2443), .ZN(n550) );
  XNOR2_X1 U603 ( .A(n551), .B(n550), .ZN(n558) );
  XOR2_X1 U604 ( .A(G2435), .B(G2446), .Z(n553) );
  XNOR2_X1 U605 ( .A(G2427), .B(G2454), .ZN(n552) );
  XNOR2_X1 U606 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U607 ( .A(n554), .B(G2438), .Z(n556) );
  XNOR2_X1 U608 ( .A(G1341), .B(G1348), .ZN(n555) );
  XNOR2_X1 U609 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U610 ( .A(n558), .B(n557), .ZN(n559) );
  AND2_X1 U611 ( .A1(n559), .A2(G14), .ZN(G401) );
  NAND2_X1 U612 ( .A1(G64), .A2(n647), .ZN(n561) );
  NAND2_X1 U613 ( .A1(G52), .A2(n648), .ZN(n560) );
  NAND2_X1 U614 ( .A1(n561), .A2(n560), .ZN(n567) );
  NAND2_X1 U615 ( .A1(n643), .A2(G90), .ZN(n562) );
  XOR2_X1 U616 ( .A(KEYINPUT71), .B(n562), .Z(n564) );
  NAND2_X1 U617 ( .A1(n644), .A2(G77), .ZN(n563) );
  NAND2_X1 U618 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U619 ( .A(KEYINPUT9), .B(n565), .Z(n566) );
  NOR2_X1 U620 ( .A1(n567), .A2(n566), .ZN(G171) );
  AND2_X1 U621 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U622 ( .A(G120), .ZN(G236) );
  INV_X1 U623 ( .A(G132), .ZN(G219) );
  INV_X1 U624 ( .A(G96), .ZN(G221) );
  NAND2_X1 U625 ( .A1(G62), .A2(n647), .ZN(n569) );
  NAND2_X1 U626 ( .A1(G88), .A2(n643), .ZN(n568) );
  NAND2_X1 U627 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U628 ( .A1(G75), .A2(n644), .ZN(n571) );
  NAND2_X1 U629 ( .A1(G50), .A2(n648), .ZN(n570) );
  NAND2_X1 U630 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U631 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U632 ( .A(KEYINPUT84), .B(n574), .Z(G303) );
  NAND2_X1 U633 ( .A1(G7), .A2(G661), .ZN(n575) );
  XNOR2_X1 U634 ( .A(n575), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U635 ( .A(G223), .ZN(n834) );
  NAND2_X1 U636 ( .A1(n834), .A2(G567), .ZN(n576) );
  XOR2_X1 U637 ( .A(KEYINPUT11), .B(n576), .Z(G234) );
  NAND2_X1 U638 ( .A1(G56), .A2(n647), .ZN(n577) );
  XOR2_X1 U639 ( .A(KEYINPUT14), .B(n577), .Z(n583) );
  NAND2_X1 U640 ( .A1(n643), .A2(G81), .ZN(n578) );
  XNOR2_X1 U641 ( .A(n578), .B(KEYINPUT12), .ZN(n580) );
  NAND2_X1 U642 ( .A1(G68), .A2(n644), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U644 ( .A(KEYINPUT13), .B(n581), .Z(n582) );
  NOR2_X1 U645 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U646 ( .A1(n648), .A2(G43), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n585), .A2(n584), .ZN(n968) );
  XNOR2_X1 U648 ( .A(G860), .B(KEYINPUT73), .ZN(n598) );
  OR2_X1 U649 ( .A1(n968), .A2(n598), .ZN(G153) );
  INV_X1 U650 ( .A(G171), .ZN(G301) );
  NAND2_X1 U651 ( .A1(G66), .A2(n647), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G92), .A2(n643), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U654 ( .A1(G79), .A2(n644), .ZN(n589) );
  NAND2_X1 U655 ( .A1(G54), .A2(n648), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U658 ( .A(KEYINPUT74), .B(KEYINPUT15), .ZN(n592) );
  XNOR2_X1 U659 ( .A(n593), .B(n592), .ZN(n965) );
  NOR2_X1 U660 ( .A1(n965), .A2(G868), .ZN(n595) );
  INV_X1 U661 ( .A(G868), .ZN(n662) );
  NOR2_X1 U662 ( .A1(n662), .A2(G301), .ZN(n594) );
  NOR2_X1 U663 ( .A1(n595), .A2(n594), .ZN(G284) );
  NOR2_X1 U664 ( .A1(G286), .A2(n662), .ZN(n597) );
  NOR2_X1 U665 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U666 ( .A1(n597), .A2(n596), .ZN(G297) );
  NAND2_X1 U667 ( .A1(n598), .A2(G559), .ZN(n599) );
  INV_X1 U668 ( .A(n965), .ZN(n615) );
  NAND2_X1 U669 ( .A1(n599), .A2(n615), .ZN(n600) );
  XNOR2_X1 U670 ( .A(n600), .B(KEYINPUT76), .ZN(n601) );
  XNOR2_X1 U671 ( .A(KEYINPUT16), .B(n601), .ZN(G148) );
  NOR2_X1 U672 ( .A1(G868), .A2(n968), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n615), .A2(G868), .ZN(n602) );
  NOR2_X1 U674 ( .A1(G559), .A2(n602), .ZN(n603) );
  NOR2_X1 U675 ( .A1(n604), .A2(n603), .ZN(G282) );
  NAND2_X1 U676 ( .A1(G99), .A2(n890), .ZN(n606) );
  NAND2_X1 U677 ( .A1(G111), .A2(n886), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n607), .B(KEYINPUT77), .ZN(n609) );
  NAND2_X1 U680 ( .A1(G135), .A2(n891), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U682 ( .A1(n887), .A2(G123), .ZN(n610) );
  XOR2_X1 U683 ( .A(KEYINPUT18), .B(n610), .Z(n611) );
  NOR2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n918) );
  XNOR2_X1 U685 ( .A(n918), .B(G2096), .ZN(n614) );
  INV_X1 U686 ( .A(G2100), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n614), .A2(n613), .ZN(G156) );
  NAND2_X1 U688 ( .A1(n615), .A2(G559), .ZN(n616) );
  XNOR2_X1 U689 ( .A(n616), .B(n968), .ZN(n660) );
  NOR2_X1 U690 ( .A1(n660), .A2(G860), .ZN(n625) );
  NAND2_X1 U691 ( .A1(G67), .A2(n647), .ZN(n618) );
  NAND2_X1 U692 ( .A1(G93), .A2(n643), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U694 ( .A1(G55), .A2(n648), .ZN(n619) );
  XNOR2_X1 U695 ( .A(KEYINPUT79), .B(n619), .ZN(n620) );
  NOR2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n644), .A2(G80), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n663) );
  XOR2_X1 U699 ( .A(n663), .B(KEYINPUT78), .Z(n624) );
  XNOR2_X1 U700 ( .A(n625), .B(n624), .ZN(G145) );
  NAND2_X1 U701 ( .A1(n647), .A2(G61), .ZN(n626) );
  XNOR2_X1 U702 ( .A(n626), .B(KEYINPUT80), .ZN(n628) );
  NAND2_X1 U703 ( .A1(G86), .A2(n643), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U705 ( .A1(G73), .A2(n644), .ZN(n629) );
  XNOR2_X1 U706 ( .A(n629), .B(KEYINPUT81), .ZN(n630) );
  XNOR2_X1 U707 ( .A(n630), .B(KEYINPUT2), .ZN(n631) );
  NOR2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U709 ( .A(KEYINPUT82), .B(n633), .ZN(n636) );
  NAND2_X1 U710 ( .A1(n648), .A2(G48), .ZN(n634) );
  XOR2_X1 U711 ( .A(KEYINPUT83), .B(n634), .Z(n635) );
  NAND2_X1 U712 ( .A1(n636), .A2(n635), .ZN(G305) );
  NAND2_X1 U713 ( .A1(G49), .A2(n648), .ZN(n638) );
  NAND2_X1 U714 ( .A1(G74), .A2(G651), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U716 ( .A1(n647), .A2(n639), .ZN(n642) );
  NAND2_X1 U717 ( .A1(G87), .A2(n640), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n642), .A2(n641), .ZN(G288) );
  NAND2_X1 U719 ( .A1(G85), .A2(n643), .ZN(n646) );
  NAND2_X1 U720 ( .A1(G72), .A2(n644), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n652) );
  NAND2_X1 U722 ( .A1(G60), .A2(n647), .ZN(n650) );
  NAND2_X1 U723 ( .A1(G47), .A2(n648), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U726 ( .A(KEYINPUT70), .B(n653), .Z(G290) );
  XNOR2_X1 U727 ( .A(G288), .B(KEYINPUT19), .ZN(n655) );
  XNOR2_X1 U728 ( .A(G290), .B(G303), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n655), .B(n654), .ZN(n656) );
  XOR2_X1 U730 ( .A(n656), .B(G299), .Z(n657) );
  XNOR2_X1 U731 ( .A(n663), .B(n657), .ZN(n658) );
  XNOR2_X1 U732 ( .A(G305), .B(n658), .ZN(n906) );
  XOR2_X1 U733 ( .A(KEYINPUT85), .B(n906), .Z(n659) );
  XNOR2_X1 U734 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U735 ( .A1(n661), .A2(G868), .ZN(n665) );
  NAND2_X1 U736 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U737 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U738 ( .A1(G2084), .A2(G2078), .ZN(n666) );
  XOR2_X1 U739 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U740 ( .A1(n667), .A2(G2090), .ZN(n668) );
  XNOR2_X1 U741 ( .A(n668), .B(KEYINPUT86), .ZN(n669) );
  XNOR2_X1 U742 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U743 ( .A1(G2072), .A2(n670), .ZN(G158) );
  XOR2_X1 U744 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  XNOR2_X1 U745 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U746 ( .A1(G220), .A2(G219), .ZN(n672) );
  XNOR2_X1 U747 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n671) );
  XNOR2_X1 U748 ( .A(n672), .B(n671), .ZN(n673) );
  NOR2_X1 U749 ( .A1(n673), .A2(G218), .ZN(n674) );
  XOR2_X1 U750 ( .A(KEYINPUT88), .B(n674), .Z(n675) );
  NOR2_X1 U751 ( .A1(G221), .A2(n675), .ZN(n676) );
  XNOR2_X1 U752 ( .A(KEYINPUT89), .B(n676), .ZN(n838) );
  NAND2_X1 U753 ( .A1(n838), .A2(G2106), .ZN(n680) );
  NAND2_X1 U754 ( .A1(G69), .A2(G108), .ZN(n677) );
  NOR2_X1 U755 ( .A1(G236), .A2(n677), .ZN(n678) );
  NAND2_X1 U756 ( .A1(G57), .A2(n678), .ZN(n839) );
  NAND2_X1 U757 ( .A1(n839), .A2(G567), .ZN(n679) );
  NAND2_X1 U758 ( .A1(n680), .A2(n679), .ZN(n840) );
  NAND2_X1 U759 ( .A1(G483), .A2(G661), .ZN(n681) );
  NOR2_X1 U760 ( .A1(n840), .A2(n681), .ZN(n837) );
  NAND2_X1 U761 ( .A1(n837), .A2(G36), .ZN(G176) );
  XNOR2_X1 U762 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n833) );
  AND2_X1 U763 ( .A1(G138), .A2(n685), .ZN(n682) );
  NAND2_X1 U764 ( .A1(n891), .A2(n682), .ZN(n687) );
  INV_X1 U765 ( .A(G1384), .ZN(n685) );
  INV_X1 U766 ( .A(n683), .ZN(n684) );
  NAND2_X1 U767 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U768 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U769 ( .A(n688), .B(KEYINPUT65), .ZN(n758) );
  INV_X1 U770 ( .A(n758), .ZN(n689) );
  NAND2_X1 U771 ( .A1(n689), .A2(n511), .ZN(n690) );
  XNOR2_X1 U772 ( .A(KEYINPUT64), .B(n690), .ZN(n692) );
  XOR2_X1 U773 ( .A(G1996), .B(KEYINPUT94), .Z(n943) );
  NOR2_X1 U774 ( .A1(n692), .A2(n943), .ZN(n691) );
  XOR2_X1 U775 ( .A(n691), .B(KEYINPUT26), .Z(n694) );
  NAND2_X1 U776 ( .A1(n736), .A2(G1341), .ZN(n693) );
  NAND2_X1 U777 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U778 ( .A1(n968), .A2(n695), .ZN(n696) );
  XOR2_X1 U779 ( .A(KEYINPUT66), .B(n696), .Z(n702) );
  NOR2_X1 U780 ( .A1(n965), .A2(n702), .ZN(n697) );
  XNOR2_X1 U781 ( .A(n697), .B(KEYINPUT95), .ZN(n701) );
  INV_X1 U782 ( .A(n736), .ZN(n718) );
  NOR2_X1 U783 ( .A1(G1348), .A2(n718), .ZN(n699) );
  NOR2_X1 U784 ( .A1(G2067), .A2(n736), .ZN(n698) );
  NOR2_X1 U785 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U786 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U787 ( .A1(n965), .A2(n702), .ZN(n703) );
  NAND2_X1 U788 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U789 ( .A(n705), .B(KEYINPUT96), .ZN(n706) );
  INV_X1 U790 ( .A(n706), .ZN(n712) );
  NAND2_X1 U791 ( .A1(G2072), .A2(n718), .ZN(n707) );
  XOR2_X1 U792 ( .A(KEYINPUT27), .B(n707), .Z(n709) );
  NAND2_X1 U793 ( .A1(n736), .A2(G1956), .ZN(n708) );
  NAND2_X1 U794 ( .A1(n709), .A2(n708), .ZN(n713) );
  NOR2_X1 U795 ( .A1(G299), .A2(n713), .ZN(n710) );
  XOR2_X1 U796 ( .A(KEYINPUT97), .B(n710), .Z(n711) );
  NOR2_X1 U797 ( .A1(n712), .A2(n711), .ZN(n716) );
  NAND2_X1 U798 ( .A1(G299), .A2(n713), .ZN(n714) );
  XOR2_X1 U799 ( .A(KEYINPUT28), .B(n714), .Z(n715) );
  NOR2_X1 U800 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U801 ( .A(n717), .B(KEYINPUT29), .ZN(n722) );
  XOR2_X1 U802 ( .A(KEYINPUT25), .B(G2078), .Z(n942) );
  NAND2_X1 U803 ( .A1(n942), .A2(n718), .ZN(n720) );
  NAND2_X1 U804 ( .A1(n736), .A2(G1961), .ZN(n719) );
  NAND2_X1 U805 ( .A1(n720), .A2(n719), .ZN(n723) );
  OR2_X1 U806 ( .A1(n723), .A2(G301), .ZN(n721) );
  NAND2_X1 U807 ( .A1(n722), .A2(n721), .ZN(n735) );
  NAND2_X1 U808 ( .A1(G301), .A2(n723), .ZN(n724) );
  XNOR2_X1 U809 ( .A(n724), .B(KEYINPUT99), .ZN(n732) );
  NAND2_X1 U810 ( .A1(n736), .A2(G8), .ZN(n824) );
  NOR2_X1 U811 ( .A1(G1966), .A2(n824), .ZN(n725) );
  XOR2_X1 U812 ( .A(KEYINPUT93), .B(n725), .Z(n750) );
  NOR2_X1 U813 ( .A1(G2084), .A2(n736), .ZN(n726) );
  XNOR2_X1 U814 ( .A(n726), .B(KEYINPUT92), .ZN(n747) );
  NOR2_X1 U815 ( .A1(n750), .A2(n747), .ZN(n727) );
  XNOR2_X1 U816 ( .A(KEYINPUT98), .B(n727), .ZN(n728) );
  NAND2_X1 U817 ( .A1(n728), .A2(G8), .ZN(n729) );
  XNOR2_X1 U818 ( .A(KEYINPUT30), .B(n729), .ZN(n730) );
  NOR2_X1 U819 ( .A1(n730), .A2(G168), .ZN(n731) );
  NOR2_X1 U820 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U821 ( .A(KEYINPUT31), .B(n733), .Z(n734) );
  NAND2_X1 U822 ( .A1(n735), .A2(n734), .ZN(n748) );
  NAND2_X1 U823 ( .A1(n748), .A2(G286), .ZN(n742) );
  NOR2_X1 U824 ( .A1(n736), .A2(G2090), .ZN(n738) );
  NOR2_X1 U825 ( .A1(G1971), .A2(n824), .ZN(n737) );
  NOR2_X1 U826 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U827 ( .A1(G303), .A2(n739), .ZN(n740) );
  XOR2_X1 U828 ( .A(KEYINPUT101), .B(n740), .Z(n741) );
  NAND2_X1 U829 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U830 ( .A(KEYINPUT102), .B(n743), .ZN(n744) );
  NAND2_X1 U831 ( .A1(n744), .A2(G8), .ZN(n746) );
  XOR2_X1 U832 ( .A(KEYINPUT32), .B(KEYINPUT103), .Z(n745) );
  XNOR2_X1 U833 ( .A(n746), .B(n745), .ZN(n815) );
  NAND2_X1 U834 ( .A1(n747), .A2(G8), .ZN(n752) );
  XOR2_X1 U835 ( .A(n748), .B(KEYINPUT100), .Z(n749) );
  NOR2_X1 U836 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U837 ( .A1(n752), .A2(n751), .ZN(n816) );
  INV_X1 U838 ( .A(n824), .ZN(n753) );
  NAND2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n974) );
  AND2_X1 U840 ( .A1(n753), .A2(n974), .ZN(n754) );
  NOR2_X1 U841 ( .A1(KEYINPUT33), .A2(n754), .ZN(n757) );
  NOR2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n973) );
  NAND2_X1 U843 ( .A1(n973), .A2(KEYINPUT33), .ZN(n755) );
  NOR2_X1 U844 ( .A1(n755), .A2(n824), .ZN(n756) );
  NOR2_X1 U845 ( .A1(n757), .A2(n756), .ZN(n791) );
  XOR2_X1 U846 ( .A(G1981), .B(G305), .Z(n962) );
  XNOR2_X1 U847 ( .A(G1986), .B(G290), .ZN(n981) );
  NAND2_X1 U848 ( .A1(n758), .A2(n511), .ZN(n785) );
  INV_X1 U849 ( .A(n785), .ZN(n809) );
  AND2_X1 U850 ( .A1(n981), .A2(n809), .ZN(n788) );
  XNOR2_X1 U851 ( .A(G2067), .B(KEYINPUT37), .ZN(n806) );
  XNOR2_X1 U852 ( .A(KEYINPUT35), .B(KEYINPUT91), .ZN(n762) );
  NAND2_X1 U853 ( .A1(G116), .A2(n886), .ZN(n760) );
  NAND2_X1 U854 ( .A1(G128), .A2(n887), .ZN(n759) );
  NAND2_X1 U855 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U856 ( .A(n762), .B(n761), .ZN(n768) );
  NAND2_X1 U857 ( .A1(n891), .A2(G140), .ZN(n763) );
  XNOR2_X1 U858 ( .A(n763), .B(KEYINPUT90), .ZN(n765) );
  NAND2_X1 U859 ( .A1(G104), .A2(n890), .ZN(n764) );
  NAND2_X1 U860 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U861 ( .A(KEYINPUT34), .B(n766), .ZN(n767) );
  NOR2_X1 U862 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U863 ( .A(KEYINPUT36), .B(n769), .ZN(n877) );
  NOR2_X1 U864 ( .A1(n806), .A2(n877), .ZN(n933) );
  NAND2_X1 U865 ( .A1(n809), .A2(n933), .ZN(n804) );
  NAND2_X1 U866 ( .A1(G95), .A2(n890), .ZN(n771) );
  NAND2_X1 U867 ( .A1(G131), .A2(n891), .ZN(n770) );
  NAND2_X1 U868 ( .A1(n771), .A2(n770), .ZN(n775) );
  NAND2_X1 U869 ( .A1(G107), .A2(n886), .ZN(n773) );
  NAND2_X1 U870 ( .A1(G119), .A2(n887), .ZN(n772) );
  NAND2_X1 U871 ( .A1(n773), .A2(n772), .ZN(n774) );
  OR2_X1 U872 ( .A1(n775), .A2(n774), .ZN(n897) );
  AND2_X1 U873 ( .A1(n897), .A2(G1991), .ZN(n784) );
  NAND2_X1 U874 ( .A1(G141), .A2(n891), .ZN(n777) );
  NAND2_X1 U875 ( .A1(G117), .A2(n886), .ZN(n776) );
  NAND2_X1 U876 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U877 ( .A1(n890), .A2(G105), .ZN(n778) );
  XOR2_X1 U878 ( .A(KEYINPUT38), .B(n778), .Z(n779) );
  NOR2_X1 U879 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U880 ( .A1(n887), .A2(G129), .ZN(n781) );
  NAND2_X1 U881 ( .A1(n782), .A2(n781), .ZN(n876) );
  AND2_X1 U882 ( .A1(G1996), .A2(n876), .ZN(n783) );
  NOR2_X1 U883 ( .A1(n784), .A2(n783), .ZN(n924) );
  NOR2_X1 U884 ( .A1(n924), .A2(n785), .ZN(n801) );
  INV_X1 U885 ( .A(n801), .ZN(n786) );
  NAND2_X1 U886 ( .A1(n804), .A2(n786), .ZN(n787) );
  OR2_X1 U887 ( .A1(n788), .A2(n787), .ZN(n827) );
  INV_X1 U888 ( .A(n827), .ZN(n789) );
  AND2_X1 U889 ( .A1(n962), .A2(n789), .ZN(n790) );
  AND2_X1 U890 ( .A1(n791), .A2(n790), .ZN(n793) );
  AND2_X1 U891 ( .A1(n816), .A2(n793), .ZN(n792) );
  NAND2_X1 U892 ( .A1(n815), .A2(n792), .ZN(n814) );
  INV_X1 U893 ( .A(n793), .ZN(n797) );
  NOR2_X1 U894 ( .A1(G303), .A2(G1971), .ZN(n977) );
  NOR2_X1 U895 ( .A1(n973), .A2(n977), .ZN(n795) );
  INV_X1 U896 ( .A(KEYINPUT33), .ZN(n794) );
  AND2_X1 U897 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U898 ( .A1(n797), .A2(n796), .ZN(n812) );
  NOR2_X1 U899 ( .A1(G1996), .A2(n876), .ZN(n926) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n799) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n897), .ZN(n798) );
  XNOR2_X1 U902 ( .A(KEYINPUT104), .B(n798), .ZN(n919) );
  NOR2_X1 U903 ( .A1(n799), .A2(n919), .ZN(n800) );
  NOR2_X1 U904 ( .A1(n801), .A2(n800), .ZN(n802) );
  NOR2_X1 U905 ( .A1(n926), .A2(n802), .ZN(n803) );
  XNOR2_X1 U906 ( .A(KEYINPUT39), .B(n803), .ZN(n805) );
  NAND2_X1 U907 ( .A1(n805), .A2(n804), .ZN(n807) );
  NAND2_X1 U908 ( .A1(n806), .A2(n877), .ZN(n934) );
  NAND2_X1 U909 ( .A1(n807), .A2(n934), .ZN(n808) );
  XOR2_X1 U910 ( .A(KEYINPUT105), .B(n808), .Z(n810) );
  AND2_X1 U911 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U912 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U913 ( .A1(n814), .A2(n813), .ZN(n831) );
  NAND2_X1 U914 ( .A1(n816), .A2(n815), .ZN(n823) );
  NOR2_X1 U915 ( .A1(G2090), .A2(G303), .ZN(n817) );
  NAND2_X1 U916 ( .A1(G8), .A2(n817), .ZN(n821) );
  NOR2_X1 U917 ( .A1(G1981), .A2(G305), .ZN(n818) );
  XOR2_X1 U918 ( .A(n818), .B(KEYINPUT24), .Z(n819) );
  NOR2_X1 U919 ( .A1(n824), .A2(n819), .ZN(n825) );
  INV_X1 U920 ( .A(n825), .ZN(n820) );
  AND2_X1 U921 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U922 ( .A1(n823), .A2(n822), .ZN(n829) );
  NOR2_X1 U923 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U924 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U925 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U926 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U927 ( .A(n833), .B(n832), .ZN(G329) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U930 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n837), .A2(n836), .ZN(G188) );
  XOR2_X1 U933 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  XOR2_X1 U934 ( .A(G108), .B(KEYINPUT116), .Z(G238) );
  NOR2_X1 U936 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  INV_X1 U938 ( .A(n840), .ZN(G319) );
  XOR2_X1 U939 ( .A(KEYINPUT42), .B(G2090), .Z(n842) );
  XNOR2_X1 U940 ( .A(G2084), .B(G2072), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U942 ( .A(n843), .B(G2100), .Z(n845) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2078), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U945 ( .A(G2096), .B(KEYINPUT43), .Z(n847) );
  XNOR2_X1 U946 ( .A(KEYINPUT109), .B(G2678), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U948 ( .A(n849), .B(n848), .Z(G227) );
  XNOR2_X1 U949 ( .A(G1991), .B(KEYINPUT41), .ZN(n859) );
  XOR2_X1 U950 ( .A(G1976), .B(G1971), .Z(n851) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1986), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U953 ( .A(G1981), .B(G1956), .Z(n853) );
  XNOR2_X1 U954 ( .A(G1966), .B(G1961), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U956 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U957 ( .A(KEYINPUT110), .B(G2474), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U960 ( .A1(G100), .A2(n890), .ZN(n861) );
  NAND2_X1 U961 ( .A1(G112), .A2(n886), .ZN(n860) );
  NAND2_X1 U962 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n862), .B(KEYINPUT111), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G136), .A2(n891), .ZN(n863) );
  NAND2_X1 U965 ( .A1(n864), .A2(n863), .ZN(n867) );
  NAND2_X1 U966 ( .A1(n887), .A2(G124), .ZN(n865) );
  XOR2_X1 U967 ( .A(KEYINPUT44), .B(n865), .Z(n866) );
  NOR2_X1 U968 ( .A1(n867), .A2(n866), .ZN(G162) );
  NAND2_X1 U969 ( .A1(G103), .A2(n890), .ZN(n869) );
  NAND2_X1 U970 ( .A1(G139), .A2(n891), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n875) );
  NAND2_X1 U972 ( .A1(n887), .A2(G127), .ZN(n870) );
  XOR2_X1 U973 ( .A(KEYINPUT113), .B(n870), .Z(n872) );
  NAND2_X1 U974 ( .A1(n886), .A2(G115), .ZN(n871) );
  NAND2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U976 ( .A(KEYINPUT47), .B(n873), .Z(n874) );
  NOR2_X1 U977 ( .A1(n875), .A2(n874), .ZN(n914) );
  XNOR2_X1 U978 ( .A(n914), .B(n918), .ZN(n879) );
  XOR2_X1 U979 ( .A(n877), .B(n876), .Z(n878) );
  XNOR2_X1 U980 ( .A(n879), .B(n878), .ZN(n883) );
  XOR2_X1 U981 ( .A(KEYINPUT114), .B(KEYINPUT112), .Z(n881) );
  XNOR2_X1 U982 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n880) );
  XNOR2_X1 U983 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U984 ( .A(n883), .B(n882), .Z(n885) );
  XNOR2_X1 U985 ( .A(G164), .B(G162), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n885), .B(n884), .ZN(n901) );
  NAND2_X1 U987 ( .A1(G118), .A2(n886), .ZN(n889) );
  NAND2_X1 U988 ( .A1(G130), .A2(n887), .ZN(n888) );
  NAND2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n896) );
  NAND2_X1 U990 ( .A1(G106), .A2(n890), .ZN(n893) );
  NAND2_X1 U991 ( .A1(G142), .A2(n891), .ZN(n892) );
  NAND2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U993 ( .A(n894), .B(KEYINPUT45), .Z(n895) );
  NOR2_X1 U994 ( .A1(n896), .A2(n895), .ZN(n898) );
  XNOR2_X1 U995 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U996 ( .A(G160), .B(n899), .Z(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U998 ( .A1(G37), .A2(n902), .ZN(n903) );
  XOR2_X1 U999 ( .A(KEYINPUT115), .B(n903), .Z(G395) );
  XNOR2_X1 U1000 ( .A(n968), .B(G286), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(G171), .B(n965), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n907) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n908), .ZN(G397) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(G401), .A2(n910), .ZN(n911) );
  AND2_X1 U1008 ( .A1(G319), .A2(n911), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1013 ( .A(G2072), .B(n914), .Z(n916) );
  XOR2_X1 U1014 ( .A(G164), .B(G2078), .Z(n915) );
  NOR2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(KEYINPUT50), .B(n917), .ZN(n931) );
  XNOR2_X1 U1017 ( .A(G160), .B(G2084), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(KEYINPUT117), .B(n922), .ZN(n923) );
  NAND2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n929) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(KEYINPUT51), .B(n927), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n935) );
  NAND2_X1 U1028 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1029 ( .A(KEYINPUT52), .B(n936), .Z(n937) );
  XOR2_X1 U1030 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n957) );
  NAND2_X1 U1031 ( .A1(n937), .A2(n957), .ZN(n938) );
  NAND2_X1 U1032 ( .A1(n938), .A2(G29), .ZN(n992) );
  XNOR2_X1 U1033 ( .A(G1991), .B(G25), .ZN(n940) );
  XNOR2_X1 U1034 ( .A(G33), .B(G2072), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n949) );
  XOR2_X1 U1036 ( .A(G2067), .B(G26), .Z(n941) );
  NAND2_X1 U1037 ( .A1(n941), .A2(G28), .ZN(n947) );
  XOR2_X1 U1038 ( .A(n942), .B(G27), .Z(n945) );
  XNOR2_X1 U1039 ( .A(n943), .B(G32), .ZN(n944) );
  NAND2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(n950), .B(KEYINPUT53), .ZN(n953) );
  XOR2_X1 U1044 ( .A(G2084), .B(G34), .Z(n951) );
  XNOR2_X1 U1045 ( .A(KEYINPUT54), .B(n951), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n955) );
  XNOR2_X1 U1047 ( .A(G35), .B(G2090), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(n957), .B(n956), .ZN(n958) );
  NOR2_X1 U1050 ( .A1(G29), .A2(n958), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(KEYINPUT119), .B(n959), .ZN(n960) );
  NAND2_X1 U1052 ( .A1(n960), .A2(G11), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(n961), .B(KEYINPUT120), .ZN(n990) );
  XNOR2_X1 U1054 ( .A(G1966), .B(G168), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(n964), .B(KEYINPUT57), .ZN(n972) );
  XOR2_X1 U1057 ( .A(n965), .B(G1348), .Z(n967) );
  XNOR2_X1 U1058 ( .A(G171), .B(G1961), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(G1341), .B(n968), .ZN(n969) );
  NOR2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1062 ( .A1(n972), .A2(n971), .ZN(n986) );
  XNOR2_X1 U1063 ( .A(KEYINPUT121), .B(n973), .ZN(n975) );
  NAND2_X1 U1064 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1065 ( .A1(n977), .A2(n976), .ZN(n983) );
  NAND2_X1 U1066 ( .A1(G303), .A2(G1971), .ZN(n979) );
  XOR2_X1 U1067 ( .A(G1956), .B(G299), .Z(n978) );
  NAND2_X1 U1068 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1069 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1070 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1071 ( .A(KEYINPUT122), .B(n984), .ZN(n985) );
  NOR2_X1 U1072 ( .A1(n986), .A2(n985), .ZN(n988) );
  XOR2_X1 U1073 ( .A(G16), .B(KEYINPUT56), .Z(n987) );
  NOR2_X1 U1074 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1075 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1076 ( .A1(n992), .A2(n991), .ZN(n1020) );
  XOR2_X1 U1077 ( .A(G1961), .B(G5), .Z(n1004) );
  XNOR2_X1 U1078 ( .A(KEYINPUT59), .B(G1348), .ZN(n993) );
  XNOR2_X1 U1079 ( .A(n993), .B(G4), .ZN(n998) );
  XOR2_X1 U1080 ( .A(G1956), .B(KEYINPUT123), .Z(n994) );
  XNOR2_X1 U1081 ( .A(G20), .B(n994), .ZN(n996) );
  XNOR2_X1 U1082 ( .A(G6), .B(G1981), .ZN(n995) );
  NOR2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n1001) );
  XNOR2_X1 U1085 ( .A(KEYINPUT124), .B(G1341), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(G19), .B(n999), .ZN(n1000) );
  NOR2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(KEYINPUT60), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1089 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XNOR2_X1 U1090 ( .A(G21), .B(G1966), .ZN(n1005) );
  NOR2_X1 U1091 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(KEYINPUT125), .B(n1007), .ZN(n1015) );
  XOR2_X1 U1093 ( .A(G1986), .B(G24), .Z(n1011) );
  XNOR2_X1 U1094 ( .A(G1971), .B(G22), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(G23), .B(G1976), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(KEYINPUT58), .B(n1012), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(KEYINPUT126), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1101 ( .A(KEYINPUT61), .B(n1016), .Z(n1017) );
  NOR2_X1 U1102 ( .A1(G16), .A2(n1017), .ZN(n1018) );
  XOR2_X1 U1103 ( .A(KEYINPUT127), .B(n1018), .Z(n1019) );
  NOR2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(n1021), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
  INV_X1 U1107 ( .A(G303), .ZN(G166) );
endmodule

