//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n629, new_n630, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n808, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938;
  XNOR2_X1  g000(.A(KEYINPUT88), .B(KEYINPUT35), .ZN(new_n202));
  XOR2_X1   g001(.A(KEYINPUT74), .B(KEYINPUT22), .Z(new_n203));
  NAND2_X1  g002(.A1(G211gat), .A2(G218gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(new_n204), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n205), .A2(new_n206), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n206), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n204), .B(new_n209), .C1(new_n212), .C2(new_n203), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G141gat), .B(G148gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n216), .A2(KEYINPUT2), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n216), .ZN(new_n219));
  NOR2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  OR3_X1    g019(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT78), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT78), .B1(new_n219), .B2(new_n220), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n218), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n220), .B1(KEYINPUT77), .B2(new_n216), .ZN(new_n224));
  OAI221_X1 g023(.A(new_n224), .B1(KEYINPUT77), .B2(new_n216), .C1(new_n217), .C2(new_n215), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n223), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT29), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n214), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT83), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n211), .A2(KEYINPUT82), .A3(new_n213), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n228), .B1(new_n211), .B2(KEYINPUT82), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n226), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n223), .A2(new_n225), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT80), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n223), .A2(new_n225), .A3(KEYINPUT80), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n229), .A2(new_n230), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n231), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G228gat), .A2(G233gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G22gat), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT29), .B1(new_n211), .B2(new_n213), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n235), .B1(new_n246), .B2(KEYINPUT3), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n247), .A2(KEYINPUT84), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(KEYINPUT84), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n229), .A2(new_n243), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n244), .A2(new_n245), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n245), .B1(new_n244), .B2(new_n251), .ZN(new_n254));
  OAI21_X1  g053(.A(G78gat), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n244), .A2(new_n251), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G22gat), .ZN(new_n257));
  INV_X1    g056(.A(G78gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n258), .A3(new_n252), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT31), .B(G50gat), .ZN(new_n260));
  INV_X1    g059(.A(G106gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n255), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n262), .B1(new_n255), .B2(new_n259), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(G15gat), .B(G43gat), .Z(new_n267));
  XNOR2_X1  g066(.A(G71gat), .B(G99gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G183gat), .A2(G190gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT24), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(G183gat), .A2(G190gat), .ZN(new_n276));
  OR3_X1    g075(.A1(new_n275), .A2(KEYINPUT64), .A3(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT64), .B1(new_n275), .B2(new_n276), .ZN(new_n278));
  INV_X1    g077(.A(G169gat), .ZN(new_n279));
  INV_X1    g078(.A(G176gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n279), .A2(new_n280), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT23), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT65), .B(G169gat), .Z(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(KEYINPUT23), .A3(new_n280), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n277), .A2(new_n278), .A3(new_n284), .A4(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT25), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT66), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(KEYINPUT66), .A3(new_n288), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n281), .A2(new_n283), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(new_n288), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT67), .B(G183gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(G190gat), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n294), .B(new_n284), .C1(new_n296), .C2(new_n275), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n291), .A2(new_n292), .A3(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT27), .B(G183gat), .ZN(new_n299));
  INV_X1    g098(.A(G190gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(KEYINPUT28), .A3(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n301), .B(KEYINPUT69), .Z(new_n302));
  NOR2_X1   g101(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n303), .B1(new_n295), .B2(KEYINPUT27), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT68), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n305), .A2(new_n306), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n302), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n282), .B1(KEYINPUT26), .B2(new_n281), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n312), .A2(KEYINPUT70), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n281), .A2(KEYINPUT26), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(new_n312), .B2(KEYINPUT70), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n313), .A2(new_n315), .B1(G183gat), .B2(G190gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n298), .A2(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(KEYINPUT71), .B(G113gat), .Z(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G120gat), .ZN(new_n320));
  XOR2_X1   g119(.A(G127gat), .B(G134gat), .Z(new_n321));
  INV_X1    g120(.A(KEYINPUT72), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G113gat), .ZN(new_n324));
  INV_X1    g123(.A(G120gat), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT1), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G127gat), .B(G134gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT72), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n320), .A2(new_n323), .A3(new_n326), .A4(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n326), .B1(new_n324), .B2(new_n325), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n321), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(G227gat), .A2(G233gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n298), .A2(new_n317), .A3(new_n332), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT33), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n270), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n335), .B1(new_n334), .B2(new_n336), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT34), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI211_X1 g142(.A(KEYINPUT34), .B(new_n335), .C1(new_n334), .C2(new_n336), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n337), .A2(KEYINPUT32), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n341), .A2(new_n342), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n339), .B1(new_n349), .B2(new_n344), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n350), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n339), .A2(new_n349), .A3(new_n344), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n347), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n266), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n356), .B(KEYINPUT75), .Z(new_n357));
  AND3_X1   g156(.A1(new_n298), .A2(new_n317), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(KEYINPUT29), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n360), .B1(new_n298), .B2(new_n317), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n214), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n318), .A2(new_n359), .ZN(new_n363));
  INV_X1    g162(.A(new_n214), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n298), .A2(new_n317), .A3(new_n357), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G8gat), .B(G36gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n367), .B(new_n368), .Z(new_n369));
  NAND3_X1  g168(.A1(new_n362), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT76), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT30), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT30), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(KEYINPUT76), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n362), .A2(new_n366), .ZN(new_n375));
  INV_X1    g174(.A(new_n369), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n372), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n329), .A2(new_n223), .A3(new_n225), .A4(new_n331), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n333), .A2(new_n237), .A3(new_n238), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n382), .B1(new_n383), .B2(new_n381), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n332), .A2(new_n227), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n226), .B1(new_n223), .B2(new_n225), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT79), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n386), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT79), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n227), .A4(new_n332), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(KEYINPUT5), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n384), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT81), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n384), .A2(new_n391), .A3(new_n397), .A4(new_n394), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n393), .B1(new_n380), .B2(new_n381), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n391), .B(new_n399), .C1(new_n381), .C2(new_n383), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT5), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n332), .A2(new_n235), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n380), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n401), .B1(new_n403), .B2(new_n393), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n396), .A2(new_n398), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT0), .ZN(new_n407));
  XOR2_X1   g206(.A(G57gat), .B(G85gat), .Z(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT6), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n410), .B1(new_n409), .B2(new_n405), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n412));
  OR3_X1    g211(.A1(new_n405), .A2(new_n412), .A3(new_n409), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n379), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n202), .B1(new_n355), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n414), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(new_n378), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n346), .A2(new_n348), .A3(new_n350), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n348), .B1(new_n346), .B2(new_n350), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT35), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(KEYINPUT88), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n418), .A2(new_n421), .A3(new_n266), .A4(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n405), .A2(new_n409), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n392), .B1(new_n384), .B2(new_n391), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n402), .A2(new_n392), .A3(new_n380), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT39), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT86), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n409), .B1(new_n430), .B2(KEYINPUT40), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT39), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n431), .B1(new_n426), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(KEYINPUT85), .A2(KEYINPUT40), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(KEYINPUT86), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n429), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n429), .B2(new_n433), .ZN(new_n437));
  NOR3_X1   g236(.A1(new_n425), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n378), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n376), .B1(new_n375), .B2(KEYINPUT37), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n363), .A2(KEYINPUT87), .A3(new_n364), .A4(new_n365), .ZN(new_n442));
  OAI211_X1 g241(.A(KEYINPUT37), .B(new_n442), .C1(new_n375), .C2(KEYINPUT87), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT38), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  AND2_X1   g244(.A1(new_n375), .A2(KEYINPUT37), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT38), .B1(new_n446), .B2(new_n440), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n411), .A2(new_n413), .A3(new_n370), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n439), .B(new_n266), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n265), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n263), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(new_n417), .B2(new_n378), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT36), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT73), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n455), .A2(KEYINPUT73), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n456), .B(new_n457), .C1(new_n419), .C2(new_n420), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n354), .A2(KEYINPUT73), .A3(new_n455), .A4(new_n351), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n416), .B(new_n424), .C1(new_n454), .C2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G15gat), .B(G22gat), .ZN(new_n462));
  INV_X1    g261(.A(G1gat), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(KEYINPUT16), .A3(new_n463), .ZN(new_n464));
  OAI221_X1 g263(.A(new_n464), .B1(KEYINPUT91), .B2(G8gat), .C1(new_n463), .C2(new_n462), .ZN(new_n465));
  NAND2_X1  g264(.A1(KEYINPUT91), .A2(G8gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(G29gat), .A2(G36gat), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT14), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(G29gat), .A2(G36gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT89), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT15), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n471), .A2(KEYINPUT15), .A3(new_n473), .ZN(new_n477));
  XNOR2_X1  g276(.A(G43gat), .B(G50gat), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  OR2_X1    g278(.A1(new_n477), .A2(new_n478), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT17), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT90), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT17), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n484), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  AOI211_X1 g285(.A(KEYINPUT90), .B(KEYINPUT17), .C1(new_n479), .C2(new_n480), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n468), .B(new_n483), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G229gat), .A2(G233gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n467), .A2(new_n481), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT18), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n488), .A2(KEYINPUT18), .A3(new_n489), .A4(new_n490), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n467), .B(new_n481), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n489), .B(KEYINPUT13), .Z(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n493), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G113gat), .B(G141gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(G197gat), .ZN(new_n500));
  XOR2_X1   g299(.A(KEYINPUT11), .B(G169gat), .Z(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(KEYINPUT12), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n493), .A2(new_n503), .A3(new_n494), .A4(new_n497), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n461), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(G71gat), .A2(G78gat), .ZN(new_n509));
  INV_X1    g308(.A(G71gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n510), .A2(new_n258), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT92), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G57gat), .B(G64gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n513), .A2(KEYINPUT9), .ZN(new_n516));
  OAI221_X1 g315(.A(new_n514), .B1(new_n513), .B2(new_n512), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT95), .ZN(new_n518));
  INV_X1    g317(.A(G57gat), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT93), .B1(new_n519), .B2(G64gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n521));
  INV_X1    g320(.A(G64gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n522), .A3(G57gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(G64gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT94), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n520), .A2(new_n523), .A3(KEYINPUT94), .A4(new_n524), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n511), .B1(KEYINPUT9), .B2(new_n509), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n518), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  AOI211_X1 g331(.A(KEYINPUT95), .B(new_n530), .C1(new_n527), .C2(new_n528), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n517), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(KEYINPUT21), .ZN(new_n536));
  NAND2_X1  g335(.A1(G231gat), .A2(G233gat), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(G127gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n535), .A2(KEYINPUT21), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n468), .ZN(new_n543));
  INV_X1    g342(.A(G127gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n538), .A2(new_n544), .A3(new_n539), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n541), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n543), .B1(new_n541), .B2(new_n545), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n549));
  INV_X1    g348(.A(G155gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G183gat), .B(G211gat), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n551), .B(new_n552), .Z(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  OR3_X1    g353(.A1(new_n547), .A2(new_n548), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n554), .B1(new_n547), .B2(new_n548), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G190gat), .B(G218gat), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G85gat), .A2(G92gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT7), .ZN(new_n561));
  NAND2_X1  g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562));
  INV_X1    g361(.A(G85gat), .ZN(new_n563));
  INV_X1    g362(.A(G92gat), .ZN(new_n564));
  AOI22_X1  g363(.A1(KEYINPUT8), .A2(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G99gat), .B(G106gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n483), .B(new_n569), .C1(new_n486), .C2(new_n487), .ZN(new_n570));
  NAND2_X1  g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n481), .A2(new_n568), .B1(KEYINPUT41), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n559), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n570), .A2(new_n559), .A3(new_n573), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n572), .A2(KEYINPUT41), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT96), .ZN(new_n579));
  XOR2_X1   g378(.A(G134gat), .B(G162gat), .Z(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n581), .B1(new_n574), .B2(KEYINPUT97), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n575), .A2(KEYINPUT97), .A3(new_n576), .A4(new_n581), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n534), .A2(new_n569), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT10), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n568), .B(new_n517), .C1(new_n532), .C2(new_n533), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n535), .A2(KEYINPUT10), .A3(new_n568), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n586), .B1(new_n588), .B2(new_n590), .ZN(new_n594));
  XNOR2_X1  g393(.A(G120gat), .B(G148gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(G176gat), .B(G204gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NOR3_X1   g397(.A1(new_n593), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n586), .B(KEYINPUT98), .Z(new_n601));
  AOI21_X1  g400(.A(new_n601), .B1(new_n591), .B2(new_n592), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n598), .B1(new_n602), .B2(new_n594), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n557), .A2(new_n585), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n508), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(new_n414), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(new_n463), .ZN(G1324gat));
  OAI21_X1  g409(.A(G8gat), .B1(new_n608), .B2(new_n379), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT42), .ZN(new_n612));
  INV_X1    g411(.A(new_n608), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT16), .B(G8gat), .Z(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(new_n378), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n616), .A3(new_n612), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n616), .B1(new_n615), .B2(new_n612), .ZN(new_n619));
  OAI221_X1 g418(.A(new_n611), .B1(new_n612), .B2(new_n615), .C1(new_n618), .C2(new_n619), .ZN(G1325gat));
  NAND3_X1  g419(.A1(new_n613), .A2(G15gat), .A3(new_n460), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n508), .A2(new_n421), .A3(new_n607), .ZN(new_n622));
  INV_X1    g421(.A(G15gat), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n622), .A2(KEYINPUT100), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT100), .B1(new_n622), .B2(new_n623), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT101), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(G1326gat));
  NOR2_X1   g427(.A1(new_n608), .A2(new_n266), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT43), .B(G22gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(G1327gat));
  NOR3_X1   g430(.A1(new_n557), .A2(new_n585), .A3(new_n604), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n508), .A2(new_n632), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n633), .A2(G29gat), .A3(new_n414), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(KEYINPUT45), .Z(new_n635));
  AND2_X1   g434(.A1(new_n583), .A2(new_n584), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n637));
  AND3_X1   g436(.A1(new_n461), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT103), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n640), .A2(KEYINPUT44), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n641), .B1(new_n461), .B2(new_n636), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n555), .A2(KEYINPUT102), .A3(new_n556), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT102), .B1(new_n555), .B2(new_n556), .ZN(new_n646));
  INV_X1    g445(.A(new_n507), .ZN(new_n647));
  NOR4_X1   g446(.A1(new_n645), .A2(new_n646), .A3(new_n647), .A4(new_n604), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(KEYINPUT104), .B1(new_n649), .B2(new_n414), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(G29gat), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n649), .A2(KEYINPUT104), .A3(new_n414), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n635), .B1(new_n651), .B2(new_n652), .ZN(G1328gat));
  NOR3_X1   g452(.A1(new_n633), .A2(G36gat), .A3(new_n379), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT46), .ZN(new_n655));
  OAI21_X1  g454(.A(G36gat), .B1(new_n649), .B2(new_n379), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(G1329gat));
  INV_X1    g456(.A(new_n421), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n633), .A2(G43gat), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n460), .A3(new_n648), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n659), .B1(new_n660), .B2(G43gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT47), .ZN(G1330gat));
  OAI211_X1 g461(.A(new_n452), .B(new_n648), .C1(new_n638), .C2(new_n642), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT105), .B1(new_n663), .B2(G50gat), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT48), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n633), .A2(G50gat), .A3(new_n266), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n667), .B1(G50gat), .B2(new_n663), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n666), .B(new_n668), .ZN(G1331gat));
  INV_X1    g468(.A(new_n557), .ZN(new_n670));
  NOR4_X1   g469(.A1(new_n670), .A2(new_n507), .A3(new_n636), .A4(new_n605), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n461), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(new_n414), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(new_n519), .ZN(G1332gat));
  NOR2_X1   g473(.A1(new_n672), .A2(new_n379), .ZN(new_n675));
  NOR2_X1   g474(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n676));
  AND2_X1   g475(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(new_n675), .B2(new_n676), .ZN(G1333gat));
  AND2_X1   g478(.A1(new_n461), .A2(new_n671), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n510), .B1(new_n680), .B2(new_n460), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(KEYINPUT106), .A3(new_n421), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n683), .B1(new_n672), .B2(new_n658), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n681), .B1(new_n685), .B2(new_n510), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1334gat));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n266), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(new_n258), .ZN(G1335gat));
  NOR2_X1   g489(.A1(new_n557), .A2(new_n507), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n604), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n692), .B1(new_n639), .B2(new_n643), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G85gat), .B1(new_n694), .B2(new_n414), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n461), .A2(new_n636), .A3(new_n691), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT51), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n461), .A2(KEYINPUT51), .A3(new_n636), .A4(new_n691), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n417), .A2(new_n563), .A3(new_n604), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n695), .B1(new_n701), .B2(new_n702), .ZN(G1336gat));
  INV_X1    g502(.A(new_n692), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n378), .B(new_n704), .C1(new_n638), .C2(new_n642), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n564), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n696), .A2(KEYINPUT108), .A3(KEYINPUT51), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT51), .B1(new_n696), .B2(KEYINPUT108), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n379), .A2(G92gat), .A3(new_n605), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT52), .B1(new_n707), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G92gat), .B1(new_n706), .B2(KEYINPUT110), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n705), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT109), .B1(new_n701), .B2(new_n711), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT52), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n700), .A2(new_n720), .A3(new_n710), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n713), .B1(new_n717), .B2(new_n722), .ZN(G1337gat));
  INV_X1    g522(.A(G99gat), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n724), .B1(new_n693), .B2(new_n460), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n421), .A2(new_n724), .A3(new_n604), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n701), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n728));
  OR3_X1    g527(.A1(new_n725), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n725), .B2(new_n727), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(G1338gat));
  NOR3_X1   g530(.A1(new_n266), .A2(G106gat), .A3(new_n605), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT53), .B1(new_n700), .B2(new_n732), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n452), .B(new_n704), .C1(new_n638), .C2(new_n642), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G106gat), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT53), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n696), .A2(KEYINPUT108), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n697), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n696), .A2(KEYINPUT108), .A3(KEYINPUT51), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n739), .A2(new_n740), .A3(new_n732), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n737), .B1(new_n735), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT112), .B1(new_n736), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n733), .A2(new_n735), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n708), .A2(new_n709), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n746), .A2(new_n732), .B1(G106gat), .B2(new_n734), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n744), .B(new_n745), .C1(new_n747), .C2(new_n737), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n743), .A2(new_n748), .ZN(G1339gat));
  NOR2_X1   g548(.A1(new_n414), .A2(new_n378), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT115), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n645), .A2(new_n646), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n591), .A2(new_n592), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n586), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n591), .A2(new_n592), .A3(new_n601), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(KEYINPUT54), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT54), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n597), .B1(new_n602), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n756), .A2(KEYINPUT55), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT113), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n756), .A2(new_n758), .A3(new_n761), .A4(KEYINPUT55), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT55), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n591), .A2(new_n592), .A3(new_n601), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n764), .A2(new_n593), .A3(new_n757), .ZN(new_n765));
  INV_X1    g564(.A(new_n601), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n753), .A2(new_n757), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n598), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n763), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n760), .A2(new_n600), .A3(new_n762), .A4(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n758), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n599), .B1(new_n773), .B2(new_n763), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n774), .A2(new_n760), .A3(KEYINPUT114), .A4(new_n762), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n772), .A2(new_n507), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n489), .B1(new_n488), .B2(new_n490), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n495), .A2(new_n496), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n502), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n604), .A2(new_n506), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n636), .B1(new_n776), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n506), .A2(new_n779), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n585), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n772), .A2(new_n775), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n752), .B1(new_n781), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n606), .A2(new_n507), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n751), .B1(new_n789), .B2(new_n266), .ZN(new_n790));
  AOI211_X1 g589(.A(KEYINPUT115), .B(new_n452), .C1(new_n786), .C2(new_n788), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n421), .B(new_n750), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(G113gat), .B1(new_n792), .B2(new_n647), .ZN(new_n793));
  INV_X1    g592(.A(new_n355), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n789), .A2(new_n417), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT116), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n414), .B1(new_n786), .B2(new_n788), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(new_n798), .A3(new_n794), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n378), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n647), .A2(new_n319), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n801), .B(KEYINPUT117), .Z(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n793), .A2(new_n803), .ZN(G1340gat));
  OAI21_X1  g603(.A(G120gat), .B1(new_n792), .B2(new_n605), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n604), .A2(new_n325), .ZN(new_n806));
  XOR2_X1   g605(.A(new_n806), .B(KEYINPUT118), .Z(new_n807));
  NAND2_X1  g606(.A1(new_n800), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(G1341gat));
  NAND3_X1  g608(.A1(new_n800), .A2(new_n544), .A3(new_n557), .ZN(new_n810));
  OAI21_X1  g609(.A(G127gat), .B1(new_n792), .B2(new_n752), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(G1342gat));
  NOR2_X1   g611(.A1(new_n585), .A2(G134gat), .ZN(new_n813));
  AND4_X1   g612(.A1(new_n798), .A2(new_n789), .A3(new_n417), .A4(new_n794), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n798), .B1(new_n797), .B2(new_n794), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n379), .B(new_n813), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT56), .ZN(new_n817));
  OAI21_X1  g616(.A(G134gat), .B1(new_n792), .B2(new_n585), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n796), .A2(new_n799), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n819), .A2(new_n820), .A3(new_n379), .A4(new_n813), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n817), .A2(new_n818), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT119), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n817), .A2(new_n818), .A3(new_n821), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(G1343gat));
  INV_X1    g625(.A(G141gat), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n460), .A2(new_n378), .A3(new_n266), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n797), .A2(new_n827), .A3(new_n507), .A4(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n507), .A2(new_n774), .A3(new_n762), .A4(new_n760), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n780), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT120), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n830), .A2(new_n833), .A3(new_n780), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n585), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n784), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n787), .B1(new_n836), .B2(new_n670), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT57), .B1(new_n837), .B2(new_n266), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n266), .B1(new_n786), .B2(new_n788), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n460), .A2(new_n414), .A3(new_n378), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n647), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n829), .B1(new_n844), .B2(new_n827), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT58), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n847), .B(new_n829), .C1(new_n844), .C2(new_n827), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1344gat));
  NOR2_X1   g648(.A1(new_n605), .A2(G148gat), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n797), .A2(new_n828), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n789), .A2(new_n452), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n636), .A2(new_n762), .A3(new_n774), .A4(new_n760), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n782), .B1(new_n854), .B2(KEYINPUT121), .ZN(new_n855));
  OR3_X1    g654(.A1(new_n770), .A2(KEYINPUT121), .A3(new_n585), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n834), .A2(new_n585), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n833), .B1(new_n830), .B2(new_n780), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n670), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n788), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n266), .A2(KEYINPUT57), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n853), .A2(KEYINPUT57), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n604), .A3(new_n842), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n852), .B1(new_n865), .B2(G148gat), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n852), .A2(G148gat), .ZN(new_n867));
  INV_X1    g666(.A(new_n843), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n868), .B2(new_n604), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n851), .B1(new_n866), .B2(new_n869), .ZN(G1345gat));
  OAI21_X1  g669(.A(G155gat), .B1(new_n843), .B2(new_n752), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n797), .A2(new_n550), .A3(new_n557), .A4(new_n828), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(G1346gat));
  OAI21_X1  g672(.A(G162gat), .B1(new_n843), .B2(new_n585), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n585), .A2(G162gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n797), .A2(new_n828), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1347gat));
  NOR2_X1   g676(.A1(new_n417), .A2(new_n379), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n421), .B(new_n878), .C1(new_n790), .C2(new_n791), .ZN(new_n879));
  OAI21_X1  g678(.A(G169gat), .B1(new_n879), .B2(new_n647), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n417), .B1(new_n786), .B2(new_n788), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n881), .A2(new_n378), .A3(new_n794), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n507), .A3(new_n285), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT122), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n880), .A2(new_n886), .A3(new_n883), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(G1348gat));
  OAI21_X1  g687(.A(G176gat), .B1(new_n879), .B2(new_n605), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n882), .A2(new_n280), .A3(new_n604), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n890), .B1(new_n889), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(G1349gat));
  OAI21_X1  g693(.A(new_n295), .B1(new_n879), .B2(new_n752), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n882), .A2(new_n299), .A3(new_n557), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT60), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT60), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n895), .A2(new_n896), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(G1350gat));
  NAND3_X1  g700(.A1(new_n882), .A2(new_n300), .A3(new_n636), .ZN(new_n902));
  XOR2_X1   g701(.A(new_n902), .B(KEYINPUT124), .Z(new_n903));
  OAI21_X1  g702(.A(G190gat), .B1(new_n879), .B2(new_n585), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(G1351gat));
  XNOR2_X1  g707(.A(KEYINPUT125), .B(G197gat), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n460), .A2(new_n379), .A3(new_n266), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n881), .A2(new_n507), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n557), .B1(new_n835), .B2(new_n857), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n863), .B1(new_n912), .B2(new_n787), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n460), .A2(new_n417), .A3(new_n379), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n913), .B(new_n914), .C1(new_n839), .C2(new_n840), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n915), .A2(new_n647), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n911), .B1(new_n916), .B2(new_n909), .ZN(G1352gat));
  NAND3_X1  g716(.A1(new_n864), .A2(new_n604), .A3(new_n914), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G204gat), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n605), .A2(G204gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n881), .A2(new_n910), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT62), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n921), .A2(KEYINPUT62), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n919), .A2(new_n922), .A3(new_n923), .ZN(G1353gat));
  NAND4_X1  g723(.A1(new_n881), .A2(new_n207), .A3(new_n557), .A4(new_n910), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n915), .A2(new_n670), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n207), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT126), .B1(new_n915), .B2(new_n670), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT63), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n864), .A2(new_n927), .A3(new_n557), .A4(new_n914), .ZN(new_n931));
  AND4_X1   g730(.A1(KEYINPUT63), .A2(new_n931), .A3(new_n929), .A4(G211gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n925), .B1(new_n930), .B2(new_n932), .ZN(G1354gat));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n585), .B1(new_n915), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n935), .B1(new_n934), .B2(new_n915), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(G218gat), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n881), .A2(new_n208), .A3(new_n636), .A4(new_n910), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1355gat));
endmodule


