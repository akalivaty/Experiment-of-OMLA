

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U556 ( .A1(G651), .A2(n627), .ZN(n652) );
  OR2_X1 U557 ( .A1(n692), .A2(n982), .ZN(n691) );
  BUF_X1 U558 ( .A(n720), .Z(n730) );
  INV_X1 U559 ( .A(G168), .ZN(n724) );
  XNOR2_X1 U560 ( .A(n711), .B(n710), .ZN(n717) );
  XNOR2_X1 U561 ( .A(KEYINPUT100), .B(KEYINPUT32), .ZN(n741) );
  OR2_X1 U562 ( .A1(n798), .A2(n687), .ZN(n720) );
  XNOR2_X1 U563 ( .A(KEYINPUT95), .B(n719), .ZN(n769) );
  NOR2_X1 U564 ( .A1(G164), .A2(G1384), .ZN(n799) );
  NOR2_X2 U565 ( .A1(G2105), .A2(n540), .ZN(n888) );
  NOR2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n536) );
  NOR2_X1 U567 ( .A1(n814), .A2(n813), .ZN(n816) );
  XOR2_X1 U568 ( .A(n522), .B(KEYINPUT1), .Z(n648) );
  OR2_X1 U569 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U570 ( .A1(n546), .A2(n545), .ZN(G160) );
  INV_X1 U571 ( .A(G651), .ZN(n529) );
  NOR2_X1 U572 ( .A1(n529), .A2(G543), .ZN(n522) );
  NAND2_X1 U573 ( .A1(n648), .A2(G63), .ZN(n523) );
  XNOR2_X1 U574 ( .A(KEYINPUT73), .B(n523), .ZN(n526) );
  XOR2_X1 U575 ( .A(KEYINPUT0), .B(G543), .Z(n627) );
  NAND2_X1 U576 ( .A1(n652), .A2(G51), .ZN(n524) );
  XOR2_X1 U577 ( .A(KEYINPUT74), .B(n524), .Z(n525) );
  NOR2_X1 U578 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U579 ( .A(n527), .B(KEYINPUT6), .ZN(n534) );
  NOR2_X1 U580 ( .A1(G651), .A2(G543), .ZN(n643) );
  NAND2_X1 U581 ( .A1(n643), .A2(G89), .ZN(n528) );
  XNOR2_X1 U582 ( .A(n528), .B(KEYINPUT4), .ZN(n531) );
  NOR2_X1 U583 ( .A1(n627), .A2(n529), .ZN(n644) );
  NAND2_X1 U584 ( .A1(G76), .A2(n644), .ZN(n530) );
  NAND2_X1 U585 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U586 ( .A(KEYINPUT5), .B(n532), .ZN(n533) );
  NAND2_X1 U587 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U588 ( .A(n535), .B(KEYINPUT7), .ZN(G168) );
  AND2_X1 U589 ( .A1(G2104), .A2(G2105), .ZN(n893) );
  NAND2_X1 U590 ( .A1(n893), .A2(G113), .ZN(n538) );
  XOR2_X2 U591 ( .A(KEYINPUT17), .B(n536), .Z(n889) );
  NAND2_X1 U592 ( .A1(n889), .A2(G137), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n538), .A2(n537), .ZN(n546) );
  INV_X1 U594 ( .A(G2104), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n888), .A2(G101), .ZN(n539) );
  XOR2_X1 U596 ( .A(KEYINPUT23), .B(n539), .Z(n542) );
  AND2_X1 U597 ( .A1(n540), .A2(G2105), .ZN(n892) );
  NAND2_X1 U598 ( .A1(n892), .A2(G125), .ZN(n541) );
  NAND2_X1 U599 ( .A1(n542), .A2(n541), .ZN(n544) );
  INV_X1 U600 ( .A(KEYINPUT65), .ZN(n543) );
  XNOR2_X1 U601 ( .A(n544), .B(n543), .ZN(n545) );
  NAND2_X1 U602 ( .A1(G78), .A2(n644), .ZN(n548) );
  NAND2_X1 U603 ( .A1(G53), .A2(n652), .ZN(n547) );
  NAND2_X1 U604 ( .A1(n548), .A2(n547), .ZN(n552) );
  NAND2_X1 U605 ( .A1(G91), .A2(n643), .ZN(n550) );
  NAND2_X1 U606 ( .A1(G65), .A2(n648), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U608 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U609 ( .A(n553), .B(KEYINPUT69), .Z(n706) );
  INV_X1 U610 ( .A(n706), .ZN(G299) );
  NAND2_X1 U611 ( .A1(G126), .A2(n892), .ZN(n555) );
  NAND2_X1 U612 ( .A1(G138), .A2(n889), .ZN(n554) );
  NAND2_X1 U613 ( .A1(n555), .A2(n554), .ZN(n559) );
  NAND2_X1 U614 ( .A1(G102), .A2(n888), .ZN(n557) );
  NAND2_X1 U615 ( .A1(G114), .A2(n893), .ZN(n556) );
  NAND2_X1 U616 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U617 ( .A(KEYINPUT89), .B(n560), .ZN(G164) );
  NAND2_X1 U618 ( .A1(G64), .A2(n648), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G52), .A2(n652), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n562), .A2(n561), .ZN(n567) );
  NAND2_X1 U621 ( .A1(G90), .A2(n643), .ZN(n564) );
  NAND2_X1 U622 ( .A1(G77), .A2(n644), .ZN(n563) );
  NAND2_X1 U623 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U624 ( .A(KEYINPUT9), .B(n565), .Z(n566) );
  NOR2_X1 U625 ( .A1(n567), .A2(n566), .ZN(G171) );
  INV_X1 U626 ( .A(G132), .ZN(G219) );
  INV_X1 U627 ( .A(G82), .ZN(G220) );
  INV_X1 U628 ( .A(G57), .ZN(G237) );
  INV_X1 U629 ( .A(G120), .ZN(G236) );
  XNOR2_X1 U630 ( .A(G168), .B(KEYINPUT8), .ZN(n568) );
  XNOR2_X1 U631 ( .A(n568), .B(KEYINPUT75), .ZN(G286) );
  NAND2_X1 U632 ( .A1(G94), .A2(G452), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT68), .B(n569), .Z(G173) );
  NAND2_X1 U634 ( .A1(G7), .A2(G661), .ZN(n570) );
  XOR2_X1 U635 ( .A(n570), .B(KEYINPUT10), .Z(n833) );
  NAND2_X1 U636 ( .A1(n833), .A2(G567), .ZN(n571) );
  XOR2_X1 U637 ( .A(KEYINPUT11), .B(n571), .Z(G234) );
  NAND2_X1 U638 ( .A1(G56), .A2(n648), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT14), .B(n572), .Z(n578) );
  NAND2_X1 U640 ( .A1(n643), .A2(G81), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n573), .B(KEYINPUT12), .ZN(n575) );
  NAND2_X1 U642 ( .A1(G68), .A2(n644), .ZN(n574) );
  NAND2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U644 ( .A(KEYINPUT13), .B(n576), .Z(n577) );
  NOR2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n652), .A2(G43), .ZN(n579) );
  NAND2_X1 U647 ( .A1(n580), .A2(n579), .ZN(n977) );
  INV_X1 U648 ( .A(G860), .ZN(n611) );
  OR2_X1 U649 ( .A1(n977), .A2(n611), .ZN(G153) );
  XOR2_X1 U650 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  INV_X1 U651 ( .A(G868), .ZN(n592) );
  NOR2_X1 U652 ( .A1(G301), .A2(n592), .ZN(n591) );
  NAND2_X1 U653 ( .A1(G79), .A2(n644), .ZN(n582) );
  NAND2_X1 U654 ( .A1(G54), .A2(n652), .ZN(n581) );
  NAND2_X1 U655 ( .A1(n582), .A2(n581), .ZN(n587) );
  NAND2_X1 U656 ( .A1(G92), .A2(n643), .ZN(n584) );
  NAND2_X1 U657 ( .A1(G66), .A2(n648), .ZN(n583) );
  NAND2_X1 U658 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U659 ( .A(n585), .B(KEYINPUT71), .Z(n586) );
  NOR2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U661 ( .A(KEYINPUT15), .B(n588), .Z(n589) );
  XNOR2_X2 U662 ( .A(KEYINPUT72), .B(n589), .ZN(n982) );
  AND2_X1 U663 ( .A1(n982), .A2(n592), .ZN(n590) );
  NOR2_X1 U664 ( .A1(n591), .A2(n590), .ZN(G284) );
  NOR2_X1 U665 ( .A1(G868), .A2(G299), .ZN(n594) );
  NOR2_X1 U666 ( .A1(G286), .A2(n592), .ZN(n593) );
  NOR2_X1 U667 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U668 ( .A(KEYINPUT76), .B(n595), .ZN(G297) );
  NAND2_X1 U669 ( .A1(n611), .A2(G559), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n596), .A2(n982), .ZN(n597) );
  XNOR2_X1 U671 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U672 ( .A1(G868), .A2(n977), .ZN(n600) );
  NAND2_X1 U673 ( .A1(n982), .A2(G868), .ZN(n598) );
  NOR2_X1 U674 ( .A1(G559), .A2(n598), .ZN(n599) );
  NOR2_X1 U675 ( .A1(n600), .A2(n599), .ZN(G282) );
  NAND2_X1 U676 ( .A1(G123), .A2(n892), .ZN(n601) );
  XNOR2_X1 U677 ( .A(n601), .B(KEYINPUT18), .ZN(n603) );
  NAND2_X1 U678 ( .A1(n888), .A2(G99), .ZN(n602) );
  NAND2_X1 U679 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U680 ( .A1(G135), .A2(n889), .ZN(n605) );
  NAND2_X1 U681 ( .A1(G111), .A2(n893), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U683 ( .A1(n607), .A2(n606), .ZN(n930) );
  XOR2_X1 U684 ( .A(G2096), .B(n930), .Z(n608) );
  NOR2_X1 U685 ( .A1(G2100), .A2(n608), .ZN(n609) );
  XNOR2_X1 U686 ( .A(KEYINPUT77), .B(n609), .ZN(G156) );
  NAND2_X1 U687 ( .A1(n982), .A2(G559), .ZN(n610) );
  XOR2_X1 U688 ( .A(n977), .B(n610), .Z(n663) );
  NAND2_X1 U689 ( .A1(n611), .A2(n663), .ZN(n619) );
  NAND2_X1 U690 ( .A1(G93), .A2(n643), .ZN(n613) );
  NAND2_X1 U691 ( .A1(G80), .A2(n644), .ZN(n612) );
  NAND2_X1 U692 ( .A1(n613), .A2(n612), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n648), .A2(G67), .ZN(n614) );
  XNOR2_X1 U694 ( .A(n614), .B(KEYINPUT78), .ZN(n616) );
  NAND2_X1 U695 ( .A1(G55), .A2(n652), .ZN(n615) );
  NAND2_X1 U696 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n666) );
  XOR2_X1 U698 ( .A(n619), .B(n666), .Z(G145) );
  NAND2_X1 U699 ( .A1(G88), .A2(n643), .ZN(n621) );
  NAND2_X1 U700 ( .A1(G62), .A2(n648), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U702 ( .A1(G50), .A2(n652), .ZN(n622) );
  XNOR2_X1 U703 ( .A(KEYINPUT81), .B(n622), .ZN(n623) );
  NOR2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n644), .A2(G75), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(G303) );
  NAND2_X1 U707 ( .A1(n627), .A2(G87), .ZN(n629) );
  NAND2_X1 U708 ( .A1(G651), .A2(G74), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U710 ( .A1(G49), .A2(n652), .ZN(n630) );
  XNOR2_X1 U711 ( .A(KEYINPUT79), .B(n630), .ZN(n631) );
  NOR2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n634) );
  INV_X1 U713 ( .A(n648), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n634), .A2(n633), .ZN(G288) );
  NAND2_X1 U715 ( .A1(G86), .A2(n643), .ZN(n636) );
  NAND2_X1 U716 ( .A1(G61), .A2(n648), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U718 ( .A(KEYINPUT80), .B(n637), .ZN(n640) );
  NAND2_X1 U719 ( .A1(G73), .A2(n644), .ZN(n638) );
  XOR2_X1 U720 ( .A(KEYINPUT2), .B(n638), .Z(n639) );
  NOR2_X1 U721 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U722 ( .A1(n652), .A2(G48), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(G305) );
  NAND2_X1 U724 ( .A1(G85), .A2(n643), .ZN(n646) );
  NAND2_X1 U725 ( .A1(G72), .A2(n644), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U727 ( .A(KEYINPUT66), .B(n647), .ZN(n651) );
  NAND2_X1 U728 ( .A1(G60), .A2(n648), .ZN(n649) );
  XNOR2_X1 U729 ( .A(KEYINPUT67), .B(n649), .ZN(n650) );
  NOR2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n654) );
  NAND2_X1 U731 ( .A1(n652), .A2(G47), .ZN(n653) );
  NAND2_X1 U732 ( .A1(n654), .A2(n653), .ZN(G290) );
  XOR2_X1 U733 ( .A(G303), .B(n666), .Z(n661) );
  XNOR2_X1 U734 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n656) );
  XNOR2_X1 U735 ( .A(G288), .B(KEYINPUT84), .ZN(n655) );
  XNOR2_X1 U736 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U737 ( .A(KEYINPUT19), .B(n657), .ZN(n659) );
  XOR2_X1 U738 ( .A(G305), .B(G299), .Z(n658) );
  XNOR2_X1 U739 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U740 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U741 ( .A(n662), .B(G290), .ZN(n905) );
  XNOR2_X1 U742 ( .A(n905), .B(n663), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n664), .A2(G868), .ZN(n665) );
  XOR2_X1 U744 ( .A(KEYINPUT85), .B(n665), .Z(n668) );
  OR2_X1 U745 ( .A1(n666), .A2(G868), .ZN(n667) );
  NAND2_X1 U746 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XOR2_X1 U748 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U749 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U750 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U751 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U753 ( .A1(G236), .A2(G237), .ZN(n673) );
  NAND2_X1 U754 ( .A1(G69), .A2(n673), .ZN(n674) );
  XNOR2_X1 U755 ( .A(KEYINPUT87), .B(n674), .ZN(n675) );
  NAND2_X1 U756 ( .A1(n675), .A2(G108), .ZN(n676) );
  XNOR2_X1 U757 ( .A(KEYINPUT88), .B(n676), .ZN(n838) );
  NAND2_X1 U758 ( .A1(G567), .A2(n838), .ZN(n682) );
  NOR2_X1 U759 ( .A1(G220), .A2(G219), .ZN(n677) );
  XOR2_X1 U760 ( .A(KEYINPUT22), .B(n677), .Z(n678) );
  NOR2_X1 U761 ( .A1(G218), .A2(n678), .ZN(n679) );
  NAND2_X1 U762 ( .A1(G96), .A2(n679), .ZN(n837) );
  NAND2_X1 U763 ( .A1(G2106), .A2(n837), .ZN(n680) );
  XNOR2_X1 U764 ( .A(KEYINPUT86), .B(n680), .ZN(n681) );
  NAND2_X1 U765 ( .A1(n682), .A2(n681), .ZN(n860) );
  NAND2_X1 U766 ( .A1(G483), .A2(G661), .ZN(n683) );
  NOR2_X1 U767 ( .A1(n860), .A2(n683), .ZN(n836) );
  NAND2_X1 U768 ( .A1(n836), .A2(G36), .ZN(G176) );
  NAND2_X1 U769 ( .A1(G160), .A2(G40), .ZN(n798) );
  INV_X1 U770 ( .A(n799), .ZN(n687) );
  NOR2_X1 U771 ( .A1(n798), .A2(n687), .ZN(n693) );
  AND2_X1 U772 ( .A1(n693), .A2(G1996), .ZN(n686) );
  XOR2_X1 U773 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n685) );
  XNOR2_X1 U774 ( .A(n686), .B(n685), .ZN(n689) );
  NAND2_X1 U775 ( .A1(n730), .A2(G1341), .ZN(n688) );
  NAND2_X1 U776 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U777 ( .A1(n977), .A2(n690), .ZN(n692) );
  XNOR2_X1 U778 ( .A(n691), .B(KEYINPUT98), .ZN(n699) );
  NAND2_X1 U779 ( .A1(n692), .A2(n982), .ZN(n697) );
  NOR2_X1 U780 ( .A1(G2067), .A2(n730), .ZN(n695) );
  BUF_X1 U781 ( .A(n693), .Z(n713) );
  NOR2_X1 U782 ( .A1(n713), .A2(G1348), .ZN(n694) );
  NOR2_X1 U783 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U784 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U785 ( .A1(n699), .A2(n698), .ZN(n704) );
  NAND2_X1 U786 ( .A1(n713), .A2(G2072), .ZN(n700) );
  XNOR2_X1 U787 ( .A(n700), .B(KEYINPUT27), .ZN(n702) );
  AND2_X1 U788 ( .A1(G1956), .A2(n730), .ZN(n701) );
  NOR2_X1 U789 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U790 ( .A1(n706), .A2(n705), .ZN(n703) );
  NAND2_X1 U791 ( .A1(n704), .A2(n703), .ZN(n709) );
  NOR2_X1 U792 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U793 ( .A(n707), .B(KEYINPUT28), .Z(n708) );
  NAND2_X1 U794 ( .A1(n709), .A2(n708), .ZN(n711) );
  INV_X1 U795 ( .A(KEYINPUT29), .ZN(n710) );
  XOR2_X1 U796 ( .A(G2078), .B(KEYINPUT25), .Z(n712) );
  XNOR2_X1 U797 ( .A(KEYINPUT97), .B(n712), .ZN(n952) );
  NOR2_X1 U798 ( .A1(n730), .A2(n952), .ZN(n715) );
  INV_X1 U799 ( .A(G1961), .ZN(n976) );
  NOR2_X1 U800 ( .A1(n713), .A2(n976), .ZN(n714) );
  NOR2_X1 U801 ( .A1(n715), .A2(n714), .ZN(n726) );
  NAND2_X1 U802 ( .A1(G171), .A2(n726), .ZN(n716) );
  NAND2_X1 U803 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U804 ( .A(KEYINPUT99), .B(n718), .ZN(n746) );
  AND2_X1 U805 ( .A1(n720), .A2(G8), .ZN(n719) );
  NOR2_X1 U806 ( .A1(G1966), .A2(n769), .ZN(n748) );
  NOR2_X1 U807 ( .A1(n720), .A2(G2084), .ZN(n721) );
  XOR2_X1 U808 ( .A(n721), .B(KEYINPUT96), .Z(n743) );
  NAND2_X1 U809 ( .A1(G8), .A2(n743), .ZN(n722) );
  NOR2_X1 U810 ( .A1(n748), .A2(n722), .ZN(n723) );
  XNOR2_X1 U811 ( .A(n723), .B(KEYINPUT30), .ZN(n725) );
  AND2_X1 U812 ( .A1(n725), .A2(n724), .ZN(n728) );
  NOR2_X1 U813 ( .A1(G171), .A2(n726), .ZN(n727) );
  NOR2_X1 U814 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U815 ( .A(n729), .B(KEYINPUT31), .ZN(n745) );
  INV_X1 U816 ( .A(G8), .ZN(n735) );
  NOR2_X1 U817 ( .A1(G1971), .A2(n769), .ZN(n732) );
  NOR2_X1 U818 ( .A1(G2090), .A2(n730), .ZN(n731) );
  NOR2_X1 U819 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U820 ( .A1(n733), .A2(G303), .ZN(n734) );
  NOR2_X1 U821 ( .A1(n735), .A2(n734), .ZN(n738) );
  OR2_X2 U822 ( .A1(n745), .A2(n738), .ZN(n736) );
  OR2_X2 U823 ( .A1(n746), .A2(n736), .ZN(n740) );
  AND2_X1 U824 ( .A1(G286), .A2(G8), .ZN(n737) );
  OR2_X1 U825 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U826 ( .A1(n740), .A2(n739), .ZN(n742) );
  XNOR2_X1 U827 ( .A(n742), .B(n741), .ZN(n752) );
  INV_X1 U828 ( .A(n743), .ZN(n744) );
  NAND2_X1 U829 ( .A1(n744), .A2(G8), .ZN(n750) );
  NOR2_X1 U830 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U831 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U832 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U833 ( .A1(n752), .A2(n751), .ZN(n768) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n774) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n753) );
  NOR2_X1 U836 ( .A1(n774), .A2(n753), .ZN(n986) );
  XOR2_X1 U837 ( .A(n986), .B(KEYINPUT101), .Z(n754) );
  NAND2_X1 U838 ( .A1(n768), .A2(n754), .ZN(n755) );
  XNOR2_X1 U839 ( .A(n755), .B(KEYINPUT102), .ZN(n760) );
  XOR2_X1 U840 ( .A(G1981), .B(G305), .Z(n994) );
  INV_X1 U841 ( .A(n994), .ZN(n756) );
  NOR2_X1 U842 ( .A1(KEYINPUT33), .A2(n756), .ZN(n758) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n985) );
  INV_X1 U844 ( .A(n769), .ZN(n773) );
  AND2_X1 U845 ( .A1(n985), .A2(n773), .ZN(n757) );
  AND2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n759) );
  AND2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n765) );
  INV_X1 U848 ( .A(n773), .ZN(n763) );
  NOR2_X1 U849 ( .A1(G1981), .A2(G305), .ZN(n761) );
  XOR2_X1 U850 ( .A(n761), .B(KEYINPUT24), .Z(n762) );
  NOR2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n780) );
  NOR2_X1 U853 ( .A1(G2090), .A2(G303), .ZN(n766) );
  NAND2_X1 U854 ( .A1(G8), .A2(n766), .ZN(n767) );
  NAND2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n770) );
  NAND2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n772) );
  INV_X1 U857 ( .A(KEYINPUT103), .ZN(n771) );
  XNOR2_X1 U858 ( .A(n772), .B(n771), .ZN(n778) );
  NAND2_X1 U859 ( .A1(n774), .A2(n773), .ZN(n776) );
  AND2_X1 U860 ( .A1(n994), .A2(KEYINPUT33), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n776), .A2(n775), .ZN(n777) );
  AND2_X1 U862 ( .A1(n778), .A2(n777), .ZN(n779) );
  AND2_X1 U863 ( .A1(n780), .A2(n779), .ZN(n814) );
  NAND2_X1 U864 ( .A1(n889), .A2(G131), .ZN(n783) );
  NAND2_X1 U865 ( .A1(G107), .A2(n893), .ZN(n781) );
  XOR2_X1 U866 ( .A(KEYINPUT93), .B(n781), .Z(n782) );
  NAND2_X1 U867 ( .A1(n783), .A2(n782), .ZN(n787) );
  NAND2_X1 U868 ( .A1(G95), .A2(n888), .ZN(n785) );
  NAND2_X1 U869 ( .A1(G119), .A2(n892), .ZN(n784) );
  NAND2_X1 U870 ( .A1(n785), .A2(n784), .ZN(n786) );
  OR2_X1 U871 ( .A1(n787), .A2(n786), .ZN(n882) );
  AND2_X1 U872 ( .A1(n882), .A2(G1991), .ZN(n797) );
  NAND2_X1 U873 ( .A1(G105), .A2(n888), .ZN(n788) );
  XNOR2_X1 U874 ( .A(n788), .B(KEYINPUT38), .ZN(n795) );
  NAND2_X1 U875 ( .A1(G129), .A2(n892), .ZN(n790) );
  NAND2_X1 U876 ( .A1(G141), .A2(n889), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U878 ( .A1(n893), .A2(G117), .ZN(n791) );
  XOR2_X1 U879 ( .A(KEYINPUT94), .B(n791), .Z(n792) );
  NOR2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U881 ( .A1(n795), .A2(n794), .ZN(n883) );
  AND2_X1 U882 ( .A1(n883), .A2(G1996), .ZN(n796) );
  NOR2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n937) );
  INV_X1 U884 ( .A(n937), .ZN(n800) );
  NOR2_X1 U885 ( .A1(n799), .A2(n798), .ZN(n828) );
  NAND2_X1 U886 ( .A1(n800), .A2(n828), .ZN(n817) );
  NAND2_X1 U887 ( .A1(G128), .A2(n892), .ZN(n802) );
  NAND2_X1 U888 ( .A1(G116), .A2(n893), .ZN(n801) );
  NAND2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U890 ( .A(KEYINPUT35), .B(n803), .Z(n811) );
  NAND2_X1 U891 ( .A1(n889), .A2(G140), .ZN(n804) );
  XNOR2_X1 U892 ( .A(KEYINPUT91), .B(n804), .ZN(n807) );
  NAND2_X1 U893 ( .A1(n888), .A2(G104), .ZN(n805) );
  XOR2_X1 U894 ( .A(n805), .B(KEYINPUT90), .Z(n806) );
  NOR2_X1 U895 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U896 ( .A(KEYINPUT34), .B(n808), .Z(n809) );
  XNOR2_X1 U897 ( .A(n809), .B(KEYINPUT92), .ZN(n810) );
  NOR2_X1 U898 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U899 ( .A(KEYINPUT36), .B(n812), .ZN(n902) );
  XNOR2_X1 U900 ( .A(G2067), .B(KEYINPUT37), .ZN(n825) );
  NOR2_X1 U901 ( .A1(n902), .A2(n825), .ZN(n946) );
  NAND2_X1 U902 ( .A1(n828), .A2(n946), .ZN(n823) );
  NAND2_X1 U903 ( .A1(n817), .A2(n823), .ZN(n813) );
  XNOR2_X1 U904 ( .A(G1986), .B(G290), .ZN(n979) );
  NAND2_X1 U905 ( .A1(n979), .A2(n828), .ZN(n815) );
  NAND2_X1 U906 ( .A1(n816), .A2(n815), .ZN(n831) );
  NOR2_X1 U907 ( .A1(G1996), .A2(n883), .ZN(n939) );
  INV_X1 U908 ( .A(n817), .ZN(n820) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U910 ( .A1(G1991), .A2(n882), .ZN(n931) );
  NOR2_X1 U911 ( .A1(n818), .A2(n931), .ZN(n819) );
  NOR2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U913 ( .A1(n939), .A2(n821), .ZN(n822) );
  XNOR2_X1 U914 ( .A(KEYINPUT39), .B(n822), .ZN(n824) );
  NAND2_X1 U915 ( .A1(n824), .A2(n823), .ZN(n826) );
  NAND2_X1 U916 ( .A1(n902), .A2(n825), .ZN(n943) );
  NAND2_X1 U917 ( .A1(n826), .A2(n943), .ZN(n827) );
  NAND2_X1 U918 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U919 ( .A(KEYINPUT104), .B(n829), .ZN(n830) );
  NAND2_X1 U920 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U921 ( .A(KEYINPUT40), .B(n832), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n833), .ZN(G217) );
  INV_X1 U923 ( .A(n833), .ZN(G223) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U925 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U927 ( .A1(n836), .A2(n835), .ZN(G188) );
  XNOR2_X1 U928 ( .A(G96), .B(KEYINPUT105), .ZN(G221) );
  INV_X1 U930 ( .A(G108), .ZN(G238) );
  NOR2_X1 U931 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  XOR2_X1 U933 ( .A(n976), .B(G2474), .Z(n849) );
  XOR2_X1 U934 ( .A(G1986), .B(G1966), .Z(n840) );
  XNOR2_X1 U935 ( .A(G1981), .B(G1956), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n840), .B(n839), .ZN(n845) );
  INV_X1 U937 ( .A(G1996), .ZN(n841) );
  XNOR2_X1 U938 ( .A(G1991), .B(n841), .ZN(n843) );
  XNOR2_X1 U939 ( .A(G1976), .B(G1971), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U941 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U942 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n846) );
  XNOR2_X1 U943 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U944 ( .A(n849), .B(n848), .ZN(G229) );
  XOR2_X1 U945 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n851) );
  XNOR2_X1 U946 ( .A(G2678), .B(KEYINPUT43), .ZN(n850) );
  XNOR2_X1 U947 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U948 ( .A(KEYINPUT42), .B(G2072), .Z(n853) );
  XNOR2_X1 U949 ( .A(G2090), .B(G2067), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U951 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U952 ( .A(G2096), .B(G2100), .ZN(n856) );
  XNOR2_X1 U953 ( .A(n857), .B(n856), .ZN(n859) );
  XOR2_X1 U954 ( .A(G2078), .B(G2084), .Z(n858) );
  XNOR2_X1 U955 ( .A(n859), .B(n858), .ZN(G227) );
  INV_X1 U956 ( .A(n860), .ZN(G319) );
  NAND2_X1 U957 ( .A1(G100), .A2(n888), .ZN(n862) );
  NAND2_X1 U958 ( .A1(G112), .A2(n893), .ZN(n861) );
  NAND2_X1 U959 ( .A1(n862), .A2(n861), .ZN(n868) );
  NAND2_X1 U960 ( .A1(n892), .A2(G124), .ZN(n863) );
  XNOR2_X1 U961 ( .A(n863), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U962 ( .A1(G136), .A2(n889), .ZN(n864) );
  NAND2_X1 U963 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U964 ( .A(KEYINPUT109), .B(n866), .Z(n867) );
  NOR2_X1 U965 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U966 ( .A(KEYINPUT110), .B(n869), .ZN(G162) );
  NAND2_X1 U967 ( .A1(G130), .A2(n892), .ZN(n871) );
  NAND2_X1 U968 ( .A1(G118), .A2(n893), .ZN(n870) );
  NAND2_X1 U969 ( .A1(n871), .A2(n870), .ZN(n876) );
  NAND2_X1 U970 ( .A1(G106), .A2(n888), .ZN(n873) );
  NAND2_X1 U971 ( .A1(G142), .A2(n889), .ZN(n872) );
  NAND2_X1 U972 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U973 ( .A(KEYINPUT45), .B(n874), .Z(n875) );
  NOR2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U975 ( .A(G160), .B(n877), .Z(n878) );
  XNOR2_X1 U976 ( .A(G162), .B(n878), .ZN(n887) );
  XOR2_X1 U977 ( .A(KEYINPUT111), .B(KEYINPUT46), .Z(n880) );
  XNOR2_X1 U978 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n879) );
  XNOR2_X1 U979 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U980 ( .A(n881), .B(n930), .Z(n885) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U983 ( .A(n887), .B(n886), .Z(n901) );
  NAND2_X1 U984 ( .A1(G103), .A2(n888), .ZN(n891) );
  NAND2_X1 U985 ( .A1(G139), .A2(n889), .ZN(n890) );
  NAND2_X1 U986 ( .A1(n891), .A2(n890), .ZN(n899) );
  NAND2_X1 U987 ( .A1(G127), .A2(n892), .ZN(n895) );
  NAND2_X1 U988 ( .A1(G115), .A2(n893), .ZN(n894) );
  NAND2_X1 U989 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U990 ( .A(KEYINPUT112), .B(n896), .Z(n897) );
  XNOR2_X1 U991 ( .A(KEYINPUT47), .B(n897), .ZN(n898) );
  NOR2_X1 U992 ( .A1(n899), .A2(n898), .ZN(n926) );
  XNOR2_X1 U993 ( .A(G164), .B(n926), .ZN(n900) );
  XNOR2_X1 U994 ( .A(n901), .B(n900), .ZN(n903) );
  XNOR2_X1 U995 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U996 ( .A1(G37), .A2(n904), .ZN(G395) );
  XNOR2_X1 U997 ( .A(n977), .B(n905), .ZN(n907) );
  XNOR2_X1 U998 ( .A(G286), .B(G171), .ZN(n906) );
  XNOR2_X1 U999 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1000 ( .A(n908), .B(n982), .ZN(n909) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n909), .ZN(G397) );
  NOR2_X1 U1002 ( .A1(G229), .A2(G227), .ZN(n911) );
  XNOR2_X1 U1003 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n910) );
  XNOR2_X1 U1004 ( .A(n911), .B(n910), .ZN(n922) );
  XOR2_X1 U1005 ( .A(G2451), .B(G2430), .Z(n913) );
  XNOR2_X1 U1006 ( .A(G2438), .B(G2443), .ZN(n912) );
  XNOR2_X1 U1007 ( .A(n913), .B(n912), .ZN(n919) );
  XOR2_X1 U1008 ( .A(G2435), .B(G2454), .Z(n915) );
  XNOR2_X1 U1009 ( .A(G1348), .B(G1341), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n915), .B(n914), .ZN(n917) );
  XOR2_X1 U1011 ( .A(G2446), .B(G2427), .Z(n916) );
  XNOR2_X1 U1012 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1013 ( .A(n919), .B(n918), .Z(n920) );
  NAND2_X1 U1014 ( .A1(G14), .A2(n920), .ZN(n925) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n925), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1018 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G303), .ZN(G166) );
  INV_X1 U1021 ( .A(G69), .ZN(G235) );
  INV_X1 U1022 ( .A(n925), .ZN(G401) );
  XOR2_X1 U1023 ( .A(G2072), .B(n926), .Z(n928) );
  XOR2_X1 U1024 ( .A(G164), .B(G2078), .Z(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(KEYINPUT50), .B(n929), .ZN(n933) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n935) );
  XOR2_X1 U1029 ( .A(G160), .B(G2084), .Z(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n942) );
  XOR2_X1 U1032 ( .A(G2090), .B(G162), .Z(n938) );
  NOR2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1034 ( .A(n940), .B(KEYINPUT51), .ZN(n941) );
  NOR2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n944) );
  NAND2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1037 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1038 ( .A(KEYINPUT52), .B(n947), .ZN(n949) );
  INV_X1 U1039 ( .A(KEYINPUT55), .ZN(n948) );
  NAND2_X1 U1040 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1041 ( .A1(n950), .A2(G29), .ZN(n1035) );
  XOR2_X1 U1042 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n951) );
  XNOR2_X1 U1043 ( .A(KEYINPUT53), .B(n951), .ZN(n964) );
  XOR2_X1 U1044 ( .A(G1996), .B(G32), .Z(n954) );
  XNOR2_X1 U1045 ( .A(n952), .B(G27), .ZN(n953) );
  NAND2_X1 U1046 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1047 ( .A(KEYINPUT115), .B(n955), .ZN(n959) );
  XNOR2_X1 U1048 ( .A(G2067), .B(G26), .ZN(n957) );
  XNOR2_X1 U1049 ( .A(G1991), .B(G25), .ZN(n956) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n962) );
  XOR2_X1 U1052 ( .A(G2072), .B(G33), .Z(n960) );
  NAND2_X1 U1053 ( .A1(G28), .A2(n960), .ZN(n961) );
  NOR2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(n964), .B(n963), .ZN(n966) );
  XNOR2_X1 U1056 ( .A(G35), .B(G2090), .ZN(n965) );
  NOR2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1058 ( .A(KEYINPUT118), .B(n967), .ZN(n971) );
  XNOR2_X1 U1059 ( .A(KEYINPUT54), .B(G34), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(n968), .B(KEYINPUT119), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(G2084), .B(n969), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1063 ( .A(KEYINPUT55), .B(n972), .Z(n974) );
  INV_X1 U1064 ( .A(G29), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1066 ( .A1(G11), .A2(n975), .ZN(n1033) );
  INV_X1 U1067 ( .A(G16), .ZN(n1029) );
  XOR2_X1 U1068 ( .A(n1029), .B(KEYINPUT56), .Z(n1001) );
  XOR2_X1 U1069 ( .A(G171), .B(n976), .Z(n981) );
  XNOR2_X1 U1070 ( .A(G1341), .B(n977), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n984) );
  XOR2_X1 U1073 ( .A(G1348), .B(n982), .Z(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n999) );
  NAND2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n990) );
  XOR2_X1 U1076 ( .A(G1956), .B(G299), .Z(n988) );
  NAND2_X1 U1077 ( .A1(G1971), .A2(G303), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1080 ( .A(n991), .B(KEYINPUT121), .ZN(n997) );
  XNOR2_X1 U1081 ( .A(G168), .B(G1966), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(n992), .B(KEYINPUT120), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1084 ( .A(KEYINPUT57), .B(n995), .Z(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1031) );
  XOR2_X1 U1088 ( .A(KEYINPUT58), .B(KEYINPUT127), .Z(n1008) );
  XNOR2_X1 U1089 ( .A(G1976), .B(G23), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(G1986), .B(G24), .ZN(n1002) );
  NOR2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1006) );
  XOR2_X1 U1092 ( .A(G1971), .B(KEYINPUT126), .Z(n1004) );
  XNOR2_X1 U1093 ( .A(G22), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(n1008), .B(n1007), .ZN(n1026) );
  XOR2_X1 U1096 ( .A(G5), .B(G1961), .Z(n1024) );
  XNOR2_X1 U1097 ( .A(G1956), .B(G20), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(G1981), .B(G6), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(n1009), .B(KEYINPUT122), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(G19), .B(G1341), .ZN(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(KEYINPUT123), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1104 ( .A(KEYINPUT124), .B(n1015), .Z(n1019) );
  XNOR2_X1 U1105 ( .A(KEYINPUT59), .B(G4), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(n1016), .B(KEYINPUT125), .ZN(n1017) );
  XNOR2_X1 U1107 ( .A(G1348), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1109 ( .A(KEYINPUT60), .B(n1020), .Z(n1022) );
  XNOR2_X1 U1110 ( .A(G1966), .B(G21), .ZN(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1114 ( .A(KEYINPUT61), .B(n1027), .ZN(n1028) );
  NAND2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1117 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1118 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1036), .ZN(G150) );
  INV_X1 U1120 ( .A(G150), .ZN(G311) );
endmodule

