//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1220, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT64), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n208), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XNOR2_X1  g0033(.A(G50), .B(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G58), .B(G77), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XOR2_X1   g0036(.A(G97), .B(G107), .Z(new_n237));
  XNOR2_X1  g0037(.A(G87), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  INV_X1    g0040(.A(G179), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT66), .B(G1698), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT3), .B(G33), .ZN(new_n243));
  NAND3_X1  g0043(.A1(new_n242), .A2(new_n243), .A3(G232), .ZN(new_n244));
  INV_X1    g0044(.A(G107), .ZN(new_n245));
  INV_X1    g0045(.A(G238), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n243), .A2(G1698), .ZN(new_n247));
  OAI221_X1 g0047(.A(new_n244), .B1(new_n245), .B2(new_n243), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G1), .A3(G13), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n250), .A2(G274), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT65), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n205), .B(KEYINPUT65), .C1(G41), .C2(G45), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n250), .A2(new_n254), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n253), .A2(new_n258), .B1(new_n259), .B2(G244), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT68), .ZN(new_n261));
  AND3_X1   g0061(.A1(new_n252), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n261), .B1(new_n252), .B2(new_n260), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n241), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n214), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT8), .B(G58), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G77), .ZN(new_n270));
  OAI22_X1  g0070(.A1(new_n267), .A2(new_n269), .B1(new_n206), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT15), .B(G87), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n206), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n266), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(new_n266), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n270), .B1(new_n205), .B2(G20), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n278), .A2(new_n279), .B1(new_n270), .B2(new_n277), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n264), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n262), .A2(new_n263), .ZN(new_n283));
  INV_X1    g0083(.A(G169), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n281), .B1(new_n283), .B2(G200), .ZN(new_n287));
  OAI21_X1  g0087(.A(G190), .B1(new_n262), .B2(new_n263), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n290), .A2(KEYINPUT69), .ZN(new_n291));
  INV_X1    g0091(.A(G68), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT70), .B1(new_n277), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT12), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(G20), .ZN(new_n295));
  INV_X1    g0095(.A(G50), .ZN(new_n296));
  OAI221_X1 g0096(.A(new_n295), .B1(new_n273), .B2(new_n270), .C1(new_n269), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n266), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT11), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n205), .A2(G20), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n278), .A2(G68), .A3(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(new_n298), .B2(new_n299), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT13), .ZN(new_n307));
  INV_X1    g0107(.A(G33), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT3), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT3), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  AND2_X1   g0112(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n313));
  NOR2_X1   g0113(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n314));
  OAI21_X1  g0114(.A(G226), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G232), .A2(G1698), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n312), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G33), .A2(G97), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n251), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n253), .A2(new_n258), .B1(new_n259), .B2(G238), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n307), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n320), .A2(new_n321), .A3(new_n307), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(G179), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n324), .ZN(new_n326));
  OAI21_X1  g0126(.A(G169), .B1(new_n326), .B2(new_n322), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n325), .B1(new_n327), .B2(KEYINPUT14), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT14), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n323), .A2(new_n324), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(G169), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n306), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n323), .A2(G190), .A3(new_n324), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n326), .A2(new_n322), .ZN(new_n334));
  INV_X1    g0134(.A(G200), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n333), .B(new_n305), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n266), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n276), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n302), .A2(G50), .ZN(new_n340));
  OAI22_X1  g0140(.A1(new_n339), .A2(new_n340), .B1(G50), .B2(new_n276), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT67), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G150), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n267), .A2(new_n273), .B1(new_n344), .B2(new_n269), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n206), .B1(new_n201), .B2(new_n296), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n266), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n242), .A2(new_n243), .A3(G222), .ZN(new_n349));
  INV_X1    g0149(.A(G223), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n349), .B1(new_n270), .B2(new_n243), .C1(new_n350), .C2(new_n247), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n251), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n253), .A2(new_n258), .B1(new_n259), .B2(G226), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n348), .B1(new_n354), .B2(G169), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n354), .A2(new_n241), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n348), .B(KEYINPUT9), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n354), .A2(new_n335), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(G190), .B2(new_n354), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT10), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT10), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n358), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n357), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n290), .A2(KEYINPUT69), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n291), .A2(new_n337), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n267), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n302), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n369), .A2(new_n339), .B1(new_n276), .B2(new_n368), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G58), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(new_n292), .ZN(new_n373));
  OAI21_X1  g0173(.A(G20), .B1(new_n373), .B2(new_n201), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n268), .A2(G159), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT7), .B1(new_n312), .B2(new_n206), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT7), .ZN(new_n378));
  AOI211_X1 g0178(.A(new_n378), .B(G20), .C1(new_n309), .C2(new_n311), .ZN(new_n379));
  OAI21_X1  g0179(.A(G68), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT71), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n376), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n378), .B1(new_n243), .B2(G20), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n312), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n292), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT71), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT16), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n376), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n380), .A2(KEYINPUT16), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n266), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n371), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n309), .A2(new_n311), .A3(G226), .A4(G1698), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n309), .B(new_n311), .C1(new_n313), .C2(new_n314), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n392), .B(new_n393), .C1(new_n394), .C2(new_n350), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n251), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n253), .A2(new_n258), .B1(new_n259), .B2(G232), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n396), .A2(new_n241), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(G169), .B1(new_n396), .B2(new_n397), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT72), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT72), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n396), .A2(new_n397), .A3(new_n241), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n396), .A2(new_n397), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n401), .B(new_n402), .C1(new_n403), .C2(G169), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n391), .A2(KEYINPUT18), .A3(new_n400), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT73), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n404), .A2(new_n400), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT73), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n407), .A2(new_n408), .A3(KEYINPUT18), .A4(new_n391), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT18), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n404), .A2(new_n400), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT16), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n380), .A2(new_n381), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n388), .B1(new_n385), .B2(KEYINPUT71), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n385), .A2(new_n376), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n338), .B1(new_n416), .B2(KEYINPUT16), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n370), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n410), .B1(new_n411), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n406), .A2(new_n409), .A3(new_n419), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n396), .A2(G190), .A3(new_n397), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n335), .B1(new_n396), .B2(new_n397), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n423), .B(new_n371), .C1(new_n387), .C2(new_n390), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT17), .B1(new_n418), .B2(new_n423), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n420), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT21), .ZN(new_n430));
  INV_X1    g0230(.A(G257), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT80), .B1(new_n394), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT80), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n242), .A2(new_n243), .A3(new_n433), .A4(G257), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n309), .A2(new_n311), .A3(G264), .A4(G1698), .ZN(new_n436));
  INV_X1    g0236(.A(G303), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n436), .B1(new_n437), .B2(new_n243), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n440), .A2(KEYINPUT81), .A3(new_n251), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT81), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n438), .B1(new_n432), .B2(new_n434), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n443), .B2(new_n250), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G1), .ZN(new_n446));
  AND2_X1   g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  NOR2_X1   g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(G270), .A3(new_n250), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT79), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT5), .B(G41), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n452), .A2(G274), .A3(new_n250), .A4(new_n446), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(new_n453), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT79), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n441), .A2(new_n444), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G116), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n277), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n308), .A2(G1), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n460), .B(KEYINPUT75), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(G116), .A3(new_n278), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G283), .ZN(new_n463));
  INV_X1    g0263(.A(G97), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n463), .B(new_n206), .C1(G33), .C2(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n465), .B(new_n266), .C1(new_n206), .C2(G116), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT20), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n466), .A2(new_n467), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n459), .B(new_n462), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G169), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n430), .B1(new_n457), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT83), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT83), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n474), .B(new_n430), .C1(new_n457), .C2(new_n471), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n456), .A2(new_n454), .ZN(new_n477));
  AOI21_X1  g0277(.A(KEYINPUT81), .B1(new_n440), .B2(new_n251), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n443), .A2(new_n442), .A3(new_n250), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n470), .B1(new_n480), .B2(G200), .ZN(new_n481));
  INV_X1    g0281(.A(G190), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(new_n480), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n480), .A2(KEYINPUT21), .A3(G169), .A4(new_n470), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n241), .B1(new_n456), .B2(new_n454), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n470), .B(new_n485), .C1(new_n478), .C2(new_n479), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n484), .A2(KEYINPUT82), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT82), .B1(new_n484), .B2(new_n486), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n476), .B(new_n483), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G87), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT78), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n490), .A2(KEYINPUT78), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n491), .A2(new_n492), .A3(new_n464), .A4(new_n245), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT19), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT77), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT77), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT19), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n318), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n493), .B1(new_n498), .B2(G20), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n495), .B(new_n497), .C1(new_n273), .C2(new_n464), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n309), .A2(new_n311), .A3(new_n206), .A4(G68), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n338), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n461), .A2(new_n278), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n490), .ZN(new_n506));
  INV_X1    g0306(.A(new_n272), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(new_n276), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n504), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT76), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n250), .A2(G274), .A3(new_n446), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n205), .A2(G45), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n250), .A2(G250), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n510), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n511), .A2(new_n513), .A3(new_n510), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G116), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n309), .A2(new_n311), .A3(G244), .A4(G1698), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n517), .B(new_n518), .C1(new_n394), .C2(new_n246), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n515), .A2(new_n516), .B1(new_n519), .B2(new_n251), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G190), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n251), .ZN(new_n522));
  INV_X1    g0322(.A(new_n516), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n522), .B1(new_n523), .B2(new_n514), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G200), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n509), .A2(new_n521), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n508), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n461), .A2(new_n278), .A3(new_n507), .ZN(new_n528));
  OR2_X1    g0328(.A1(new_n498), .A2(G20), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n502), .B1(new_n529), .B2(new_n493), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n527), .B(new_n528), .C1(new_n530), .C2(new_n338), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n522), .B(new_n241), .C1(new_n514), .C2(new_n523), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n531), .B(new_n532), .C1(G169), .C2(new_n520), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n277), .A2(new_n464), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n505), .B2(new_n464), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  XNOR2_X1  g0337(.A(G97), .B(G107), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT6), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n539), .A2(new_n464), .A3(G107), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n543), .A2(G20), .B1(G77), .B2(new_n268), .ZN(new_n544));
  OAI21_X1  g0344(.A(G107), .B1(new_n377), .B2(new_n379), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n338), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT74), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n541), .B1(new_n539), .B2(new_n538), .ZN(new_n549));
  OAI22_X1  g0349(.A1(new_n549), .A2(new_n206), .B1(new_n270), .B2(new_n269), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n245), .B1(new_n383), .B2(new_n384), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n266), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n552), .A2(KEYINPUT74), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n537), .B1(new_n548), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n449), .A2(G257), .A3(new_n250), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n453), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT4), .ZN(new_n557));
  INV_X1    g0357(.A(G244), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n557), .B1(new_n394), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n242), .A2(new_n243), .A3(KEYINPUT4), .A4(G244), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n243), .A2(G250), .A3(G1698), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n559), .A2(new_n463), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n556), .B1(new_n562), .B2(new_n251), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(G169), .ZN(new_n564));
  AOI211_X1 g0364(.A(G179), .B(new_n556), .C1(new_n562), .C2(new_n251), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n554), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n546), .A2(new_n547), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n552), .A2(KEYINPUT74), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n536), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n563), .A2(new_n482), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(G200), .B2(new_n563), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n534), .A2(new_n567), .A3(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(G250), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n394), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n309), .A2(new_n311), .A3(G257), .A4(G1698), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G294), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n251), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n449), .A2(G264), .A3(new_n250), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT88), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT88), .B1(new_n580), .B2(new_n581), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n453), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n335), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT87), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(KEYINPUT87), .B(new_n251), .C1(new_n576), .C2(new_n579), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n587), .A2(new_n453), .A3(new_n588), .A4(new_n581), .ZN(new_n589));
  OR2_X1    g0389(.A1(new_n589), .A2(G190), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  OR3_X1    g0391(.A1(new_n206), .A2(KEYINPUT23), .A3(G107), .ZN(new_n592));
  OAI21_X1  g0392(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT24), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n592), .B(new_n593), .C1(KEYINPUT86), .C2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n206), .A2(G33), .A3(G116), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT85), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  AND2_X1   g0399(.A1(KEYINPUT84), .A2(G87), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n243), .A2(new_n206), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT22), .ZN(new_n602));
  OR2_X1    g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n602), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n599), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n594), .A2(KEYINPUT86), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n266), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n505), .A2(new_n245), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT25), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n276), .B2(G107), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n277), .A2(KEYINPUT25), .A3(new_n245), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n591), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(G179), .B(new_n453), .C1(new_n582), .C2(new_n583), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n589), .A2(G169), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT89), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n609), .A2(new_n614), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n616), .A2(new_n617), .A3(KEYINPUT89), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n574), .A2(new_n615), .A3(new_n623), .ZN(new_n624));
  NOR4_X1   g0424(.A1(new_n367), .A2(new_n429), .A3(new_n489), .A4(new_n624), .ZN(G372));
  NOR2_X1   g0425(.A1(new_n367), .A2(new_n429), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT91), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n520), .A2(KEYINPUT90), .A3(G169), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT90), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n524), .B2(new_n284), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n532), .B(new_n531), .C1(new_n628), .C2(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n567), .A2(new_n573), .A3(new_n526), .A4(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n621), .B1(new_n590), .B2(new_n585), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n627), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n567), .A2(new_n573), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n631), .A2(new_n526), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n635), .A2(new_n636), .A3(KEYINPUT91), .A4(new_n615), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n484), .A2(new_n486), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n621), .A2(new_n618), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n476), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n634), .A2(new_n637), .A3(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n570), .A2(new_n565), .A3(new_n564), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n534), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT26), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n636), .A2(new_n646), .A3(new_n643), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n645), .A2(new_n647), .A3(new_n631), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n626), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n419), .A2(new_n405), .ZN(new_n651));
  INV_X1    g0451(.A(new_n332), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n282), .A2(new_n285), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n652), .B1(new_n653), .B2(new_n336), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n424), .A2(new_n425), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n418), .A2(KEYINPUT17), .A3(new_n423), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n651), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n364), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n363), .B1(new_n358), .B2(new_n360), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n357), .B1(new_n658), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n650), .A2(new_n663), .ZN(G369));
  NAND2_X1  g0464(.A1(new_n476), .A2(new_n639), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n470), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n489), .B2(new_n672), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT92), .Z(new_n675));
  NAND2_X1  g0475(.A1(new_n621), .A2(new_n671), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n623), .A2(new_n615), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n671), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n677), .B1(new_n623), .B2(new_n678), .ZN(new_n679));
  XOR2_X1   g0479(.A(new_n679), .B(KEYINPUT93), .Z(new_n680));
  NAND3_X1  g0480(.A1(new_n675), .A2(G330), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT94), .ZN(new_n682));
  INV_X1    g0482(.A(new_n488), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n484), .A2(KEYINPUT82), .A3(new_n486), .ZN(new_n684));
  AOI22_X1  g0484(.A1(new_n683), .A2(new_n684), .B1(new_n475), .B2(new_n473), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n671), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n621), .A2(new_n618), .A3(new_n678), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n682), .A2(new_n689), .ZN(G399));
  INV_X1    g0490(.A(new_n209), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G41), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n493), .A2(G116), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G1), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n212), .B2(new_n693), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT28), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n476), .B(new_n623), .C1(new_n487), .C2(new_n488), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(new_n615), .A3(new_n635), .A4(new_n636), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n631), .B1(new_n644), .B2(KEYINPUT26), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n646), .B1(new_n636), .B2(new_n643), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n671), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT29), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(G330), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n480), .A2(new_n241), .A3(new_n524), .ZN(new_n707));
  INV_X1    g0507(.A(new_n453), .ZN(new_n708));
  INV_X1    g0508(.A(new_n583), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT88), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT96), .B1(new_n711), .B2(new_n563), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT96), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n562), .A2(new_n251), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n584), .B(new_n713), .C1(new_n714), .C2(new_n556), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n707), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT95), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(KEYINPUT30), .ZN(new_n718));
  OAI22_X1  g0518(.A1(new_n478), .A2(new_n479), .B1(new_n582), .B2(new_n583), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n485), .A2(new_n563), .A3(new_n520), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n709), .A2(new_n710), .B1(new_n441), .B2(new_n444), .ZN(new_n722));
  INV_X1    g0522(.A(new_n720), .ZN(new_n723));
  INV_X1    g0523(.A(new_n718), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n671), .B1(new_n716), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT31), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI211_X1 g0529(.A(KEYINPUT31), .B(new_n671), .C1(new_n716), .C2(new_n726), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n624), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n733), .A2(new_n685), .A3(new_n483), .A4(new_n678), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n706), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n649), .A2(new_n704), .A3(new_n678), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n705), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n697), .B1(new_n738), .B2(G1), .ZN(G364));
  AND2_X1   g0539(.A1(new_n206), .A2(G13), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n205), .B1(new_n740), .B2(G45), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n693), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(new_n675), .B2(G330), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(G330), .B2(new_n675), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n214), .B1(G20), .B2(new_n284), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n209), .A2(new_n312), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n236), .A2(new_n445), .ZN(new_n752));
  XOR2_X1   g0552(.A(new_n752), .B(KEYINPUT97), .Z(new_n753));
  AOI211_X1 g0553(.A(new_n751), .B(new_n753), .C1(new_n445), .C2(new_n213), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n209), .A2(new_n243), .ZN(new_n755));
  INV_X1    g0555(.A(G355), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n755), .A2(new_n756), .B1(G116), .B2(new_n209), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n750), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n743), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n206), .A2(new_n241), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G190), .ZN(new_n762));
  INV_X1    g0562(.A(G317), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(KEYINPUT33), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n763), .A2(KEYINPUT33), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n762), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G294), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n482), .A2(G179), .A3(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n206), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n206), .A2(G179), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n766), .B1(new_n767), .B2(new_n769), .C1(new_n437), .C2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G190), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n243), .B1(new_n775), .B2(G329), .ZN(new_n776));
  INV_X1    g0576(.A(G311), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n760), .A2(new_n773), .ZN(new_n778));
  INV_X1    g0578(.A(G322), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n760), .A2(G190), .A3(new_n335), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n776), .B1(new_n777), .B2(new_n778), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n761), .A2(new_n482), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(KEYINPUT98), .B(G326), .Z(new_n784));
  NAND3_X1  g0584(.A1(new_n770), .A2(new_n482), .A3(G200), .ZN(new_n785));
  INV_X1    g0585(.A(G283), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n783), .A2(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n772), .A2(new_n781), .A3(new_n787), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n788), .A2(KEYINPUT99), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(KEYINPUT99), .ZN(new_n790));
  INV_X1    g0590(.A(new_n762), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT32), .ZN(new_n792));
  INV_X1    g0592(.A(G159), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n774), .A2(new_n793), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n791), .A2(new_n292), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(new_n792), .B2(new_n794), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n243), .B1(new_n780), .B2(new_n372), .ZN(new_n797));
  INV_X1    g0597(.A(new_n778), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(G77), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n771), .B1(new_n491), .B2(new_n492), .ZN(new_n800));
  INV_X1    g0600(.A(new_n769), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n800), .B1(G97), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n785), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n782), .A2(G50), .B1(new_n803), .B2(G107), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n796), .A2(new_n799), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n789), .A2(new_n790), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n759), .B1(new_n749), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n748), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n674), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n745), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G396));
  NAND2_X1  g0611(.A1(new_n649), .A2(new_n678), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n282), .A2(new_n285), .A3(new_n678), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n287), .A2(new_n288), .B1(new_n281), .B2(new_n671), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n653), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  AND3_X1   g0616(.A1(new_n282), .A2(new_n285), .A3(new_n678), .ZN(new_n817));
  INV_X1    g0617(.A(new_n814), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(new_n818), .B2(new_n286), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n649), .A2(new_n678), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n732), .A2(new_n734), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(G330), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n743), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n823), .B2(new_n821), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n749), .A2(new_n746), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n742), .B1(new_n270), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n749), .ZN(new_n828));
  INV_X1    g0628(.A(new_n780), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n829), .A2(G143), .B1(new_n798), .B2(G159), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n830), .B1(new_n791), .B2(new_n344), .C1(new_n831), .C2(new_n783), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT34), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n803), .A2(G68), .ZN(new_n835));
  INV_X1    g0635(.A(G132), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n835), .B(new_n243), .C1(new_n836), .C2(new_n774), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n769), .A2(new_n372), .B1(new_n771), .B2(new_n296), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n834), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n833), .B2(new_n832), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n786), .A2(new_n791), .B1(new_n783), .B2(new_n437), .ZN(new_n841));
  INV_X1    g0641(.A(new_n771), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(G107), .B2(new_n842), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n780), .A2(new_n767), .B1(new_n774), .B2(new_n777), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n243), .B(new_n844), .C1(G116), .C2(new_n798), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n785), .A2(new_n490), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G97), .B2(new_n801), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n843), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n840), .A2(new_n848), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n827), .B1(new_n828), .B2(new_n849), .C1(new_n819), .C2(new_n747), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n825), .A2(new_n850), .ZN(G384));
  OAI21_X1  g0651(.A(new_n412), .B1(new_n385), .B2(new_n376), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n370), .B1(new_n417), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n669), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n429), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n391), .B1(new_n407), .B2(new_n855), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n859), .A2(new_n860), .A3(new_n424), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n855), .B1(new_n404), .B2(new_n400), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n424), .B1(new_n862), .B2(new_n853), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n858), .A2(KEYINPUT38), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT101), .B1(new_n862), .B2(new_n418), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n867), .A2(new_n859), .A3(KEYINPUT37), .A4(new_n424), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(KEYINPUT37), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n424), .B1(new_n862), .B2(new_n418), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n657), .B1(new_n405), .B2(new_n419), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n418), .A2(new_n669), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n868), .B(new_n871), .C1(new_n872), .C2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n866), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n856), .B1(new_n420), .B2(new_n428), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n861), .A2(new_n864), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n876), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n878), .B1(new_n866), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT102), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n652), .A2(new_n678), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n858), .B2(new_n865), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n880), .A2(new_n881), .A3(new_n876), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT39), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT102), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n866), .A2(new_n877), .A3(new_n878), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n884), .A2(new_n886), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n651), .A2(new_n855), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n327), .A2(KEYINPUT14), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n330), .A2(new_n329), .A3(G169), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n336), .A2(new_n895), .A3(new_n325), .A4(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT100), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n305), .A2(new_n678), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n899), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n332), .A2(new_n336), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n898), .B1(new_n897), .B2(new_n899), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n820), .B2(new_n813), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n866), .A2(new_n882), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n894), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n893), .A2(KEYINPUT103), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT103), .B1(new_n893), .B2(new_n908), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n626), .B1(new_n705), .B2(new_n737), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n663), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT104), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n911), .B(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n428), .A2(new_n651), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n916), .A2(new_n873), .B1(new_n870), .B2(new_n869), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n917), .B2(new_n868), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(new_n888), .ZN(new_n919));
  INV_X1    g0719(.A(new_n905), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n489), .A2(new_n624), .A3(new_n671), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n920), .B(new_n819), .C1(new_n921), .C2(new_n731), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT40), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT40), .B1(new_n866), .B2(new_n882), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n819), .B1(new_n904), .B2(new_n903), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n732), .B2(new_n734), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n626), .A2(new_n822), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n706), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n929), .B2(new_n928), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n915), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n932), .A2(KEYINPUT105), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(KEYINPUT105), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n915), .A2(new_n931), .B1(new_n205), .B2(new_n740), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n543), .A2(KEYINPUT35), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n543), .A2(KEYINPUT35), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n937), .A2(G116), .A3(new_n215), .A4(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT36), .Z(new_n940));
  OR3_X1    g0740(.A1(new_n212), .A2(new_n270), .A3(new_n373), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n296), .A2(G68), .ZN(new_n942));
  AOI211_X1 g0742(.A(new_n205), .B(G13), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  OR3_X1    g0743(.A1(new_n936), .A2(new_n940), .A3(new_n943), .ZN(G367));
  OR2_X1    g0744(.A1(new_n509), .A2(new_n678), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n636), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT106), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(KEYINPUT106), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n947), .B(new_n948), .C1(new_n631), .C2(new_n945), .ZN(new_n949));
  XOR2_X1   g0749(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(KEYINPUT43), .B2(new_n949), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n635), .B1(new_n570), .B2(new_n678), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n567), .B1(new_n953), .B2(new_n623), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n678), .ZN(new_n955));
  INV_X1    g0755(.A(new_n687), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n643), .A2(new_n671), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n956), .A2(KEYINPUT42), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(KEYINPUT42), .B1(new_n956), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n955), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  MUX2_X1   g0761(.A(new_n951), .B(new_n952), .S(new_n961), .Z(new_n962));
  INV_X1    g0762(.A(new_n682), .ZN(new_n963));
  INV_X1    g0763(.A(new_n958), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n962), .B(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n692), .B(KEYINPUT41), .Z(new_n967));
  OAI211_X1 g0767(.A(new_n689), .B(new_n964), .C1(KEYINPUT108), .C2(KEYINPUT44), .ZN(new_n968));
  NAND2_X1  g0768(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n689), .A2(new_n964), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n682), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n970), .A2(new_n963), .A3(new_n972), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n680), .A2(new_n686), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n956), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n675), .A2(G330), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n974), .A2(new_n738), .A3(new_n975), .A4(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n967), .B1(new_n980), .B2(new_n738), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n741), .B(KEYINPUT109), .Z(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n966), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n750), .B1(new_n209), .B2(new_n272), .C1(new_n232), .C2(new_n751), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n743), .A2(new_n985), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n791), .A2(new_n793), .B1(new_n771), .B2(new_n372), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G68), .B2(new_n801), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n780), .A2(new_n344), .B1(new_n778), .B2(new_n296), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n312), .B(new_n989), .C1(G137), .C2(new_n775), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n782), .A2(G143), .B1(new_n803), .B2(G77), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n988), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n791), .A2(new_n767), .B1(new_n785), .B2(new_n464), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G311), .B2(new_n782), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n769), .A2(new_n245), .B1(new_n778), .B2(new_n786), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n995), .A2(KEYINPUT110), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(KEYINPUT110), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n842), .A2(KEYINPUT46), .A3(G116), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n243), .B1(new_n775), .B2(G317), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n829), .A2(G303), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT46), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n771), .B2(new_n458), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n992), .B1(new_n998), .B2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT47), .Z(new_n1006));
  OAI221_X1 g0806(.A(new_n986), .B1(new_n828), .B2(new_n1006), .C1(new_n949), .C2(new_n808), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n984), .A2(new_n1007), .ZN(G387));
  NOR2_X1   g0808(.A1(new_n979), .A2(new_n738), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n979), .A2(new_n738), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n692), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1009), .B1(new_n1011), .B2(KEYINPUT112), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(KEYINPUT112), .B2(new_n1011), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n979), .A2(new_n983), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n829), .A2(G317), .B1(new_n798), .B2(G303), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n791), .B2(new_n777), .C1(new_n779), .C2(new_n783), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT48), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n786), .B2(new_n769), .C1(new_n767), .C2(new_n771), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1021), .A2(KEYINPUT49), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n312), .B1(new_n785), .B2(new_n458), .C1(new_n774), .C2(new_n784), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(KEYINPUT49), .B2(new_n1021), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n778), .A2(new_n292), .B1(new_n774), .B2(new_n344), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n312), .B(new_n1026), .C1(G50), .C2(new_n829), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n842), .A2(G77), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n507), .A2(new_n801), .B1(new_n762), .B2(new_n368), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n782), .A2(G159), .B1(new_n803), .B2(G97), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n828), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n229), .A2(new_n445), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n1033), .A2(new_n751), .B1(new_n694), .B2(new_n755), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n267), .A2(G50), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n694), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1034), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(G107), .B2(new_n209), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n742), .B(new_n1032), .C1(new_n750), .C2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n680), .B2(new_n808), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1013), .A2(new_n1014), .A3(new_n1043), .ZN(G393));
  NAND2_X1  g0844(.A1(new_n974), .A2(new_n975), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n1010), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1046), .A2(new_n692), .A3(new_n980), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n974), .A2(new_n975), .A3(new_n983), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n750), .B1(new_n464), .B2(new_n209), .C1(new_n239), .C2(new_n751), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n743), .A2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT113), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n791), .A2(new_n296), .B1(new_n771), .B2(new_n292), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n846), .B(new_n1052), .C1(G77), .C2(new_n801), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n775), .A2(G143), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n312), .B1(new_n798), .B2(new_n368), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n783), .A2(new_n344), .B1(new_n793), .B2(new_n780), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT51), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G317), .A2(new_n782), .B1(new_n829), .B2(G311), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n791), .A2(new_n437), .B1(new_n785), .B2(new_n245), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n312), .B1(new_n774), .B2(new_n779), .C1(new_n767), .C2(new_n778), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n769), .A2(new_n458), .B1(new_n771), .B2(new_n786), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1056), .A2(new_n1058), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1051), .B1(new_n828), .B2(new_n1066), .C1(new_n958), .C2(new_n808), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1047), .A2(new_n1048), .A3(new_n1067), .ZN(G390));
  NAND3_X1  g0868(.A1(new_n735), .A2(new_n819), .A3(new_n920), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n820), .A2(new_n813), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n920), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n884), .A2(new_n892), .B1(new_n1072), .B2(new_n885), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n866), .A2(new_n877), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n653), .A2(new_n814), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n817), .B1(new_n703), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n885), .B(new_n1074), .C1(new_n1077), .C2(new_n905), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1070), .B1(new_n1073), .B2(new_n1079), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n879), .A2(new_n883), .A3(KEYINPUT102), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n890), .B1(new_n889), .B2(new_n891), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n1081), .A2(new_n1082), .B1(new_n886), .B2(new_n906), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1083), .A2(new_n1078), .A3(new_n1069), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n626), .A2(new_n735), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n912), .A2(new_n663), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n920), .B1(new_n735), .B2(new_n819), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1071), .B1(new_n1070), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1088), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(new_n1077), .A3(new_n1069), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1087), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1085), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1080), .A2(new_n1084), .A3(new_n1092), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(new_n692), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1080), .A2(new_n1084), .A3(new_n983), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n746), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n826), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n743), .B1(new_n368), .B2(new_n1099), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n245), .A2(new_n791), .B1(new_n783), .B2(new_n786), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G87), .B2(new_n842), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n801), .A2(G77), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n780), .A2(new_n458), .B1(new_n778), .B2(new_n464), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n243), .B(new_n1104), .C1(G294), .C2(new_n775), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1102), .A2(new_n835), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n842), .A2(G150), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT53), .ZN(new_n1108));
  INV_X1    g0908(.A(G125), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n243), .B1(new_n774), .B2(new_n1109), .C1(new_n780), .C2(new_n836), .ZN(new_n1110));
  INV_X1    g0910(.A(G128), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n783), .A2(new_n1111), .B1(new_n793), .B2(new_n769), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n785), .A2(new_n296), .ZN(new_n1113));
  OR4_X1    g0913(.A1(new_n1108), .A2(new_n1110), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT54), .B(G143), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n791), .A2(new_n831), .B1(new_n778), .B2(new_n1115), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT115), .Z(new_n1117));
  OAI21_X1  g0917(.A(new_n1106), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1100), .B1(new_n1118), .B2(new_n749), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1098), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1096), .A2(new_n1097), .A3(new_n1120), .ZN(G378));
  NAND2_X1  g0921(.A1(new_n348), .A2(new_n855), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n661), .B2(new_n357), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n365), .A2(new_n1122), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n928), .B2(G330), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n706), .B(new_n1129), .C1(new_n923), .C2(new_n927), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n893), .A2(new_n908), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT103), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n893), .A2(KEYINPUT103), .A3(new_n908), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1133), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n926), .A2(new_n1074), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1139), .A2(KEYINPUT40), .B1(new_n926), .B2(new_n924), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1129), .B1(new_n1140), .B2(new_n706), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n928), .A2(G330), .A3(new_n1130), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n909), .B2(new_n910), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1138), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1087), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1095), .A2(new_n1147), .A3(KEYINPUT119), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT119), .B1(new_n1095), .B2(new_n1147), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT57), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n693), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n1138), .A2(new_n1144), .A3(KEYINPUT57), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT120), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT120), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1153), .B(new_n1156), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1152), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1146), .A2(new_n983), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n762), .A2(G132), .B1(new_n798), .B2(G137), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT116), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n769), .A2(new_n344), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n780), .A2(new_n1111), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n783), .A2(new_n1109), .B1(new_n771), .B2(new_n1115), .ZN(new_n1164));
  NOR4_X1   g0964(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1168));
  AOI211_X1 g0968(.A(G33), .B(G41), .C1(new_n775), .C2(G124), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n793), .B2(new_n785), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT117), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1167), .A2(new_n1168), .A3(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n783), .A2(new_n458), .B1(new_n785), .B2(new_n372), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G97), .B2(new_n762), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n243), .A2(G41), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G283), .B2(new_n775), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n829), .A2(G107), .B1(new_n798), .B2(new_n507), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n801), .A2(G68), .B1(new_n842), .B2(G77), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1174), .A2(new_n1176), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT58), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1175), .B(new_n296), .C1(G33), .C2(G41), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n749), .B1(new_n1172), .B2(new_n1184), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT118), .Z(new_n1186));
  AOI21_X1  g0986(.A(new_n742), .B1(new_n296), .B2(new_n826), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n1130), .C2(new_n747), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1159), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1158), .A2(new_n1189), .ZN(G375));
  NAND2_X1  g0990(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n982), .B(KEYINPUT121), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n905), .A2(new_n746), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n743), .B1(G68), .B2(new_n1099), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n769), .A2(new_n296), .B1(new_n778), .B2(new_n344), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT123), .Z(new_n1196));
  OAI221_X1 g0996(.A(new_n243), .B1(new_n774), .B2(new_n1111), .C1(new_n780), .C2(new_n831), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n783), .A2(new_n836), .B1(new_n785), .B2(new_n372), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n791), .A2(new_n1115), .B1(new_n771), .B2(new_n793), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n769), .A2(new_n272), .B1(new_n780), .B2(new_n786), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT122), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n312), .B1(new_n774), .B2(new_n437), .C1(new_n245), .C2(new_n778), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n458), .A2(new_n791), .B1(new_n783), .B2(new_n767), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n270), .A2(new_n785), .B1(new_n771), .B2(new_n464), .ZN(new_n1205));
  NOR4_X1   g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1200), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1194), .B1(new_n1207), .B2(new_n749), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1191), .A2(new_n1192), .B1(new_n1193), .B2(new_n1208), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1092), .A2(new_n967), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1191), .A2(new_n1147), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1209), .B1(new_n1210), .B2(new_n1211), .ZN(G381));
  NOR4_X1   g1012(.A1(G393), .A2(G396), .A3(G384), .A4(G381), .ZN(new_n1213));
  INV_X1    g1013(.A(G390), .ZN(new_n1214));
  INV_X1    g1014(.A(G378), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  OR3_X1    g1016(.A1(new_n1216), .A2(G387), .A3(G375), .ZN(G407));
  NAND2_X1  g1017(.A1(new_n670), .A2(G213), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT124), .Z(new_n1219));
  NAND2_X1  g1019(.A1(new_n1215), .A2(new_n1219), .ZN(new_n1220));
  OAI211_X1 g1020(.A(G407), .B(G213), .C1(G375), .C2(new_n1220), .ZN(G409));
  INV_X1    g1021(.A(KEYINPUT126), .ZN(new_n1222));
  AOI21_X1  g1022(.A(G390), .B1(new_n984), .B2(new_n1007), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(G393), .B(new_n810), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(G390), .A2(new_n984), .A3(new_n1007), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1225), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1226), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1228), .B1(new_n1229), .B2(new_n1223), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1093), .A2(KEYINPUT60), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n1147), .B2(new_n1191), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1093), .A2(new_n1211), .A3(KEYINPUT60), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n692), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1209), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1237), .A2(new_n825), .A3(new_n850), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(G384), .A3(new_n1209), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1219), .A2(G2897), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1240), .B(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1095), .A2(new_n1147), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT119), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1095), .A2(new_n1147), .A3(KEYINPUT119), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1145), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n692), .B1(new_n1248), .B2(KEYINPUT57), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G378), .B(new_n1189), .C1(new_n1243), .C2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT125), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT125), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1158), .A2(new_n1252), .A3(G378), .A4(new_n1189), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1146), .A2(new_n1192), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1188), .B(new_n1254), .C1(new_n1150), .C2(new_n967), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1251), .A2(new_n1253), .B1(new_n1215), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1242), .B1(new_n1256), .B2(new_n1219), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT61), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT62), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1255), .A2(new_n1215), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1219), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1240), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1260), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1259), .A2(new_n1265), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1256), .A2(new_n1219), .A3(new_n1240), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1260), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1232), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1263), .A2(KEYINPUT63), .A3(new_n1264), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1270), .A2(new_n1258), .A3(new_n1257), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1232), .B1(new_n1267), .B2(KEYINPUT63), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1222), .B1(new_n1269), .B2(new_n1273), .ZN(new_n1274));
  OR2_X1    g1074(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1268), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1258), .B(new_n1257), .C1(new_n1267), .C2(new_n1260), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1231), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1275), .A2(new_n1278), .A3(KEYINPUT126), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1274), .A2(new_n1279), .ZN(G405));
  NAND2_X1  g1080(.A1(G375), .A2(new_n1215), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1261), .A2(new_n1281), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1282), .B(new_n1264), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(KEYINPUT127), .A3(new_n1232), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n1232), .B2(new_n1283), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT127), .B1(new_n1283), .B2(new_n1232), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(G402));
endmodule


