//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955;
  XNOR2_X1  g000(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(G101), .ZN(new_n188));
  NOR2_X1   g002(.A1(G237), .A2(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  INV_X1    g006(.A(G134), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G137), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(G137), .ZN(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT11), .A3(G134), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G131), .ZN(new_n199));
  INV_X1    g013(.A(G131), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n194), .A2(new_n197), .A3(new_n200), .A4(new_n195), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT0), .A2(G128), .ZN(new_n203));
  XNOR2_X1  g017(.A(G143), .B(G146), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT0), .B(G128), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT64), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n206), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n202), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G128), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(new_n208), .A3(new_n210), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n207), .A3(G143), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n209), .B(G146), .C1(new_n216), .C2(KEYINPUT1), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n196), .A2(G134), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n193), .A2(G137), .ZN(new_n223));
  OAI21_X1  g037(.A(G131), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n201), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n215), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g040(.A(G116), .B(G119), .Z(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT2), .B(G113), .ZN(new_n228));
  XOR2_X1   g042(.A(new_n227), .B(new_n228), .Z(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  OR2_X1    g045(.A1(new_n231), .A2(KEYINPUT28), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n229), .B1(new_n215), .B2(new_n225), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT28), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n191), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n231), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n191), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n199), .A2(new_n201), .B1(new_n206), .B2(new_n213), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n201), .A2(new_n224), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT30), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT30), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n215), .A2(new_n243), .A3(new_n225), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT65), .B1(new_n245), .B2(new_n229), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n242), .A2(new_n244), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(new_n230), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n237), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  XOR2_X1   g064(.A(KEYINPUT67), .B(KEYINPUT31), .Z(new_n251));
  AOI21_X1  g065(.A(new_n235), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n191), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n231), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n248), .B1(new_n247), .B2(new_n230), .ZN(new_n255));
  AOI211_X1 g069(.A(KEYINPUT65), .B(new_n229), .C1(new_n242), .C2(new_n244), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n257), .A2(KEYINPUT66), .A3(KEYINPUT31), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT66), .B1(new_n257), .B2(KEYINPUT31), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n252), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT68), .ZN(new_n261));
  NOR2_X1   g075(.A1(G472), .A2(G902), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n252), .B(new_n263), .C1(new_n258), .C2(new_n259), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n261), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT32), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT32), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n261), .A2(new_n267), .A3(new_n262), .A4(new_n264), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G902), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n232), .A2(new_n234), .A3(new_n191), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT29), .ZN(new_n272));
  OR2_X1    g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n246), .A2(new_n249), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n191), .B1(new_n274), .B2(new_n236), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n271), .A2(new_n272), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n270), .B(new_n273), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G472), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n269), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G953), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n280), .A2(G952), .ZN(new_n281));
  NAND2_X1  g095(.A1(G234), .A2(G237), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g097(.A(KEYINPUT21), .B(G898), .Z(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(G902), .A3(G953), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G214), .B1(G237), .B2(G902), .ZN(new_n287));
  INV_X1    g101(.A(G104), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT3), .B1(new_n288), .B2(G107), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n290));
  INV_X1    g104(.A(G107), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n291), .A3(G104), .ZN(new_n292));
  INV_X1    g106(.A(G101), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n288), .A2(G107), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n289), .A2(new_n292), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n291), .A2(G104), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n288), .A2(G107), .ZN(new_n297));
  OAI21_X1  g111(.A(G101), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  OR2_X1    g113(.A1(new_n227), .A2(new_n228), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT5), .ZN(new_n301));
  INV_X1    g115(.A(G119), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n302), .A3(G116), .ZN(new_n303));
  OAI211_X1 g117(.A(G113), .B(new_n303), .C1(new_n227), .C2(new_n301), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n299), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n289), .A2(new_n292), .A3(new_n294), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT76), .B(KEYINPUT4), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n306), .A2(G101), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n295), .A2(KEYINPUT75), .A3(KEYINPUT4), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n295), .A2(new_n310), .A3(KEYINPUT4), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n306), .A2(G101), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n308), .A2(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n305), .B1(new_n313), .B2(new_n229), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT6), .ZN(new_n315));
  XNOR2_X1  g129(.A(G110), .B(G122), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT81), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT81), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n314), .A2(new_n320), .A3(new_n315), .A4(new_n317), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n214), .A2(G125), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n221), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(G224), .A3(new_n280), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n280), .A2(G224), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n323), .A2(new_n328), .A3(new_n325), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n314), .A2(new_n317), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n305), .B(new_n316), .C1(new_n313), .C2(new_n229), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(KEYINPUT6), .A3(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n322), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT7), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n328), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n327), .A2(new_n329), .A3(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n316), .B(KEYINPUT8), .ZN(new_n338));
  INV_X1    g152(.A(new_n305), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n299), .B1(new_n300), .B2(new_n304), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n323), .A2(new_n335), .A3(new_n328), .A4(new_n325), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n337), .A2(new_n332), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n343), .A2(new_n270), .ZN(new_n344));
  OAI21_X1  g158(.A(G210), .B1(G237), .B2(G902), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n334), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n345), .B(KEYINPUT82), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n348), .B1(new_n334), .B2(new_n344), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n286), .B(new_n287), .C1(new_n347), .C2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G125), .B(G140), .ZN(new_n351));
  NAND2_X1  g165(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n353), .B(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n207), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT16), .ZN(new_n357));
  INV_X1    g171(.A(G140), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(G125), .ZN(new_n359));
  INV_X1    g173(.A(new_n351), .ZN(new_n360));
  OAI211_X1 g174(.A(G146), .B(new_n359), .C1(new_n360), .C2(new_n357), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n189), .A2(G143), .A3(G214), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(G143), .B1(new_n189), .B2(G214), .ZN(new_n364));
  OAI21_X1  g178(.A(G131), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n364), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n200), .A3(new_n362), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n356), .A2(new_n361), .A3(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n351), .B(new_n207), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n366), .A2(new_n362), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT18), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(new_n200), .ZN(new_n373));
  OAI221_X1 g187(.A(new_n370), .B1(new_n371), .B2(new_n373), .C1(new_n365), .C2(new_n372), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G113), .B(G122), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(new_n288), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n377), .B(KEYINPUT84), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT17), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n365), .A2(new_n367), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n359), .B1(new_n360), .B2(new_n357), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n207), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n371), .A2(KEYINPUT17), .A3(G131), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n382), .A2(new_n361), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n380), .A2(new_n386), .A3(new_n374), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n379), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT20), .ZN(new_n389));
  INV_X1    g203(.A(G475), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .A4(new_n270), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n377), .B1(new_n369), .B2(new_n374), .ZN(new_n392));
  INV_X1    g206(.A(new_n387), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n390), .B(new_n270), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT20), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n386), .A2(new_n374), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n397), .A2(KEYINPUT85), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n377), .B1(new_n397), .B2(KEYINPUT85), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n393), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G475), .B1(new_n400), .B2(G902), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G478), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(KEYINPUT15), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  XOR2_X1   g220(.A(KEYINPUT9), .B(G234), .Z(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G217), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n408), .A2(new_n409), .A3(G953), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G116), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G122), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(KEYINPUT14), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT90), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT86), .B1(new_n412), .B2(G122), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT86), .ZN(new_n417));
  INV_X1    g231(.A(G122), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n418), .A3(G116), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n416), .A2(new_n419), .B1(new_n413), .B2(KEYINPUT14), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n291), .B1(new_n415), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n416), .A2(new_n419), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n413), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT87), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT87), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n422), .A2(new_n425), .A3(new_n413), .ZN(new_n426));
  AOI21_X1  g240(.A(G107), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n421), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(G128), .B(G143), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(G134), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT89), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NOR3_X1   g248(.A1(new_n216), .A2(KEYINPUT13), .A3(G143), .ZN(new_n435));
  AOI211_X1 g249(.A(new_n193), .B(new_n435), .C1(KEYINPUT13), .C2(new_n429), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n429), .A2(new_n193), .ZN(new_n437));
  XOR2_X1   g251(.A(new_n437), .B(KEYINPUT88), .Z(new_n438));
  INV_X1    g252(.A(new_n427), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n424), .A2(G107), .A3(new_n426), .ZN(new_n440));
  AOI211_X1 g254(.A(new_n436), .B(new_n438), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n411), .B1(new_n434), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n443));
  INV_X1    g257(.A(new_n438), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n410), .A3(new_n433), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n406), .B1(new_n447), .B2(new_n270), .ZN(new_n448));
  AOI211_X1 g262(.A(G902), .B(new_n405), .C1(new_n442), .C2(new_n446), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n403), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n350), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n384), .A2(new_n361), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n302), .A2(G128), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT23), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(G119), .B2(new_n216), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n302), .A2(KEYINPUT23), .A3(G128), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G110), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n216), .A2(G119), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT24), .B(G110), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n453), .B(new_n459), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n462), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n458), .B2(G110), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n351), .A2(new_n207), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n361), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n467), .A2(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(KEYINPUT69), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n463), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n280), .A2(G221), .A3(G234), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(KEYINPUT22), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(new_n196), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT70), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n472), .A2(new_n196), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n196), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT70), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n470), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT71), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n481), .B(new_n482), .C1(new_n470), .C2(new_n473), .ZN(new_n483));
  OR3_X1    g297(.A1(new_n470), .A2(new_n482), .A3(new_n473), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n409), .B1(G234), .B2(new_n270), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n486), .A2(G902), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(G902), .B1(new_n483), .B2(new_n484), .ZN(new_n489));
  XOR2_X1   g303(.A(KEYINPUT72), .B(KEYINPUT25), .Z(new_n490));
  AND2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(KEYINPUT72), .A2(KEYINPUT25), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n486), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n488), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT73), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n489), .A2(new_n490), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n496), .B(new_n486), .C1(new_n492), .C2(new_n489), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT73), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n498), .A3(new_n488), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G221), .B1(new_n408), .B2(G902), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n308), .A2(new_n309), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n311), .A2(new_n312), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n214), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n299), .A2(KEYINPUT10), .A3(new_n221), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT77), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n299), .A2(new_n507), .A3(new_n221), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n295), .A2(new_n298), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT77), .B1(new_n239), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT10), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n505), .A2(new_n506), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n202), .ZN(new_n514));
  INV_X1    g328(.A(new_n202), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n505), .A2(new_n515), .A3(new_n506), .A4(new_n512), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n280), .A2(G227), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(new_n358), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT74), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(G110), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT79), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n299), .B2(new_n221), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n239), .A2(new_n509), .A3(KEYINPUT79), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n523), .A2(new_n508), .A3(new_n510), .A4(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n515), .A2(KEYINPUT78), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT12), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n516), .A2(new_n521), .ZN(new_n529));
  OAI22_X1  g343(.A1(new_n517), .A2(new_n521), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G469), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n270), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT12), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n527), .B(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n521), .B1(new_n535), .B2(new_n516), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n516), .A2(new_n521), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n514), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT80), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n521), .ZN(new_n541));
  INV_X1    g355(.A(new_n516), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n541), .B1(new_n528), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT80), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n538), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n533), .B1(new_n546), .B2(G469), .ZN(new_n547));
  NAND2_X1  g361(.A1(G469), .A2(G902), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n502), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n279), .A2(new_n452), .A3(new_n500), .A4(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(G101), .ZN(G3));
  AND2_X1   g365(.A1(new_n495), .A2(new_n499), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n261), .A2(new_n270), .A3(new_n264), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G472), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n265), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n540), .A2(new_n545), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n548), .B(new_n532), .C1(new_n556), .C2(new_n531), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n501), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n552), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n447), .A2(KEYINPUT33), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT33), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n442), .A2(new_n561), .A3(new_n446), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(G478), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n447), .A2(new_n404), .A3(new_n270), .ZN(new_n564));
  NAND2_X1  g378(.A1(G478), .A2(G902), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(new_n403), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n567), .A2(new_n286), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n345), .B1(new_n334), .B2(new_n344), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n287), .B1(new_n347), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n559), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(G104), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n573), .B(new_n575), .ZN(G6));
  XNOR2_X1  g390(.A(new_n401), .B(KEYINPUT92), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n577), .A2(new_n396), .ZN(new_n578));
  INV_X1    g392(.A(new_n450), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n579), .A3(new_n286), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT93), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n580), .A2(new_n581), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n582), .A2(new_n583), .A3(new_n570), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n559), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT35), .B(G107), .Z(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(G9));
  AND2_X1   g401(.A1(new_n261), .A2(new_n264), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n588), .A2(new_n262), .B1(new_n553), .B2(G472), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT94), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT36), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n479), .B2(new_n591), .ZN(new_n592));
  AOI211_X1 g406(.A(KEYINPUT94), .B(KEYINPUT36), .C1(new_n475), .C2(new_n478), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n470), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n478), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT70), .B1(new_n476), .B2(new_n477), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n591), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT94), .ZN(new_n598));
  INV_X1    g412(.A(new_n470), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n479), .A2(new_n590), .A3(new_n591), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n594), .A2(new_n601), .A3(new_n487), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT95), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n603), .B1(new_n493), .B2(new_n491), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT96), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT96), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n497), .A2(new_n606), .A3(new_n603), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n589), .A2(new_n608), .A3(new_n549), .A4(new_n452), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT97), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT37), .B(G110), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G12));
  INV_X1    g426(.A(new_n608), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n266), .A2(new_n268), .B1(G472), .B2(new_n277), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n613), .A2(new_n614), .A3(new_n558), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n283), .B1(new_n285), .B2(G900), .ZN(new_n616));
  AND4_X1   g430(.A1(new_n579), .A2(new_n578), .A3(new_n571), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G128), .ZN(G30));
  NOR3_X1   g433(.A1(new_n231), .A2(new_n233), .A3(new_n191), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n274), .A2(new_n236), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n620), .B1(new_n621), .B2(new_n191), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n622), .A2(KEYINPUT98), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n270), .B1(new_n622), .B2(KEYINPUT98), .ZN(new_n624));
  OAI21_X1  g438(.A(G472), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n269), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(new_n604), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n347), .A2(new_n349), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT38), .ZN(new_n630));
  INV_X1    g444(.A(new_n287), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n579), .A2(new_n402), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(KEYINPUT99), .B1(new_n628), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n604), .ZN(new_n635));
  AND4_X1   g449(.A1(KEYINPUT99), .A2(new_n626), .A3(new_n633), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n616), .B(KEYINPUT39), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n549), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT40), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n634), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(new_n209), .ZN(G45));
  INV_X1    g455(.A(new_n566), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n402), .A3(new_n616), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT100), .B1(new_n643), .B2(new_n570), .ZN(new_n644));
  INV_X1    g458(.A(new_n616), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n566), .A2(new_n403), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(new_n571), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n615), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G146), .ZN(G48));
  NAND2_X1  g465(.A1(new_n530), .A2(new_n270), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(G469), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n653), .A2(new_n532), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n501), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n614), .A2(new_n552), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT101), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n657), .A3(new_n572), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n657), .B1(new_n656), .B2(new_n572), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT41), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n662), .B(G113), .Z(G15));
  NAND2_X1  g477(.A1(new_n584), .A2(new_n656), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G116), .ZN(G18));
  NOR2_X1   g479(.A1(new_n655), .A2(new_n570), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n286), .ZN(new_n667));
  NOR4_X1   g481(.A1(new_n667), .A2(new_n613), .A3(new_n614), .A4(new_n451), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(new_n302), .ZN(G21));
  XNOR2_X1  g483(.A(new_n262), .B(KEYINPUT102), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n257), .A2(KEYINPUT31), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n670), .B1(new_n252), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n554), .A2(KEYINPUT103), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n553), .A2(new_n674), .A3(G472), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n672), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n494), .ZN(new_n677));
  INV_X1    g491(.A(new_n632), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n679), .A2(new_n667), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G122), .ZN(G24));
  NAND4_X1  g495(.A1(new_n676), .A2(new_n604), .A3(new_n646), .A4(new_n666), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT104), .B(G125), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G27));
  NOR2_X1   g498(.A1(new_n614), .A2(new_n552), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n548), .B(KEYINPUT105), .Z(new_n687));
  NAND3_X1  g501(.A1(new_n543), .A2(G469), .A3(new_n538), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n532), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n501), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT106), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n347), .A2(new_n349), .A3(new_n631), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n643), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n685), .A2(new_n686), .A3(new_n691), .A4(new_n694), .ZN(new_n695));
  AND4_X1   g509(.A1(new_n279), .A2(new_n691), .A3(new_n677), .A4(new_n694), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n695), .B1(new_n696), .B2(new_n686), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n200), .ZN(G33));
  AND3_X1   g512(.A1(new_n578), .A2(new_n579), .A3(new_n616), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n685), .A2(new_n699), .A3(new_n691), .A4(new_n692), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT107), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n193), .ZN(G36));
  NAND3_X1  g516(.A1(new_n543), .A2(KEYINPUT45), .A3(new_n538), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n703), .B(G469), .C1(new_n546), .C2(KEYINPUT45), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(KEYINPUT46), .A3(new_n687), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n532), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n705), .A2(KEYINPUT108), .A3(new_n532), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n704), .A2(new_n687), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n708), .B(new_n709), .C1(new_n710), .C2(KEYINPUT46), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n501), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n566), .A2(new_n402), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT43), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n555), .A3(new_n604), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n713), .A2(new_n637), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n692), .B1(new_n716), .B2(new_n717), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n720), .A2(KEYINPUT109), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(KEYINPUT109), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n196), .ZN(G39));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n711), .A2(new_n726), .A3(new_n501), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n726), .B1(new_n711), .B2(new_n501), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n725), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n712), .A2(KEYINPUT110), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(KEYINPUT47), .A3(new_n727), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n279), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n500), .A2(new_n643), .A3(new_n693), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G140), .ZN(G42));
  INV_X1    g550(.A(new_n283), .ZN(new_n737));
  AND4_X1   g551(.A1(new_n737), .A2(new_n676), .A3(new_n677), .A4(new_n715), .ZN(new_n738));
  INV_X1    g552(.A(new_n655), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n739), .A2(new_n630), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(new_n631), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT117), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT117), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n738), .A2(new_n744), .A3(new_n631), .A4(new_n740), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT118), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT118), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n742), .A2(new_n748), .A3(new_n743), .A4(new_n745), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n747), .B(new_n749), .C1(new_n743), .C2(new_n741), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n626), .A2(new_n655), .A3(new_n693), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n737), .A3(new_n500), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n752), .A2(new_n402), .A3(new_n642), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n676), .A2(new_n604), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  AND4_X1   g569(.A1(new_n737), .A2(new_n715), .A3(new_n739), .A4(new_n692), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n654), .A2(new_n502), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n730), .A2(new_n732), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n692), .A3(new_n738), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n750), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n750), .A2(KEYINPUT51), .A3(new_n757), .A4(new_n760), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n396), .B(new_n401), .C1(new_n448), .C2(new_n449), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT113), .B1(new_n350), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n450), .A2(new_n402), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n334), .A2(new_n344), .ZN(new_n769));
  INV_X1    g583(.A(new_n348), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n631), .B1(new_n771), .B2(new_n346), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n768), .A2(new_n772), .A3(new_n773), .A4(new_n286), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n767), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n775), .A2(new_n589), .A3(new_n500), .A4(new_n549), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n609), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n776), .A2(new_n609), .A3(KEYINPUT114), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n668), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n555), .A2(new_n558), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n772), .A3(new_n500), .A4(new_n568), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n784), .A2(new_n550), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n781), .A2(new_n680), .A3(new_n782), .A4(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n664), .B1(new_n659), .B2(new_n660), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n615), .A2(new_n450), .A3(new_n578), .A4(new_n616), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n676), .A2(new_n604), .A3(new_n646), .A4(new_n691), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n693), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n700), .B(new_n695), .C1(new_n696), .C2(new_n686), .ZN(new_n791));
  NOR4_X1   g605(.A1(new_n786), .A2(new_n787), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n558), .B1(new_n269), .B2(new_n278), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n793), .B(new_n608), .C1(new_n617), .C2(new_n649), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n690), .A2(new_n645), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n678), .A2(new_n571), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n626), .A2(new_n635), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n794), .A2(new_n682), .A3(KEYINPUT52), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n794), .A2(new_n682), .A3(new_n798), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n801), .B(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT53), .B1(new_n792), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n799), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n804), .A2(KEYINPUT116), .A3(new_n799), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n776), .A2(new_n609), .A3(KEYINPUT114), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT114), .B1(new_n776), .B2(new_n609), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n550), .B(new_n784), .C1(new_n679), .C2(new_n667), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n814), .A2(new_n815), .A3(new_n668), .ZN(new_n816));
  INV_X1    g630(.A(new_n790), .ZN(new_n817));
  INV_X1    g631(.A(new_n660), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n818), .A2(new_n658), .B1(new_n584), .B2(new_n656), .ZN(new_n819));
  INV_X1    g633(.A(new_n791), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n816), .A2(new_n817), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n811), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT54), .B1(new_n806), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n822), .B1(new_n811), .B2(new_n821), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n786), .A2(new_n787), .A3(new_n791), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n805), .A2(new_n826), .A3(KEYINPUT53), .A4(new_n817), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n825), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n614), .A2(new_n494), .ZN(new_n830));
  NAND2_X1  g644(.A1(KEYINPUT119), .A2(KEYINPUT48), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n756), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(KEYINPUT119), .A2(KEYINPUT48), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n752), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n567), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n281), .ZN(new_n837));
  AOI211_X1 g651(.A(new_n834), .B(new_n837), .C1(new_n666), .C2(new_n738), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n824), .A2(new_n829), .A3(new_n838), .ZN(new_n839));
  OAI22_X1  g653(.A1(new_n765), .A2(new_n839), .B1(G952), .B2(G953), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT49), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n654), .A2(new_n841), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n627), .A2(new_n630), .A3(new_n714), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n677), .A2(new_n287), .A3(new_n501), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT111), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n843), .B(new_n845), .C1(new_n841), .C2(new_n654), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(KEYINPUT112), .Z(new_n847));
  NAND2_X1  g661(.A1(new_n840), .A2(new_n847), .ZN(G75));
  NOR2_X1   g662(.A1(new_n280), .A2(G952), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n270), .B1(new_n825), .B2(new_n827), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT56), .B1(new_n851), .B2(G210), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n322), .A2(new_n333), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(new_n330), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT55), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n850), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT56), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n851), .B2(new_n770), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n859), .A2(KEYINPUT120), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(KEYINPUT120), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n856), .B1(new_n860), .B2(new_n861), .ZN(G51));
  XOR2_X1   g676(.A(new_n687), .B(KEYINPUT57), .Z(new_n863));
  INV_X1    g677(.A(new_n829), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n828), .B1(new_n825), .B2(new_n827), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n530), .ZN(new_n867));
  INV_X1    g681(.A(new_n704), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n851), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n849), .B1(new_n867), .B2(new_n869), .ZN(G54));
  NAND2_X1  g684(.A1(new_n825), .A2(new_n827), .ZN(new_n871));
  AND2_X1   g685(.A1(KEYINPUT58), .A2(G475), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n871), .A2(G902), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n850), .B1(new_n873), .B2(new_n388), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n851), .A2(new_n872), .ZN(new_n875));
  INV_X1    g689(.A(new_n388), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT121), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n873), .A2(new_n878), .A3(new_n388), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n874), .B1(new_n877), .B2(new_n879), .ZN(G60));
  XOR2_X1   g694(.A(new_n565), .B(KEYINPUT59), .Z(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n824), .B2(new_n829), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n560), .A2(new_n562), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT122), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n850), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n865), .ZN(new_n887));
  AOI211_X1 g701(.A(new_n884), .B(new_n881), .C1(new_n887), .C2(new_n829), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n886), .A2(new_n888), .ZN(G63));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n890));
  NAND2_X1  g704(.A1(G217), .A2(G902), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT123), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT60), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n871), .A2(new_n601), .A3(new_n594), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n850), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n485), .B1(new_n871), .B2(new_n893), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n890), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n896), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n898), .A2(KEYINPUT61), .A3(new_n850), .A4(new_n894), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n899), .ZN(G66));
  NAND2_X1  g714(.A1(new_n284), .A2(G224), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(G953), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n786), .A2(new_n787), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n902), .B1(new_n903), .B2(G953), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT124), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n853), .B1(G898), .B2(new_n280), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n905), .B(new_n906), .ZN(G69));
  XNOR2_X1  g721(.A(new_n245), .B(new_n355), .ZN(new_n908));
  INV_X1    g722(.A(G227), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n280), .B1(new_n910), .B2(G900), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n723), .B1(new_n733), .B2(new_n734), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n567), .A2(new_n768), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n638), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT125), .B1(new_n567), .B2(new_n768), .ZN(new_n916));
  AND4_X1   g730(.A1(new_n685), .A2(new_n915), .A3(new_n692), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n794), .A2(new_n682), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n628), .A2(new_n633), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT99), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n636), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g738(.A(KEYINPUT62), .B(new_n919), .C1(new_n924), .C2(new_n639), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n640), .B2(new_n918), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n917), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(G953), .B1(new_n912), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n911), .B1(new_n929), .B2(new_n908), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n713), .A2(new_n637), .A3(new_n830), .A4(new_n797), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n912), .A2(new_n919), .A3(new_n931), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n932), .A2(G953), .A3(new_n791), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(G227), .B2(G953), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n930), .B1(new_n934), .B2(new_n908), .ZN(G72));
  NAND3_X1  g749(.A1(new_n274), .A2(new_n236), .A3(new_n253), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT126), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n912), .A2(new_n826), .A3(new_n919), .A4(new_n931), .ZN(new_n938));
  NAND2_X1  g752(.A1(G472), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT63), .Z(new_n940));
  AOI21_X1  g754(.A(new_n937), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n621), .A2(new_n191), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n912), .A2(new_n903), .A3(new_n928), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(new_n940), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n941), .A2(new_n944), .A3(new_n849), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n792), .A2(new_n805), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n822), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n792), .A2(KEYINPUT53), .A3(new_n809), .A4(new_n810), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n949), .A2(new_n942), .A3(new_n940), .A4(new_n936), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n936), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n947), .B2(new_n948), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n954), .A2(KEYINPUT127), .A3(new_n942), .A4(new_n940), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n945), .A2(new_n952), .A3(new_n955), .ZN(G57));
endmodule


