//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n819, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT98), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n204), .A2(G1gat), .ZN(new_n205));
  INV_X1    g004(.A(G8gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(new_n207), .B2(G1gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n205), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT100), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n205), .A2(KEYINPUT99), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(new_n208), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n205), .A2(KEYINPUT99), .ZN(new_n214));
  OAI21_X1  g013(.A(G8gat), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n211), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT14), .ZN(new_n218));
  XOR2_X1   g017(.A(KEYINPUT97), .B(G29gat), .Z(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n218), .B1(G36gat), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n221), .A2(KEYINPUT15), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(KEYINPUT15), .ZN(new_n223));
  XNOR2_X1  g022(.A(G43gat), .B(G50gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(KEYINPUT17), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n216), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G229gat), .A2(G233gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n211), .A2(new_n215), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n227), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT101), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n234), .A2(KEYINPUT18), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT102), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n211), .A2(new_n215), .A3(new_n225), .A4(new_n226), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n232), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n230), .B(KEYINPUT13), .Z(new_n240));
  NAND3_X1  g039(.A1(new_n231), .A2(KEYINPUT102), .A3(new_n227), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n235), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n229), .A2(new_n232), .A3(new_n230), .A4(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n236), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G113gat), .B(G141gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(G197gat), .ZN(new_n247));
  XOR2_X1   g046(.A(KEYINPUT11), .B(G169gat), .Z(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n249), .B(KEYINPUT12), .Z(new_n250));
  NAND2_X1  g049(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n250), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n236), .A2(new_n242), .A3(new_n252), .A4(new_n244), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT35), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT94), .ZN(new_n257));
  XNOR2_X1  g056(.A(G78gat), .B(G106gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT31), .B(G50gat), .ZN(new_n259));
  XOR2_X1   g058(.A(new_n258), .B(new_n259), .Z(new_n260));
  NAND2_X1  g059(.A1(G211gat), .A2(G218gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT22), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G197gat), .A2(G204gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(G197gat), .A2(G204gat), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n263), .B(KEYINPUT77), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G211gat), .ZN(new_n268));
  INV_X1    g067(.A(G218gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT76), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n271), .A3(new_n261), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n271), .B1(new_n270), .B2(new_n261), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n267), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n266), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n276), .A2(new_n264), .B1(new_n262), .B2(new_n261), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(KEYINPUT77), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n274), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n280), .A2(new_n277), .A3(KEYINPUT77), .A4(new_n272), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G141gat), .B(G148gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285));
  INV_X1    g084(.A(G155gat), .ZN(new_n286));
  INV_X1    g085(.A(G162gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n284), .A2(KEYINPUT83), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(G141gat), .B(G148gat), .Z(new_n290));
  INV_X1    g089(.A(KEYINPUT83), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT84), .B(G155gat), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT2), .B1(new_n293), .B2(new_n287), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n289), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  OR2_X1    g094(.A1(KEYINPUT81), .A2(KEYINPUT2), .ZN(new_n296));
  NAND2_X1  g095(.A1(KEYINPUT81), .A2(KEYINPUT2), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n296), .A2(new_n297), .A3(new_n285), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n290), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT80), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(KEYINPUT80), .A2(G155gat), .A3(G162gat), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n301), .A2(new_n302), .A3(new_n288), .ZN(new_n303));
  AND3_X1   g102(.A1(new_n299), .A2(KEYINPUT82), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT82), .B1(new_n299), .B2(new_n303), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n295), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT85), .B1(new_n306), .B2(KEYINPUT3), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n299), .A2(new_n303), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT82), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n299), .A2(KEYINPUT82), .A3(new_n303), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT85), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .A4(new_n295), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT29), .B1(new_n307), .B2(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n289), .A2(new_n292), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n310), .A2(new_n311), .B1(new_n317), .B2(new_n294), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT87), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n306), .A2(KEYINPUT87), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n281), .B(new_n323), .C1(new_n275), .C2(new_n278), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT90), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT3), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n279), .A2(KEYINPUT90), .A3(new_n323), .A4(new_n281), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI22_X1  g127(.A1(new_n283), .A2(new_n316), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(G228gat), .A2(G233gat), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n307), .A2(new_n315), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n323), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n282), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT91), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT3), .B1(new_n324), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(new_n335), .B2(new_n324), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n331), .B1(new_n337), .B2(new_n306), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n329), .A2(new_n331), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT92), .B(G22gat), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n260), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT93), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n334), .A2(new_n338), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n283), .B1(new_n332), .B2(new_n323), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n320), .A2(new_n321), .B1(new_n326), .B2(new_n327), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n331), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n342), .B1(new_n347), .B2(G22gat), .ZN(new_n348));
  INV_X1    g147(.A(G22gat), .ZN(new_n349));
  AOI211_X1 g148(.A(KEYINPUT93), .B(new_n349), .C1(new_n343), .C2(new_n346), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n257), .B(new_n341), .C1(new_n348), .C2(new_n350), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n343), .A2(new_n346), .A3(new_n340), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n340), .B1(new_n343), .B2(new_n346), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n260), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT94), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n343), .A2(new_n346), .A3(new_n340), .ZN(new_n356));
  INV_X1    g155(.A(new_n260), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT93), .B1(new_n339), .B2(new_n349), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n347), .A2(new_n342), .A3(G22gat), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n351), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT32), .ZN(new_n363));
  XNOR2_X1  g162(.A(G15gat), .B(G43gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(G71gat), .B(G99gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT33), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OR2_X1    g167(.A1(G113gat), .A2(G120gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(G113gat), .A2(G120gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(KEYINPUT69), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT69), .ZN(new_n372));
  AND2_X1   g171(.A1(G113gat), .A2(G120gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(G113gat), .A2(G120gat), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT1), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n371), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G127gat), .B(G134gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT70), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n369), .A2(new_n381), .A3(new_n370), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT70), .B1(new_n373), .B2(new_n374), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n382), .A2(new_n383), .A3(new_n376), .A4(new_n378), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT24), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT24), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n388), .A2(G183gat), .A3(G190gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  OR2_X1    g189(.A1(G183gat), .A2(G190gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G169gat), .ZN(new_n393));
  INV_X1    g192(.A(G176gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT66), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n396), .B1(new_n397), .B2(KEYINPUT23), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT23), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n399), .A2(KEYINPUT66), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n395), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT65), .B(G169gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n399), .A2(G176gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n392), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  XOR2_X1   g204(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT23), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT25), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n397), .A2(KEYINPUT23), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n399), .A2(KEYINPUT66), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n411), .A3(new_n396), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n409), .B1(new_n395), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT67), .B(G190gat), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n390), .B1(new_n414), .B2(G183gat), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n405), .A2(new_n407), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT26), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n395), .A2(new_n417), .A3(new_n396), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT26), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n418), .A2(new_n386), .A3(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n421));
  XOR2_X1   g220(.A(KEYINPUT27), .B(G183gat), .Z(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(new_n414), .ZN(new_n423));
  XOR2_X1   g222(.A(KEYINPUT67), .B(G190gat), .Z(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT27), .B(G183gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n421), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n420), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n385), .B1(new_n416), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n380), .A2(new_n384), .ZN(new_n432));
  INV_X1    g231(.A(new_n420), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n422), .A2(new_n414), .A3(new_n421), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n426), .B1(new_n424), .B2(new_n425), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n390), .A2(new_n391), .B1(new_n402), .B2(new_n403), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n406), .B1(new_n437), .B2(new_n401), .ZN(new_n438));
  INV_X1    g237(.A(new_n409), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n415), .A2(new_n401), .A3(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n432), .B(new_n436), .C1(new_n438), .C2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n429), .A2(new_n431), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT71), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT71), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n429), .A2(new_n441), .A3(new_n444), .A4(new_n431), .ZN(new_n445));
  AOI211_X1 g244(.A(new_n363), .B(new_n368), .C1(new_n443), .C2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n431), .B1(new_n429), .B2(new_n441), .ZN(new_n447));
  NOR2_X1   g246(.A1(KEYINPUT74), .A2(KEYINPUT34), .ZN(new_n448));
  AND2_X1   g247(.A1(KEYINPUT74), .A2(KEYINPUT34), .ZN(new_n449));
  NOR3_X1   g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n447), .A2(new_n449), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n443), .A2(new_n445), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n366), .B1(new_n453), .B2(new_n367), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT72), .B1(new_n453), .B2(KEYINPUT32), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT72), .ZN(new_n456));
  AOI211_X1 g255(.A(new_n456), .B(new_n363), .C1(new_n443), .C2(new_n445), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n454), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT73), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT73), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n460), .B(new_n454), .C1(new_n455), .C2(new_n457), .ZN(new_n461));
  AOI211_X1 g260(.A(new_n446), .B(new_n452), .C1(new_n459), .C2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n452), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n459), .A2(new_n461), .ZN(new_n464));
  INV_X1    g263(.A(new_n446), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR3_X1   g265(.A1(new_n362), .A2(new_n462), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(G226gat), .A2(G233gat), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n416), .A2(new_n428), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(KEYINPUT29), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT78), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n436), .B1(new_n438), .B2(new_n440), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n472), .A2(new_n323), .B1(G226gat), .B2(G233gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n469), .A2(new_n468), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n283), .B(new_n471), .C1(new_n475), .C2(KEYINPUT78), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n470), .B1(new_n469), .B2(new_n468), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n282), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G8gat), .B(G36gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(G64gat), .B(G92gat), .ZN(new_n481));
  XOR2_X1   g280(.A(new_n480), .B(new_n481), .Z(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT30), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n476), .A2(new_n478), .A3(new_n482), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT79), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n486), .B2(new_n485), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n486), .A2(new_n488), .A3(new_n485), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT96), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n318), .A2(new_n385), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT4), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n320), .A2(new_n385), .A3(new_n321), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n496), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(G225gat), .A2(G233gat), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n385), .B1(new_n306), .B2(KEYINPUT3), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n332), .A2(KEYINPUT86), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT86), .B1(new_n332), .B2(new_n502), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n498), .B(new_n501), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(G1gat), .B(G29gat), .Z(new_n506));
  XNOR2_X1  g305(.A(G57gat), .B(G85gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT89), .B(KEYINPUT0), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n500), .B1(new_n494), .B2(new_n495), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(new_n497), .B2(new_n495), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n332), .A2(new_n502), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT86), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n332), .A2(KEYINPUT86), .A3(new_n502), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n306), .A2(new_n432), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n494), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT88), .B1(new_n520), .B2(new_n500), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n522));
  AOI211_X1 g321(.A(new_n522), .B(new_n499), .C1(new_n494), .C2(new_n519), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT5), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n505), .B(new_n511), .C1(new_n518), .C2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT6), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n322), .A2(KEYINPUT4), .A3(new_n385), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n528), .B(new_n512), .C1(new_n503), .C2(new_n504), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT5), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n494), .A2(new_n519), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n522), .B1(new_n531), .B2(new_n499), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n520), .A2(KEYINPUT88), .A3(new_n500), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n511), .B1(new_n535), .B2(new_n505), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n527), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n505), .B1(new_n518), .B2(new_n524), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n538), .A2(KEYINPUT6), .A3(new_n510), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n492), .B(new_n493), .C1(new_n537), .C2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n256), .B1(new_n467), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n464), .A2(new_n465), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n452), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n464), .A2(new_n465), .A3(new_n463), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR4_X1   g345(.A1(new_n546), .A2(new_n540), .A3(new_n362), .A4(KEYINPUT35), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT36), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n544), .A2(KEYINPUT75), .A3(new_n549), .A4(new_n545), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(KEYINPUT75), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n549), .A2(KEYINPUT75), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n551), .B(new_n552), .C1(new_n466), .C2(new_n462), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n492), .B1(new_n537), .B2(new_n539), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n362), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n550), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT95), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT95), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n550), .A2(new_n553), .A3(new_n555), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n538), .A2(new_n510), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(new_n526), .A3(new_n525), .ZN(new_n561));
  INV_X1    g360(.A(new_n486), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n483), .B1(new_n479), .B2(KEYINPUT37), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n282), .B(new_n471), .C1(new_n475), .C2(KEYINPUT78), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT37), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n566), .B1(new_n477), .B2(new_n283), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT38), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n562), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n527), .A2(new_n536), .ZN(new_n570));
  INV_X1    g369(.A(new_n479), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n571), .A2(new_n566), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT38), .B1(new_n572), .B2(new_n563), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n561), .A2(new_n569), .A3(new_n570), .A4(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n482), .B1(new_n476), .B2(new_n478), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n575), .B1(new_n562), .B2(KEYINPUT30), .ZN(new_n576));
  INV_X1    g375(.A(new_n491), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n576), .B1(new_n577), .B2(new_n489), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT40), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n498), .B1(new_n503), .B2(new_n504), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT39), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(new_n581), .A3(new_n500), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n511), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n531), .A2(new_n499), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT39), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n585), .B1(new_n580), .B2(new_n500), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n579), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n588), .A2(KEYINPUT40), .A3(new_n511), .A4(new_n582), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n578), .A2(new_n587), .A3(new_n589), .A4(new_n560), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n341), .B1(new_n348), .B2(new_n350), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n591), .A2(KEYINPUT94), .A3(new_n354), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n574), .A2(new_n590), .A3(new_n592), .A4(new_n351), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n557), .A2(new_n559), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n255), .B1(new_n548), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(G57gat), .B(G64gat), .ZN(new_n597));
  XOR2_X1   g396(.A(G71gat), .B(G78gat), .Z(new_n598));
  INV_X1    g397(.A(KEYINPUT103), .ZN(new_n599));
  AOI211_X1 g398(.A(new_n596), .B(new_n597), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n598), .A2(new_n599), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(KEYINPUT21), .ZN(new_n603));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(G127gat), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n231), .B1(KEYINPUT21), .B2(new_n602), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(new_n286), .ZN(new_n610));
  XNOR2_X1  g409(.A(G183gat), .B(G211gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n608), .B(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT104), .B(KEYINPUT7), .ZN(new_n615));
  NAND2_X1  g414(.A1(G85gat), .A2(G92gat), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  AND2_X1   g417(.A1(G99gat), .A2(G106gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(G85gat), .ZN(new_n621));
  INV_X1    g420(.A(G92gat), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n620), .A2(KEYINPUT8), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n617), .A2(new_n618), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(G99gat), .A2(G106gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n619), .A2(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n228), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n627), .A2(new_n628), .ZN(new_n631));
  AND2_X1   g430(.A1(G232gat), .A2(G233gat), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n227), .A2(new_n631), .B1(KEYINPUT41), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G190gat), .B(G218gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT105), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n634), .B(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n638));
  XNOR2_X1  g437(.A(G134gat), .B(G162gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(G230gat), .ZN(new_n645));
  INV_X1    g444(.A(G233gat), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n602), .ZN(new_n648));
  INV_X1    g447(.A(new_n602), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n629), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n651), .A2(KEYINPUT10), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n631), .A2(KEYINPUT10), .A3(new_n602), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n647), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n656), .B(new_n657), .Z(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n651), .A2(new_n647), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n655), .B(new_n663), .C1(new_n662), .C2(new_n661), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n659), .B1(new_n654), .B2(new_n661), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n614), .A2(new_n644), .A3(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n668), .A2(KEYINPUT107), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(KEYINPUT107), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n595), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n537), .A2(new_n539), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g474(.A(KEYINPUT16), .B(G8gat), .Z(new_n676));
  NAND3_X1  g475(.A1(new_n672), .A2(new_n578), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(KEYINPUT108), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n679), .A2(KEYINPUT108), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n206), .B1(new_n672), .B2(new_n578), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n677), .B1(new_n682), .B2(new_n678), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n680), .B1(new_n681), .B2(new_n683), .ZN(G1325gat));
  INV_X1    g483(.A(new_n672), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n550), .A2(new_n553), .A3(KEYINPUT109), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT109), .B1(new_n550), .B2(new_n553), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(G15gat), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n546), .A2(G15gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n685), .B2(new_n690), .ZN(G1326gat));
  NAND2_X1  g490(.A1(new_n672), .A2(new_n362), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT43), .B(G22gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  NOR3_X1   g493(.A1(new_n614), .A2(new_n644), .A3(new_n666), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n595), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n673), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n696), .A2(new_n697), .A3(new_n220), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT45), .Z(new_n699));
  NAND2_X1  g498(.A1(new_n593), .A2(new_n555), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n686), .A2(new_n687), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n542), .A2(new_n547), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n643), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n548), .A2(new_n594), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n644), .A2(new_n704), .ZN(new_n706));
  AOI22_X1  g505(.A1(new_n703), .A2(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT110), .B1(new_n251), .B2(new_n253), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n251), .A2(KEYINPUT110), .A3(new_n253), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n614), .A2(new_n666), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n707), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n220), .B1(new_n713), .B2(new_n697), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n714), .ZN(G1328gat));
  NOR3_X1   g514(.A1(new_n696), .A2(G36gat), .A3(new_n492), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT46), .ZN(new_n717));
  OAI21_X1  g516(.A(G36gat), .B1(new_n713), .B2(new_n492), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(G1329gat));
  NOR3_X1   g518(.A1(new_n696), .A2(G43gat), .A3(new_n546), .ZN(new_n720));
  INV_X1    g519(.A(new_n688), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n707), .A2(new_n721), .A3(new_n711), .A4(new_n712), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n720), .B1(new_n722), .B2(G43gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g523(.A(new_n362), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n696), .A2(G50gat), .A3(new_n725), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n707), .A2(new_n362), .A3(new_n711), .A4(new_n712), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(G50gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g528(.A1(new_n701), .A2(new_n702), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n614), .A2(new_n644), .ZN(new_n731));
  NOR4_X1   g530(.A1(new_n730), .A2(new_n731), .A3(new_n667), .A4(new_n711), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n673), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g533(.A(new_n492), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n736), .B(new_n737), .Z(G1333gat));
  NAND2_X1  g537(.A1(new_n732), .A2(new_n721), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n546), .A2(G71gat), .ZN(new_n740));
  AOI22_X1  g539(.A1(new_n739), .A2(G71gat), .B1(new_n732), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g541(.A1(new_n732), .A2(new_n362), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g543(.A1(new_n711), .A2(new_n614), .A3(new_n667), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n707), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G85gat), .B1(new_n746), .B2(new_n697), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n711), .A2(new_n614), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n643), .B(new_n748), .C1(new_n701), .C2(new_n702), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT51), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n673), .A2(new_n621), .A3(new_n666), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n747), .B1(new_n750), .B2(new_n751), .ZN(G1336gat));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n749), .B(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n754), .A2(new_n622), .A3(new_n578), .A4(new_n666), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n746), .A2(new_n492), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n622), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n755), .B(new_n758), .C1(new_n756), .C2(new_n622), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(G1337gat));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n688), .ZN(new_n763));
  XOR2_X1   g562(.A(KEYINPUT112), .B(G99gat), .Z(new_n764));
  NAND4_X1  g563(.A1(new_n544), .A2(new_n545), .A3(new_n666), .A4(new_n764), .ZN(new_n765));
  OAI22_X1  g564(.A1(new_n763), .A2(new_n764), .B1(new_n750), .B2(new_n765), .ZN(G1338gat));
  NOR3_X1   g565(.A1(new_n725), .A2(G106gat), .A3(new_n667), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n754), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n703), .A2(new_n704), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n705), .A2(new_n706), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n769), .A2(new_n362), .A3(new_n770), .A4(new_n745), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n771), .A2(G106gat), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT53), .B1(new_n768), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(KEYINPUT113), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n707), .A2(new_n775), .A3(new_n362), .A4(new_n745), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n774), .A2(G106gat), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT53), .B1(new_n754), .B2(new_n767), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n778), .B1(new_n777), .B2(new_n779), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n773), .B1(new_n780), .B2(new_n781), .ZN(G1339gat));
  NAND3_X1  g581(.A1(new_n652), .A2(new_n647), .A3(new_n653), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n655), .A2(KEYINPUT54), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n658), .B1(new_n654), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n784), .A2(KEYINPUT55), .A3(new_n786), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n664), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n710), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n793), .B2(new_n708), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n240), .B1(new_n239), .B2(new_n241), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n230), .B1(new_n229), .B2(new_n232), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n249), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n253), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n667), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n643), .B1(new_n794), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n798), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n792), .A2(new_n643), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n613), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n668), .A2(new_n711), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n697), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n546), .A2(new_n362), .A3(new_n578), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n811), .A2(G113gat), .A3(new_n254), .ZN(new_n812));
  AOI21_X1  g611(.A(G113gat), .B1(new_n811), .B2(new_n711), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(G1340gat));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815));
  OAI22_X1  g614(.A1(new_n810), .A2(new_n667), .B1(new_n815), .B2(G120gat), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(G120gat), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n816), .B(new_n817), .ZN(G1341gat));
  NAND2_X1  g617(.A1(new_n811), .A2(new_n614), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(G127gat), .ZN(G1342gat));
  AOI211_X1 g619(.A(new_n644), .B(new_n810), .C1(KEYINPUT56), .C2(G134gat), .ZN(new_n821));
  NOR2_X1   g620(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n821), .B(new_n822), .ZN(G1343gat));
  NAND2_X1  g622(.A1(new_n805), .A2(new_n807), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n725), .A2(new_n578), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n673), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n255), .A2(G141gat), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT118), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n826), .A2(new_n721), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(KEYINPUT58), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n255), .A2(new_n791), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n644), .B1(new_n831), .B2(new_n799), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n614), .B1(new_n832), .B2(new_n803), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n362), .B1(new_n833), .B2(new_n806), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT57), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n791), .B1(new_n709), .B2(new_n710), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n644), .B1(new_n837), .B2(new_n799), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n614), .B1(new_n838), .B2(new_n803), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n836), .B(new_n362), .C1(new_n839), .C2(new_n806), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n721), .A2(new_n697), .A3(new_n578), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n835), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G141gat), .B1(new_n842), .B2(new_n255), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n830), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n835), .A2(new_n840), .A3(new_n711), .A4(new_n841), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n845), .A2(KEYINPUT117), .A3(G141gat), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT117), .B1(new_n845), .B2(G141gat), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n846), .A2(new_n847), .A3(new_n829), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n844), .B1(new_n848), .B2(new_n849), .ZN(G1344gat));
  NOR2_X1   g649(.A1(new_n826), .A2(new_n721), .ZN(new_n851));
  INV_X1    g650(.A(G148gat), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n852), .A3(new_n666), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT119), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n824), .A2(new_n362), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT57), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n669), .A2(new_n255), .A3(new_n670), .ZN(new_n858));
  OR3_X1    g657(.A1(new_n644), .A2(KEYINPUT120), .A3(new_n791), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT120), .B1(new_n644), .B2(new_n791), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n802), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n614), .B1(new_n861), .B2(new_n832), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n836), .B(new_n362), .C1(new_n858), .C2(new_n862), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n857), .A2(new_n666), .A3(new_n841), .A4(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n855), .B1(new_n864), .B2(G148gat), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n842), .A2(new_n667), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n866), .A2(KEYINPUT59), .A3(new_n852), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n854), .B1(new_n865), .B2(new_n867), .ZN(G1345gat));
  INV_X1    g667(.A(new_n293), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(new_n851), .B2(new_n614), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n842), .A2(new_n293), .A3(new_n613), .ZN(new_n871));
  OR3_X1    g670(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT121), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT121), .B1(new_n870), .B2(new_n871), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1346gat));
  AOI21_X1  g673(.A(G162gat), .B1(new_n851), .B2(new_n643), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n842), .A2(new_n287), .A3(new_n644), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(G1347gat));
  AOI21_X1  g676(.A(new_n362), .B1(new_n805), .B2(new_n807), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n546), .A2(new_n673), .A3(new_n492), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n402), .A3(new_n711), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n879), .B(KEYINPUT122), .Z(new_n882));
  NAND2_X1  g681(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(G169gat), .B1(new_n883), .B2(new_n255), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(new_n884), .ZN(G1348gat));
  NAND3_X1  g684(.A1(new_n880), .A2(new_n394), .A3(new_n666), .ZN(new_n886));
  OAI21_X1  g685(.A(G176gat), .B1(new_n883), .B2(new_n667), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT123), .ZN(G1349gat));
  NAND3_X1  g688(.A1(new_n880), .A2(new_n425), .A3(new_n614), .ZN(new_n890));
  OAI21_X1  g689(.A(G183gat), .B1(new_n883), .B2(new_n613), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g692(.A1(new_n880), .A2(new_n424), .A3(new_n643), .ZN(new_n894));
  OAI21_X1  g693(.A(G190gat), .B1(new_n883), .B2(new_n644), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n895), .A2(KEYINPUT61), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(KEYINPUT61), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(G1351gat));
  NOR2_X1   g697(.A1(new_n673), .A2(new_n492), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n688), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n857), .A2(new_n254), .A3(new_n863), .A4(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(KEYINPUT124), .B(G197gat), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n856), .A2(new_n900), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n711), .A3(new_n903), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT125), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n905), .A2(new_n910), .A3(new_n907), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(G1352gat));
  INV_X1    g711(.A(G204gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n906), .A2(new_n913), .A3(new_n666), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n914), .A2(KEYINPUT62), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n857), .A2(new_n666), .A3(new_n863), .ZN(new_n916));
  OAI21_X1  g715(.A(G204gat), .B1(new_n916), .B2(new_n900), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n914), .A2(KEYINPUT62), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(G1353gat));
  NAND3_X1  g718(.A1(new_n906), .A2(new_n268), .A3(new_n614), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n857), .A2(new_n614), .A3(new_n863), .A4(new_n901), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT63), .B1(new_n921), .B2(G211gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(G1354gat));
  NOR2_X1   g723(.A1(new_n644), .A2(new_n269), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n857), .A2(new_n863), .A3(new_n901), .A4(new_n925), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n824), .A2(new_n362), .A3(new_n643), .A4(new_n901), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n927), .A2(KEYINPUT126), .A3(new_n269), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT126), .B1(new_n927), .B2(new_n269), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n930), .B(new_n931), .ZN(G1355gat));
endmodule


