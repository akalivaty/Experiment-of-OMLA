//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1325, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  AOI211_X1 g0011(.A(new_n206), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n201), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n212), .A2(KEYINPUT0), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT64), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G68), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G87), .A2(G250), .ZN(new_n230));
  NAND4_X1  g0030(.A1(new_n227), .A2(new_n228), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n207), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT1), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n219), .B(new_n233), .C1(KEYINPUT0), .C2(new_n212), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT65), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G58), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND2_X1  g0050(.A1(new_n203), .A2(G20), .ZN(new_n251));
  INV_X1    g0051(.A(G150), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n214), .A2(G33), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n251), .B1(new_n252), .B2(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n213), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G50), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n259), .B1(new_n261), .B2(G20), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n263), .B1(new_n264), .B2(G50), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT9), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n260), .A2(KEYINPUT9), .A3(new_n265), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT68), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n271), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n272), .A2(G33), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT68), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(G222), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(G223), .A3(G1698), .ZN(new_n283));
  INV_X1    g0083(.A(G77), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n282), .B(new_n283), .C1(new_n284), .C2(new_n280), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(G1), .A3(G13), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G45), .ZN(new_n290));
  NAND2_X1  g0090(.A1(KEYINPUT66), .A2(G41), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(KEYINPUT66), .A2(G41), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n290), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G274), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(G1), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G226), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n287), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n297), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT67), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n289), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n270), .B1(new_n304), .B2(G190), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT73), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n303), .B2(G200), .ZN(new_n307));
  INV_X1    g0107(.A(G200), .ZN(new_n308));
  AOI211_X1 g0108(.A(KEYINPUT73), .B(new_n308), .C1(new_n289), .C2(new_n302), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n305), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n305), .B(new_n312), .C1(new_n307), .C2(new_n309), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT69), .B(G179), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n304), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n266), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n318), .B1(new_n303), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n314), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(KEYINPUT75), .A2(G169), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT13), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT68), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT68), .B1(new_n277), .B2(new_n278), .ZN(new_n327));
  OAI211_X1 g0127(.A(G232), .B(G1698), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  OAI211_X1 g0128(.A(G226), .B(new_n281), .C1(new_n326), .C2(new_n327), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G97), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n288), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n297), .B1(new_n225), .B2(new_n300), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n325), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  AOI211_X1 g0135(.A(KEYINPUT13), .B(new_n333), .C1(new_n331), .C2(new_n288), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n324), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT14), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n332), .A2(new_n334), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT13), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n332), .A2(new_n325), .A3(new_n334), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT14), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n343), .A3(new_n324), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n335), .A2(new_n336), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT76), .B1(new_n345), .B2(G179), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT76), .ZN(new_n347));
  INV_X1    g0147(.A(G179), .ZN(new_n348));
  NOR4_X1   g0148(.A1(new_n335), .A2(new_n336), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n338), .B(new_n344), .C1(new_n346), .C2(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT64), .B(G68), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n351), .A2(new_n214), .B1(new_n284), .B2(new_n255), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(KEYINPUT74), .B1(G50), .B2(new_n253), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(KEYINPUT74), .B2(new_n352), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n259), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT11), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT12), .ZN(new_n358));
  OAI21_X1  g0158(.A(G68), .B1(new_n264), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n262), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n224), .A2(new_n360), .A3(KEYINPUT12), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n359), .B(new_n361), .C1(KEYINPUT12), .C2(new_n360), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n350), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n345), .A2(G190), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n342), .A2(G200), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n363), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G159), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n254), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G58), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n217), .B1(new_n224), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n372), .B1(new_n374), .B2(G20), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  AOI211_X1 g0176(.A(new_n376), .B(G20), .C1(new_n277), .C2(new_n278), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n276), .A2(new_n214), .A3(new_n279), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n377), .B1(new_n378), .B2(new_n376), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n375), .B1(new_n379), .B2(new_n224), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT16), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n277), .A2(new_n278), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT7), .B1(new_n383), .B2(new_n214), .ZN(new_n384));
  OAI21_X1  g0184(.A(G68), .B1(new_n384), .B2(new_n377), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(new_n375), .A3(KEYINPUT16), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n386), .A2(new_n259), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT78), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n287), .A2(G232), .A3(new_n299), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT66), .ZN(new_n391));
  INV_X1    g0191(.A(G41), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(G45), .B1(new_n393), .B2(new_n291), .ZN(new_n394));
  INV_X1    g0194(.A(new_n296), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n390), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  OR2_X1    g0197(.A1(G223), .A2(G1698), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n298), .A2(G1698), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n277), .A2(new_n398), .A3(new_n278), .A4(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G87), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n288), .ZN(new_n403));
  AOI21_X1  g0203(.A(G200), .B1(new_n397), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n287), .B1(new_n400), .B2(new_n401), .ZN(new_n405));
  NOR3_X1   g0205(.A1(new_n405), .A2(new_n396), .A3(G190), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n389), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n308), .B1(new_n405), .B2(new_n396), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n397), .A2(new_n403), .ZN(new_n409));
  OAI211_X1 g0209(.A(KEYINPUT78), .B(new_n408), .C1(new_n409), .C2(G190), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n256), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(new_n360), .ZN(new_n413));
  INV_X1    g0213(.A(new_n264), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n413), .B1(new_n414), .B2(new_n412), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n388), .A2(new_n411), .A3(KEYINPUT79), .A4(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n415), .B1(new_n382), .B2(new_n387), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n420), .A2(KEYINPUT79), .A3(KEYINPUT17), .A4(new_n411), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n397), .A2(new_n403), .A3(new_n315), .ZN(new_n422));
  OAI21_X1  g0222(.A(G169), .B1(new_n405), .B2(new_n396), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT77), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n422), .A2(KEYINPUT77), .A3(new_n423), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT18), .B1(new_n420), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n426), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(new_n424), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT18), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n386), .A2(new_n259), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n381), .B2(new_n380), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n430), .B(new_n431), .C1(new_n433), .C2(new_n415), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n419), .A2(new_n421), .A3(new_n428), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n259), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n412), .A2(KEYINPUT71), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT71), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n256), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n253), .A3(new_n439), .ZN(new_n440));
  XOR2_X1   g0240(.A(KEYINPUT15), .B(G87), .Z(new_n441));
  INV_X1    g0241(.A(new_n255), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n441), .A2(new_n442), .B1(G20), .B2(G77), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n436), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT72), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n360), .A2(new_n284), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n414), .B2(new_n284), .ZN(new_n447));
  OR3_X1    g0247(.A1(new_n444), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n445), .B1(new_n444), .B2(new_n447), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n280), .A2(G232), .A3(new_n281), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n280), .A2(G238), .A3(G1698), .ZN(new_n453));
  INV_X1    g0253(.A(G107), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n452), .B(new_n453), .C1(new_n454), .C2(new_n280), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n288), .ZN(new_n456));
  INV_X1    g0256(.A(G244), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n297), .B1(new_n457), .B2(new_n300), .ZN(new_n458));
  XNOR2_X1  g0258(.A(new_n458), .B(KEYINPUT70), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G190), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n451), .B(new_n461), .C1(new_n308), .C2(new_n460), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n456), .A2(new_n459), .A3(new_n316), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n450), .B(new_n463), .C1(new_n460), .C2(G169), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NOR4_X1   g0265(.A1(new_n322), .A2(new_n370), .A3(new_n435), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n261), .A2(G33), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n262), .A2(new_n467), .A3(new_n213), .A4(new_n258), .ZN(new_n468));
  INV_X1    g0268(.A(G116), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(KEYINPUT86), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT86), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n468), .A2(new_n472), .A3(new_n469), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n360), .A2(new_n469), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G283), .ZN(new_n476));
  INV_X1    g0276(.A(G97), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n476), .B(new_n214), .C1(G33), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n469), .A2(G20), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n478), .A2(new_n259), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT20), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n480), .A2(new_n481), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n475), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n474), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT5), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n261), .B(G45), .C1(new_n486), .C2(G41), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n393), .A2(new_n486), .A3(new_n291), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n288), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G270), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n488), .A2(new_n489), .A3(G274), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n276), .A2(G303), .A3(new_n279), .ZN(new_n494));
  XNOR2_X1  g0294(.A(KEYINPUT3), .B(G33), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n211), .A2(G1698), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n495), .B(new_n496), .C1(G257), .C2(G1698), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n287), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(G169), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n485), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT21), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n493), .A2(new_n498), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G190), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n503), .B(new_n485), .C1(new_n308), .C2(new_n502), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT21), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n485), .B2(new_n499), .ZN(new_n506));
  INV_X1    g0306(.A(new_n485), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n493), .A2(new_n498), .A3(new_n348), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n501), .A2(new_n504), .A3(new_n506), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT87), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n500), .A2(KEYINPUT21), .B1(new_n507), .B2(new_n508), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT87), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n512), .A2(new_n513), .A3(new_n506), .A4(new_n504), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n225), .A2(new_n281), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n457), .A2(G1698), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n277), .A2(new_n516), .A3(new_n278), .A4(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n274), .A2(new_n469), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n287), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n261), .A2(G45), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G250), .ZN(new_n523));
  OAI22_X1  g0323(.A1(new_n288), .A2(new_n523), .B1(new_n295), .B2(new_n522), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT83), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n522), .A2(new_n295), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n206), .B1(new_n261), .B2(G45), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n526), .B1(new_n287), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT83), .ZN(new_n529));
  NOR2_X1   g0329(.A1(G238), .A2(G1698), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n530), .B1(new_n457), .B2(G1698), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n519), .B1(new_n531), .B2(new_n495), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n528), .B(new_n529), .C1(new_n532), .C2(new_n287), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n525), .A2(new_n533), .A3(new_n319), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n315), .B1(new_n525), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT84), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n525), .A2(new_n533), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n316), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT84), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n525), .A2(new_n533), .A3(new_n319), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n495), .A2(new_n214), .A3(G68), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT19), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n214), .B1(new_n330), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(G87), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n545), .A2(new_n477), .A3(new_n454), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n543), .B1(new_n255), .B2(new_n477), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n542), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n441), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n549), .A2(new_n259), .B1(new_n360), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n468), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n441), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n536), .A2(new_n541), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n549), .A2(new_n259), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(G87), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n550), .A2(new_n360), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(G190), .B2(new_n537), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n308), .B2(new_n537), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n555), .A2(KEYINPUT85), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT85), .B1(new_n555), .B2(new_n561), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(G250), .B(G1698), .C1(new_n326), .C2(new_n327), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT4), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n566), .A2(new_n457), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n281), .B(new_n567), .C1(new_n326), .C2(new_n327), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n457), .A2(G1698), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n570), .A2(new_n277), .A3(new_n278), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT82), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n572), .A3(new_n566), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n572), .B1(new_n571), .B2(new_n566), .ZN(new_n575));
  INV_X1    g0375(.A(new_n476), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n287), .B1(new_n569), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n490), .A2(G257), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n492), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n319), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n575), .A2(new_n576), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n582), .A2(new_n573), .A3(new_n565), .A4(new_n568), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n288), .ZN(new_n584));
  INV_X1    g0384(.A(new_n580), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n316), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n378), .A2(new_n376), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n383), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n254), .A2(new_n284), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n477), .A2(new_n454), .A3(KEYINPUT6), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT6), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G97), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n454), .A2(KEYINPUT80), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT80), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G107), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n591), .A2(new_n593), .A3(new_n595), .A4(new_n597), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n590), .B1(new_n601), .B2(G20), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT81), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n589), .A2(G107), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n214), .B1(new_n599), .B2(new_n600), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT81), .B1(new_n605), .B2(new_n590), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n436), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n360), .A2(new_n477), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n468), .B2(new_n477), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n581), .B(new_n586), .C1(new_n607), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n584), .A2(new_n585), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(G200), .ZN(new_n612));
  INV_X1    g0412(.A(new_n600), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n591), .A2(new_n593), .B1(new_n595), .B2(new_n597), .ZN(new_n614));
  OAI21_X1  g0414(.A(G20), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n590), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n603), .A3(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n617), .B(new_n606), .C1(new_n454), .C2(new_n379), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n609), .B1(new_n618), .B2(new_n259), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n584), .A2(G190), .A3(new_n585), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n612), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT24), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n454), .A2(G20), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT88), .B1(new_n623), .B2(KEYINPUT23), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT88), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT23), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n625), .A2(new_n626), .A3(new_n454), .A4(G20), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n624), .A2(new_n627), .B1(KEYINPUT23), .B2(new_n623), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT22), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(new_n545), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n519), .B1(new_n495), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n628), .B1(new_n631), .B2(G20), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n545), .A2(G20), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT22), .B1(new_n280), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n622), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n326), .A2(new_n327), .ZN(new_n636));
  INV_X1    g0436(.A(new_n633), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n629), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n631), .A2(G20), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n638), .A2(new_n639), .A3(KEYINPUT24), .A4(new_n628), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n635), .A2(new_n640), .A3(new_n259), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n360), .A2(KEYINPUT25), .A3(new_n454), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n642), .A2(KEYINPUT89), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT25), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(new_n262), .B2(G107), .ZN(new_n645));
  OAI22_X1  g0445(.A1(new_n643), .A2(new_n645), .B1(new_n454), .B2(new_n468), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n643), .B2(new_n645), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n210), .A2(G1698), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(G250), .B2(G1698), .ZN(new_n650));
  INV_X1    g0450(.A(G294), .ZN(new_n651));
  OAI22_X1  g0451(.A1(new_n650), .A2(new_n383), .B1(new_n274), .B2(new_n651), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n490), .A2(G264), .B1(new_n652), .B2(new_n288), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n653), .A2(G179), .A3(new_n492), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n319), .B1(new_n653), .B2(new_n492), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT90), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n656), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT90), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(new_n654), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n648), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n653), .A2(G190), .A3(new_n492), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n653), .A2(new_n492), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G200), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n641), .A2(new_n647), .A3(new_n662), .A4(new_n664), .ZN(new_n665));
  AND4_X1   g0465(.A1(new_n610), .A2(new_n621), .A3(new_n661), .A4(new_n665), .ZN(new_n666));
  AND4_X1   g0466(.A1(new_n466), .A2(new_n515), .A3(new_n564), .A4(new_n666), .ZN(G372));
  NAND2_X1  g0467(.A1(new_n419), .A2(new_n421), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n368), .A2(new_n464), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n668), .B1(new_n669), .B2(new_n365), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n388), .A2(new_n416), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n422), .A2(new_n423), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT18), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n672), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n420), .A2(new_n431), .A3(new_n674), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n314), .B1(new_n670), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n321), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(G169), .B1(new_n584), .B2(new_n585), .ZN(new_n681));
  AOI211_X1 g0481(.A(new_n315), .B(new_n580), .C1(new_n583), .C2(new_n288), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n528), .B1(new_n532), .B2(new_n287), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G200), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n551), .A2(new_n553), .B1(new_n319), .B2(new_n684), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n560), .A2(new_n685), .B1(new_n538), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n618), .A2(new_n259), .ZN(new_n688));
  INV_X1    g0488(.A(new_n609), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT26), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n683), .A2(new_n687), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n538), .A2(new_n686), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AND4_X1   g0494(.A1(new_n610), .A2(new_n621), .A3(new_n665), .A4(new_n687), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n648), .B1(new_n656), .B2(new_n655), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(new_n512), .A3(new_n506), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n694), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n555), .A2(new_n561), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT85), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n555), .A2(KEYINPUT85), .A3(new_n561), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n619), .A2(new_n681), .A3(new_n682), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT26), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n698), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n466), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n680), .A2(new_n707), .ZN(G369));
  INV_X1    g0508(.A(G13), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G20), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n261), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n711), .A2(KEYINPUT27), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(KEYINPUT27), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G213), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(G343), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n515), .B1(new_n485), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n512), .A2(new_n506), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(new_n507), .A3(new_n716), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(G330), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n661), .A2(new_n665), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n648), .A2(new_n716), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n661), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n716), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n724), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n719), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n716), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n725), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n696), .A2(new_n716), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n731), .A2(new_n737), .ZN(G399));
  NAND2_X1  g0538(.A1(new_n393), .A2(new_n291), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n209), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n546), .A2(G116), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n742), .A2(G1), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(new_n218), .B2(new_n742), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT91), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT28), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n716), .B1(new_n698), .B2(new_n705), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT29), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n701), .A2(new_n691), .A3(new_n702), .A4(new_n703), .ZN(new_n751));
  INV_X1    g0551(.A(new_n693), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n703), .A2(new_n687), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n752), .B1(new_n753), .B2(KEYINPUT26), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT92), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n732), .A2(new_n661), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n755), .A2(new_n756), .B1(new_n695), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n751), .A2(new_n754), .A3(KEYINPUT92), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n716), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n750), .B1(new_n760), .B2(new_n749), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n578), .A2(new_n580), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n763), .A2(new_n508), .A3(new_n537), .A4(new_n653), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT30), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n663), .A2(new_n316), .A3(new_n684), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n502), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n764), .A2(new_n765), .B1(new_n611), .B2(new_n768), .ZN(new_n769));
  AOI211_X1 g0569(.A(KEYINPUT31), .B(new_n717), .C1(new_n766), .C2(new_n769), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n515), .A2(new_n564), .A3(new_n666), .A4(new_n717), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT31), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n766), .A2(new_n769), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n772), .B1(new_n773), .B2(new_n716), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n770), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G330), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n762), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n747), .B1(new_n778), .B2(G1), .ZN(G364));
  AOI21_X1  g0579(.A(new_n261), .B1(new_n710), .B2(G45), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n741), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n724), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(G330), .B2(new_n721), .ZN(new_n784));
  INV_X1    g0584(.A(new_n782), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n280), .A2(G355), .A3(new_n208), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n249), .A2(new_n290), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n209), .A2(new_n495), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(G45), .B2(new_n218), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n786), .B1(G116), .B2(new_n208), .C1(new_n787), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n213), .B1(G20), .B2(new_n319), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n785), .B1(new_n790), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n794), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n315), .A2(G20), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G190), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G200), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n798), .A2(new_n800), .A3(new_n308), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n803), .A2(G322), .B1(G326), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G329), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n214), .A2(G179), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G190), .A2(G200), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT96), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n805), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n800), .A2(new_n308), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n807), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n308), .A2(G190), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n807), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G303), .A2(new_n814), .B1(new_n817), .B2(G283), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n801), .A2(new_n348), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(G20), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n818), .B(new_n636), .C1(new_n651), .C2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(G311), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n799), .A2(new_n808), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n799), .A2(new_n815), .ZN(new_n825));
  XOR2_X1   g0625(.A(KEYINPUT33), .B(G317), .Z(new_n826));
  OAI22_X1  g0626(.A1(new_n823), .A2(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n811), .A2(new_n822), .A3(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n804), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n829), .A2(new_n202), .B1(new_n373), .B2(new_n802), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n824), .A2(KEYINPUT93), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n798), .A2(G190), .A3(G200), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT93), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n830), .B1(new_n836), .B2(G77), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(KEYINPUT94), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n813), .A2(new_n545), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n839), .B(new_n636), .C1(G107), .C2(new_n817), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n840), .B1(new_n220), .B2(new_n825), .C1(new_n477), .C2(new_n821), .ZN(new_n841));
  INV_X1    g0641(.A(new_n809), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(G159), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT95), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT32), .Z(new_n845));
  NOR3_X1   g0645(.A1(new_n838), .A2(new_n841), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n837), .A2(KEYINPUT94), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n828), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n793), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n796), .B1(new_n797), .B2(new_n848), .C1(new_n721), .C2(new_n849), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n784), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(G396));
  NAND2_X1  g0652(.A1(new_n836), .A2(G116), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n813), .A2(new_n454), .B1(new_n816), .B2(new_n545), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n280), .B(new_n854), .C1(G97), .C2(new_n820), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n803), .A2(G294), .B1(G303), .B2(new_n804), .ZN(new_n856));
  INV_X1    g0656(.A(new_n810), .ZN(new_n857));
  INV_X1    g0657(.A(new_n825), .ZN(new_n858));
  AOI22_X1  g0658(.A1(G311), .A2(new_n857), .B1(new_n858), .B2(G283), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n853), .A2(new_n855), .A3(new_n856), .A4(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n803), .A2(G143), .B1(G137), .B2(new_n804), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n252), .B2(new_n825), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(G159), .B2(new_n836), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT34), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n816), .A2(new_n220), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(G50), .B2(new_n814), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n373), .B2(new_n821), .ZN(new_n867));
  INV_X1    g0667(.A(G132), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n495), .B1(new_n810), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n867), .B1(new_n869), .B2(KEYINPUT97), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n864), .B(new_n870), .C1(KEYINPUT97), .C2(new_n869), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n863), .A2(KEYINPUT34), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n860), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT98), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n875), .A2(new_n876), .A3(new_n797), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n794), .A2(new_n791), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n782), .B1(G77), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n882), .A2(KEYINPUT99), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(KEYINPUT99), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n464), .A2(new_n716), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n462), .B1(new_n451), .B2(new_n717), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n885), .B1(new_n886), .B2(new_n464), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n887), .A2(new_n792), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n883), .A2(new_n884), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n748), .B(new_n887), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n890), .A2(new_n776), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n782), .B1(new_n890), .B2(new_n776), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(G384));
  INV_X1    g0695(.A(KEYINPUT104), .ZN(new_n896));
  INV_X1    g0696(.A(new_n714), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n676), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n368), .B1(new_n350), .B2(new_n364), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n364), .A2(new_n716), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n346), .A2(new_n349), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n344), .A2(new_n338), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n363), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n899), .A2(new_n900), .B1(new_n903), .B2(new_n716), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n691), .B1(new_n564), .B2(new_n703), .ZN(new_n905));
  INV_X1    g0705(.A(new_n694), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n687), .A2(new_n665), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n697), .A2(new_n907), .A3(new_n610), .A4(new_n621), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n717), .B(new_n887), .C1(new_n905), .C2(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n885), .B(KEYINPUT100), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n904), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT38), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT37), .B1(new_n420), .B2(new_n411), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n671), .A2(new_n430), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n897), .B1(new_n433), .B2(new_n415), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n386), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n385), .A2(new_n375), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n436), .B1(new_n919), .B2(new_n381), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n918), .B1(new_n920), .B2(KEYINPUT101), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT101), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT16), .B1(new_n385), .B2(new_n375), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n922), .B1(new_n923), .B2(new_n436), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n415), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT102), .B1(new_n925), .B2(new_n714), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n201), .B1(new_n351), .B2(G58), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n927), .A2(new_n214), .B1(new_n371), .B2(new_n254), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n376), .B1(new_n495), .B2(G20), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n220), .B1(new_n929), .B2(new_n588), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n381), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(KEYINPUT101), .A3(new_n259), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n924), .A2(new_n386), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n416), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n934), .A2(new_n672), .B1(new_n420), .B2(new_n411), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT102), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n934), .A2(new_n936), .A3(new_n897), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n926), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n917), .B1(new_n938), .B2(KEYINPUT37), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n926), .A2(new_n937), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n940), .A2(new_n435), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n913), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n435), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT37), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n936), .B1(new_n934), .B2(new_n897), .ZN(new_n945));
  AOI211_X1 g0745(.A(KEYINPUT102), .B(new_n714), .C1(new_n933), .C2(new_n416), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n944), .B1(new_n947), .B2(new_n935), .ZN(new_n948));
  OAI211_X1 g0748(.A(KEYINPUT38), .B(new_n943), .C1(new_n948), .C2(new_n917), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n942), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n898), .B1(new_n912), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n903), .A2(new_n717), .ZN(new_n953));
  INV_X1    g0753(.A(new_n916), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n421), .B(new_n419), .C1(new_n673), .C2(new_n675), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n672), .B1(new_n433), .B2(new_n415), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n420), .A2(new_n411), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n956), .A2(new_n916), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT37), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n954), .A2(new_n955), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT103), .B1(new_n961), .B2(KEYINPUT38), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(new_n942), .A3(new_n949), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT39), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n955), .A2(new_n954), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n959), .A2(new_n960), .ZN(new_n966));
  AOI21_X1  g0766(.A(KEYINPUT38), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n938), .A2(KEYINPUT37), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n968), .A2(new_n960), .B1(new_n435), .B2(new_n940), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n967), .B1(new_n969), .B2(KEYINPUT38), .ZN(new_n970));
  NOR2_X1   g0770(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n953), .B1(new_n964), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n896), .B1(new_n952), .B2(new_n973), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n963), .A2(KEYINPUT39), .B1(new_n970), .B2(new_n971), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n951), .B(KEYINPUT104), .C1(new_n975), .C2(new_n953), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n679), .B1(new_n761), .B2(new_n466), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT40), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n942), .A2(new_n949), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n365), .A2(new_n369), .A3(new_n900), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n365), .B2(new_n717), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n983), .A2(new_n775), .A3(new_n887), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n980), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  AND3_X1   g0785(.A1(new_n983), .A2(new_n775), .A3(new_n887), .ZN(new_n986));
  INV_X1    g0786(.A(new_n967), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n980), .B1(new_n987), .B2(new_n949), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n985), .A2(G330), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n466), .A2(G330), .A3(new_n775), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n950), .A2(new_n775), .A3(new_n887), .A4(new_n983), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n993), .A2(new_n980), .B1(new_n986), .B2(new_n988), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n994), .A2(new_n466), .A3(new_n775), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n979), .A2(new_n996), .B1(new_n261), .B2(new_n710), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT105), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n979), .A2(new_n996), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n997), .A2(new_n998), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n601), .A2(KEYINPUT35), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1003), .A2(G116), .A3(new_n215), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(KEYINPUT35), .B2(new_n601), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(KEYINPUT36), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1005), .A2(KEYINPUT36), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n284), .B(new_n218), .C1(new_n351), .C2(G58), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n220), .A2(G50), .ZN(new_n1009));
  OAI211_X1 g0809(.A(G1), .B(new_n709), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1002), .A2(new_n1006), .A3(new_n1007), .A4(new_n1010), .ZN(G367));
  INV_X1    g0811(.A(new_n788), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n241), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n795), .B1(new_n208), .B2(new_n550), .ZN(new_n1014));
  INV_X1    g0814(.A(G143), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n829), .A2(new_n1015), .B1(new_n371), .B2(new_n825), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G150), .B2(new_n803), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n836), .A2(G50), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n813), .A2(new_n373), .B1(new_n816), .B2(new_n284), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G137), .B2(new_n842), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n820), .A2(G68), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1021), .A2(new_n280), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n817), .A2(G97), .ZN(new_n1024));
  INV_X1    g0824(.A(G317), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1024), .B(new_n383), .C1(new_n1025), .C2(new_n809), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G107), .B2(new_n820), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n803), .A2(G303), .B1(G311), .B2(new_n804), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT110), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT46), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n813), .B2(new_n469), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n814), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(new_n825), .C2(new_n651), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1027), .B(new_n1028), .C1(new_n1029), .C2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1029), .ZN(new_n1035));
  INV_X1    g0835(.A(G283), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1035), .B1(new_n835), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1023), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT47), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n794), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n782), .B1(new_n1013), .B2(new_n1014), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT111), .Z(new_n1043));
  NAND2_X1  g0843(.A1(new_n559), .A2(new_n716), .ZN(new_n1044));
  MUX2_X1   g0844(.A(new_n752), .B(new_n687), .S(new_n1044), .Z(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT106), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n793), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT112), .Z(new_n1049));
  OAI211_X1 g0849(.A(new_n610), .B(new_n621), .C1(new_n619), .C2(new_n717), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n610), .B2(new_n717), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT107), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n735), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT42), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n728), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n716), .B1(new_n1055), .B2(new_n610), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT43), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n1058), .A3(new_n1046), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n731), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1046), .A2(new_n1058), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1046), .A2(new_n1058), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(new_n1054), .C2(new_n1056), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1059), .A2(new_n1060), .A3(new_n1052), .A4(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT108), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1059), .A2(new_n1063), .B1(new_n1060), .B2(new_n1052), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT45), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1051), .A2(KEYINPUT107), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1051), .A2(KEYINPUT107), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n734), .B1(new_n696), .B2(new_n716), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1070), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1052), .A2(new_n737), .A3(KEYINPUT45), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT44), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n1052), .B2(new_n737), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1073), .A2(KEYINPUT44), .A3(new_n1074), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n1060), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1077), .A2(new_n1081), .A3(new_n731), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT109), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n722), .B2(new_n723), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n734), .B1(new_n730), .B2(new_n733), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1087), .B(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n778), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n741), .B(KEYINPUT41), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n780), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1049), .B1(new_n1069), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(G387));
  NAND2_X1  g0896(.A1(new_n778), .A2(new_n1089), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1097), .A2(KEYINPUT117), .A3(new_n741), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT117), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1090), .A2(new_n777), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n742), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1098), .B(new_n1101), .C1(new_n778), .C2(new_n1089), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n727), .A2(new_n729), .A3(new_n793), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n238), .A2(G45), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1105), .A2(KEYINPUT113), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(KEYINPUT113), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n437), .A2(new_n439), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1108), .A2(G50), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n1110), .A2(KEYINPUT50), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(KEYINPUT50), .ZN(new_n1112));
  AOI21_X1  g0912(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1111), .A2(new_n743), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1106), .A2(new_n788), .A3(new_n1107), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n280), .A2(new_n208), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1115), .B1(G107), .B2(new_n208), .C1(new_n743), .C2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n785), .B1(new_n1117), .B2(new_n795), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n814), .A2(G77), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n842), .A2(G150), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1119), .A2(new_n1024), .A3(new_n1120), .A4(new_n495), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n858), .A2(new_n412), .B1(G159), .B2(new_n804), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n202), .B2(new_n802), .C1(new_n220), .C2(new_n824), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1121), .B(new_n1123), .C1(new_n441), .C2(new_n820), .ZN(new_n1124));
  INV_X1    g0924(.A(G303), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n835), .A2(new_n1125), .B1(new_n1025), .B2(new_n802), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT114), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n858), .A2(G311), .B1(G322), .B2(new_n804), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT115), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT48), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT115), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1129), .B(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(KEYINPUT48), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G283), .A2(new_n820), .B1(new_n814), .B2(G294), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1132), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT49), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n495), .B1(new_n842), .B2(G326), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n469), .B2(new_n816), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1124), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1103), .B(new_n1118), .C1(new_n1143), .C2(new_n797), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT116), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1090), .A2(new_n780), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1102), .A2(new_n1147), .ZN(G393));
  NOR2_X1   g0948(.A1(new_n246), .A2(new_n1012), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n795), .B1(new_n477), .B2(new_n208), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n782), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n803), .A2(G159), .B1(G150), .B2(new_n804), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT51), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n821), .A2(new_n284), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n495), .B1(new_n816), .B2(new_n545), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n813), .A2(new_n224), .B1(new_n809), .B2(new_n1015), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n202), .B2(new_n825), .C1(new_n835), .C2(new_n1108), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1153), .A2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT120), .Z(new_n1160));
  OAI22_X1  g0960(.A1(new_n829), .A2(new_n1025), .B1(new_n823), .B2(new_n802), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT52), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G107), .A2(new_n817), .B1(new_n842), .B2(G322), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n1036), .B2(new_n813), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n280), .B(new_n1164), .C1(G116), .C2(new_n820), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n858), .A2(G303), .B1(G294), .B2(new_n832), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1162), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(KEYINPUT121), .B1(new_n1160), .B2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1168), .A2(new_n797), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1160), .A2(KEYINPUT121), .A3(new_n1167), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1151), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n1052), .B2(new_n849), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT119), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1083), .B(new_n1173), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1084), .B(KEYINPUT118), .Z(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1100), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n741), .B1(new_n1097), .B2(new_n1085), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1172), .B1(new_n1176), .B2(new_n780), .C1(new_n1177), .C2(new_n1178), .ZN(G390));
  NAND4_X1  g0979(.A1(new_n983), .A2(new_n775), .A3(G330), .A4(new_n887), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n911), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n748), .B2(new_n887), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n953), .B1(new_n1183), .B2(new_n904), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1184), .A2(new_n964), .A3(new_n972), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n987), .A2(new_n949), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n953), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n755), .A2(new_n756), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n757), .A2(new_n695), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(new_n759), .A3(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(new_n717), .A3(new_n887), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n911), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1187), .B1(new_n1192), .B2(new_n983), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1181), .B1(new_n1185), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1187), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1182), .B1(new_n760), .B2(new_n887), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1195), .B1(new_n1196), .B2(new_n904), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n975), .A2(new_n1184), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1197), .A2(new_n1198), .A3(new_n1180), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1194), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n761), .A2(new_n466), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1201), .A2(new_n680), .A3(new_n991), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n887), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n904), .B1(new_n776), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n1180), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1183), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1196), .A2(new_n1180), .A3(new_n1204), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1202), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1200), .A2(new_n1210), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1194), .A2(new_n1199), .A3(new_n1202), .A4(new_n1209), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1211), .A2(new_n741), .A3(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1194), .A2(new_n781), .A3(new_n1199), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n782), .B1(new_n412), .B2(new_n879), .ZN(new_n1215));
  INV_X1    g1015(.A(G137), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n825), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n814), .A2(G150), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT53), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1217), .B(new_n1219), .C1(G128), .C2(new_n804), .ZN(new_n1220));
  XOR2_X1   g1020(.A(KEYINPUT54), .B(G143), .Z(new_n1221));
  NAND2_X1  g1021(.A1(new_n836), .A2(new_n1221), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n280), .B1(new_n202), .B2(new_n816), .C1(new_n821), .C2(new_n371), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G125), .A2(new_n857), .B1(new_n803), .B2(G132), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1220), .A2(new_n1222), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n835), .A2(new_n477), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(G107), .A2(new_n858), .B1(new_n803), .B2(G116), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(new_n1154), .A2(new_n280), .A3(new_n839), .A4(new_n865), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n857), .A2(G294), .B1(G283), .B2(new_n804), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1226), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1215), .B1(new_n1232), .B2(new_n794), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n964), .A2(new_n972), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1233), .B1(new_n1234), .B2(new_n792), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1214), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1213), .A2(new_n1236), .ZN(G378));
  NOR2_X1   g1037(.A1(new_n318), .A2(new_n714), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n322), .A2(new_n1238), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n314), .B(new_n321), .C1(new_n318), .C2(new_n714), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1241), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1239), .A2(new_n1240), .A3(new_n1242), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n994), .A2(G330), .A3(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1246), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n990), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n953), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1234), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT104), .B1(new_n1251), .B2(new_n951), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n976), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1247), .B(new_n1249), .C1(new_n1252), .C2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1246), .B1(new_n994), .B2(G330), .ZN(new_n1255));
  AND4_X1   g1055(.A1(G330), .A2(new_n985), .A3(new_n989), .A4(new_n1246), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n974), .B(new_n976), .C1(new_n1255), .C2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1254), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n781), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n803), .A2(G128), .B1(new_n814), .B2(new_n1221), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT122), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(G125), .A2(new_n804), .B1(new_n832), .B2(G137), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n1262), .B1(new_n868), .B2(new_n825), .C1(new_n252), .C2(new_n821), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  XOR2_X1   g1064(.A(new_n1264), .B(KEYINPUT59), .Z(new_n1265));
  AOI211_X1 g1065(.A(G33), .B(G41), .C1(new_n842), .C2(G124), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n371), .B2(new_n816), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(G283), .A2(new_n857), .B1(new_n803), .B2(G107), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n550), .B2(new_n824), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n817), .A2(G58), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n740), .A2(new_n495), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1021), .A2(new_n1119), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n829), .A2(new_n469), .B1(new_n477), .B2(new_n825), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1270), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1275), .A2(KEYINPUT58), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(KEYINPUT58), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1276), .B(new_n1277), .C1(new_n1272), .C2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n794), .B1(new_n1268), .B2(new_n1279), .ZN(new_n1280));
  XOR2_X1   g1080(.A(new_n1280), .B(KEYINPUT123), .Z(new_n1281));
  OAI21_X1  g1081(.A(new_n782), .B1(G50), .B2(new_n879), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1282), .B(KEYINPUT124), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1281), .B(new_n1283), .C1(new_n792), .C2(new_n1246), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1259), .A2(new_n1284), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n1254), .A2(new_n1257), .B1(new_n1212), .B2(new_n1202), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n741), .B1(new_n1286), .B2(KEYINPUT57), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT57), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(new_n1212), .B2(new_n1202), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1254), .A2(KEYINPUT125), .A3(new_n1257), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT125), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n977), .A2(new_n1291), .A3(new_n1247), .A4(new_n1249), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1289), .A2(new_n1290), .A3(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1285), .B1(new_n1287), .B2(new_n1293), .ZN(G375));
  AOI22_X1  g1094(.A1(G97), .A2(new_n814), .B1(new_n817), .B2(G77), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1295), .B(new_n636), .C1(new_n550), .C2(new_n821), .ZN(new_n1296));
  AOI22_X1  g1096(.A1(new_n858), .A2(G116), .B1(G294), .B2(new_n804), .ZN(new_n1297));
  OAI221_X1 g1097(.A(new_n1297), .B1(new_n1036), .B2(new_n802), .C1(new_n1125), .C2(new_n810), .ZN(new_n1298));
  AOI211_X1 g1098(.A(new_n1296), .B(new_n1298), .C1(G107), .C2(new_n836), .ZN(new_n1299));
  AOI22_X1  g1099(.A1(new_n858), .A2(new_n1221), .B1(G132), .B2(new_n804), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1300), .B1(new_n252), .B2(new_n824), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n383), .B1(new_n817), .B2(G58), .ZN(new_n1302));
  OAI221_X1 g1102(.A(new_n1302), .B1(new_n371), .B2(new_n813), .C1(new_n202), .C2(new_n821), .ZN(new_n1303));
  INV_X1    g1103(.A(G128), .ZN(new_n1304));
  OAI22_X1  g1104(.A1(new_n810), .A2(new_n1304), .B1(new_n802), .B2(new_n1216), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1301), .A2(new_n1303), .A3(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n794), .B1(new_n1299), .B2(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1307), .B(new_n782), .C1(G68), .C2(new_n879), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1308), .B1(new_n904), .B2(new_n791), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1309), .B1(new_n1209), .B2(new_n781), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1210), .A2(new_n1092), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1202), .A2(new_n1209), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1310), .B1(new_n1311), .B2(new_n1312), .ZN(G381));
  NOR4_X1   g1113(.A1(G387), .A2(G384), .A3(G390), .A4(G381), .ZN(new_n1314));
  INV_X1    g1114(.A(G378), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1259), .A2(new_n1284), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1212), .A2(new_n1202), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1258), .A2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n742), .B1(new_n1318), .B2(new_n1288), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1289), .A2(new_n1290), .A3(new_n1292), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1316), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1102), .A2(new_n851), .A3(new_n1147), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1314), .A2(new_n1315), .A3(new_n1321), .A4(new_n1323), .ZN(G407));
  NAND2_X1  g1124(.A1(new_n1321), .A2(new_n1315), .ZN(new_n1325));
  OAI211_X1 g1125(.A(G407), .B(G213), .C1(G343), .C2(new_n1325), .ZN(G409));
  NAND3_X1  g1126(.A1(new_n1290), .A2(new_n781), .A3(new_n1292), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1258), .A2(new_n1317), .A3(new_n1092), .ZN(new_n1328));
  AND2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1213), .A2(new_n1236), .A3(new_n1284), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(G213), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1332), .A2(G343), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  OAI211_X1 g1134(.A(new_n1331), .B(new_n1334), .C1(new_n1321), .C2(new_n1315), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT60), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1336), .B1(new_n1202), .B2(new_n1209), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n978), .A2(new_n991), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1338), .A2(KEYINPUT60), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1337), .A2(new_n1339), .A3(new_n741), .A4(new_n1210), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n1310), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n894), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1340), .A2(G384), .A3(new_n1310), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1333), .A2(G2897), .ZN(new_n1345));
  XNOR2_X1  g1145(.A(new_n1344), .B(new_n1345), .ZN(new_n1346));
  AOI21_X1  g1146(.A(KEYINPUT61), .B1(new_n1335), .B2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(G375), .A2(G378), .ZN(new_n1348));
  AND2_X1   g1148(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1333), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1348), .A2(new_n1349), .A3(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(KEYINPUT62), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT62), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1348), .A2(new_n1353), .A3(new_n1350), .A4(new_n1349), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1347), .A2(new_n1352), .A3(new_n1354), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1172), .B1(new_n1176), .B2(new_n780), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n851), .B1(new_n1102), .B2(new_n1147), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1358), .B1(new_n1323), .B2(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(G393), .A2(G396), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1361), .A2(G390), .A3(new_n1322), .ZN(new_n1362));
  AND3_X1   g1162(.A1(new_n1360), .A2(new_n1362), .A3(new_n1095), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1095), .B1(new_n1360), .B2(new_n1362), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1355), .A2(new_n1366), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT63), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1351), .A2(new_n1368), .ZN(new_n1369));
  NAND4_X1  g1169(.A1(new_n1348), .A2(KEYINPUT63), .A3(new_n1350), .A4(new_n1349), .ZN(new_n1370));
  NAND4_X1  g1170(.A1(new_n1347), .A2(new_n1365), .A3(new_n1369), .A4(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1367), .A2(new_n1371), .ZN(G405));
  NOR2_X1   g1172(.A1(new_n1349), .A2(KEYINPUT126), .ZN(new_n1373));
  INV_X1    g1173(.A(KEYINPUT126), .ZN(new_n1374));
  NOR2_X1   g1174(.A1(new_n1344), .A2(new_n1374), .ZN(new_n1375));
  NOR2_X1   g1175(.A1(new_n1373), .A2(new_n1375), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1325), .A2(new_n1348), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1376), .A2(new_n1377), .ZN(new_n1378));
  OAI211_X1 g1178(.A(new_n1325), .B(new_n1348), .C1(new_n1373), .C2(new_n1375), .ZN(new_n1379));
  AND3_X1   g1179(.A1(new_n1365), .A2(new_n1378), .A3(new_n1379), .ZN(new_n1380));
  AOI21_X1  g1180(.A(new_n1365), .B1(new_n1379), .B2(new_n1378), .ZN(new_n1381));
  NOR2_X1   g1181(.A1(new_n1380), .A2(new_n1381), .ZN(G402));
endmodule


