

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593;

  NAND2_X1 U323 ( .A1(n577), .A2(n557), .ZN(n381) );
  INV_X1 U324 ( .A(n523), .ZN(n464) );
  XNOR2_X2 U325 ( .A(n452), .B(n451), .ZN(n455) );
  NOR2_X1 U326 ( .A1(n456), .A2(n545), .ZN(n459) );
  BUF_X1 U327 ( .A(n400), .Z(n348) );
  XNOR2_X1 U328 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U329 ( .A(G211GAT), .B(KEYINPUT21), .Z(n291) );
  XOR2_X1 U330 ( .A(n371), .B(n370), .Z(n292) );
  XOR2_X1 U331 ( .A(KEYINPUT36), .B(KEYINPUT92), .Z(n293) );
  XOR2_X1 U332 ( .A(n427), .B(n343), .Z(n294) );
  XNOR2_X1 U333 ( .A(n381), .B(KEYINPUT46), .ZN(n397) );
  XNOR2_X1 U334 ( .A(G162GAT), .B(KEYINPUT65), .ZN(n338) );
  NOR2_X1 U335 ( .A1(n577), .A2(n405), .ZN(n406) );
  INV_X1 U336 ( .A(KEYINPUT70), .ZN(n374) );
  INV_X1 U337 ( .A(n393), .ZN(n319) );
  XNOR2_X1 U338 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U339 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U340 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U341 ( .A(n347), .B(n346), .ZN(n400) );
  XNOR2_X1 U342 ( .A(n322), .B(n321), .ZN(n324) );
  XNOR2_X1 U343 ( .A(n400), .B(n293), .ZN(n591) );
  NOR2_X1 U344 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U345 ( .A(n328), .B(n437), .ZN(n523) );
  XNOR2_X1 U346 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n453) );
  XNOR2_X1 U347 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XOR2_X1 U348 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n296) );
  XNOR2_X1 U349 ( .A(KEYINPUT84), .B(KEYINPUT82), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n296), .B(n295), .ZN(n313) );
  XOR2_X1 U351 ( .A(KEYINPUT83), .B(KEYINPUT1), .Z(n298) );
  XNOR2_X1 U352 ( .A(KEYINPUT85), .B(KEYINPUT6), .ZN(n297) );
  XNOR2_X1 U353 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U354 ( .A(n299), .B(G85GAT), .Z(n301) );
  XOR2_X1 U355 ( .A(G120GAT), .B(G148GAT), .Z(n371) );
  XNOR2_X1 U356 ( .A(n371), .B(G57GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n306) );
  XOR2_X1 U358 ( .A(G29GAT), .B(G134GAT), .Z(n342) );
  XNOR2_X1 U359 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n302), .B(KEYINPUT75), .ZN(n436) );
  XOR2_X1 U361 ( .A(n342), .B(n436), .Z(n304) );
  NAND2_X1 U362 ( .A1(G225GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U363 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U364 ( .A(n306), .B(n305), .Z(n311) );
  XNOR2_X1 U365 ( .A(G1GAT), .B(G127GAT), .ZN(n307) );
  XNOR2_X1 U366 ( .A(n307), .B(G155GAT), .ZN(n385) );
  XOR2_X1 U367 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n309) );
  XNOR2_X1 U368 ( .A(G141GAT), .B(G162GAT), .ZN(n308) );
  XNOR2_X1 U369 ( .A(n309), .B(n308), .ZN(n426) );
  XNOR2_X1 U370 ( .A(n385), .B(n426), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U372 ( .A(n313), .B(n312), .Z(n475) );
  XNOR2_X1 U373 ( .A(KEYINPUT86), .B(n475), .ZN(n520) );
  XNOR2_X1 U374 ( .A(G197GAT), .B(KEYINPUT80), .ZN(n314) );
  XNOR2_X1 U375 ( .A(n291), .B(n314), .ZN(n427) );
  XOR2_X1 U376 ( .A(G36GAT), .B(G190GAT), .Z(n343) );
  NAND2_X1 U377 ( .A1(G226GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U378 ( .A(n294), .B(n315), .ZN(n316) );
  XOR2_X1 U379 ( .A(n316), .B(KEYINPUT88), .Z(n322) );
  XOR2_X1 U380 ( .A(G64GAT), .B(G204GAT), .Z(n318) );
  XNOR2_X1 U381 ( .A(G176GAT), .B(KEYINPUT71), .ZN(n317) );
  XNOR2_X1 U382 ( .A(n318), .B(n317), .ZN(n367) );
  XNOR2_X1 U383 ( .A(n367), .B(KEYINPUT87), .ZN(n320) );
  XOR2_X1 U384 ( .A(G8GAT), .B(G183GAT), .Z(n393) );
  XNOR2_X1 U385 ( .A(G218GAT), .B(G92GAT), .ZN(n323) );
  XNOR2_X1 U386 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U387 ( .A(KEYINPUT19), .B(KEYINPUT77), .Z(n326) );
  XNOR2_X1 U388 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n325) );
  XNOR2_X1 U389 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U390 ( .A(G169GAT), .B(n327), .Z(n437) );
  XNOR2_X1 U391 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n329) );
  XNOR2_X1 U392 ( .A(n329), .B(KEYINPUT7), .ZN(n351) );
  INV_X1 U393 ( .A(G106GAT), .ZN(n330) );
  NAND2_X1 U394 ( .A1(n330), .A2(G85GAT), .ZN(n333) );
  INV_X1 U395 ( .A(G85GAT), .ZN(n331) );
  NAND2_X1 U396 ( .A1(n331), .A2(G106GAT), .ZN(n332) );
  NAND2_X1 U397 ( .A1(n333), .A2(n332), .ZN(n335) );
  XNOR2_X1 U398 ( .A(G99GAT), .B(G92GAT), .ZN(n334) );
  XNOR2_X1 U399 ( .A(n335), .B(n334), .ZN(n373) );
  XNOR2_X1 U400 ( .A(n351), .B(n373), .ZN(n336) );
  XNOR2_X1 U401 ( .A(n336), .B(KEYINPUT11), .ZN(n341) );
  AND2_X1 U402 ( .A1(G232GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U404 ( .A(KEYINPUT9), .B(n339), .Z(n340) );
  XNOR2_X1 U405 ( .A(n341), .B(n340), .ZN(n347) );
  XOR2_X1 U406 ( .A(KEYINPUT10), .B(n342), .Z(n345) );
  XOR2_X1 U407 ( .A(G50GAT), .B(G218GAT), .Z(n417) );
  XNOR2_X1 U408 ( .A(n343), .B(n417), .ZN(n344) );
  XOR2_X1 U409 ( .A(G8GAT), .B(G197GAT), .Z(n350) );
  XNOR2_X1 U410 ( .A(G169GAT), .B(G29GAT), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n364) );
  XOR2_X1 U412 ( .A(G22GAT), .B(G15GAT), .Z(n394) );
  XOR2_X1 U413 ( .A(n394), .B(n351), .Z(n353) );
  XNOR2_X1 U414 ( .A(G50GAT), .B(G36GAT), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U416 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n355) );
  NAND2_X1 U417 ( .A1(G229GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U418 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U419 ( .A(n357), .B(n356), .Z(n362) );
  XOR2_X1 U420 ( .A(KEYINPUT29), .B(G113GAT), .Z(n359) );
  XNOR2_X1 U421 ( .A(G1GAT), .B(G141GAT), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n360), .B(KEYINPUT30), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n577) );
  XOR2_X1 U426 ( .A(G57GAT), .B(G78GAT), .Z(n366) );
  XNOR2_X1 U427 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n366), .B(n365), .ZN(n386) );
  XNOR2_X1 U429 ( .A(n367), .B(n386), .ZN(n379) );
  XOR2_X1 U430 ( .A(KEYINPUT33), .B(KEYINPUT69), .Z(n369) );
  XNOR2_X1 U431 ( .A(KEYINPUT32), .B(KEYINPUT72), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n370) );
  NAND2_X1 U433 ( .A1(G230GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n292), .B(n372), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n373), .B(KEYINPUT31), .ZN(n375) );
  XOR2_X1 U436 ( .A(n379), .B(n378), .Z(n582) );
  INV_X1 U437 ( .A(KEYINPUT41), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n582), .B(n380), .ZN(n557) );
  XOR2_X1 U439 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n383) );
  NAND2_X1 U440 ( .A1(G231GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U442 ( .A(n384), .B(KEYINPUT73), .Z(n388) );
  XNOR2_X1 U443 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U445 ( .A(KEYINPUT74), .B(KEYINPUT15), .Z(n390) );
  XNOR2_X1 U446 ( .A(G64GAT), .B(G211GAT), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U448 ( .A(n392), .B(n391), .Z(n396) );
  XNOR2_X1 U449 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U450 ( .A(n396), .B(n395), .ZN(n562) );
  XOR2_X1 U451 ( .A(n562), .B(KEYINPUT105), .Z(n545) );
  NAND2_X1 U452 ( .A1(n397), .A2(n545), .ZN(n398) );
  NOR2_X1 U453 ( .A1(n348), .A2(n398), .ZN(n399) );
  XOR2_X1 U454 ( .A(KEYINPUT47), .B(n399), .Z(n408) );
  INV_X1 U455 ( .A(KEYINPUT45), .ZN(n402) );
  NOR2_X1 U456 ( .A1(n562), .A2(n591), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n402), .B(n401), .ZN(n403) );
  NOR2_X1 U458 ( .A1(n582), .A2(n403), .ZN(n404) );
  XOR2_X1 U459 ( .A(KEYINPUT106), .B(n404), .Z(n405) );
  XOR2_X1 U460 ( .A(KEYINPUT107), .B(n406), .Z(n407) );
  NOR2_X1 U461 ( .A1(n408), .A2(n407), .ZN(n409) );
  XNOR2_X1 U462 ( .A(KEYINPUT48), .B(n409), .ZN(n532) );
  NOR2_X1 U463 ( .A1(n464), .A2(n532), .ZN(n411) );
  XNOR2_X1 U464 ( .A(KEYINPUT54), .B(KEYINPUT117), .ZN(n410) );
  XNOR2_X1 U465 ( .A(n411), .B(n410), .ZN(n412) );
  NOR2_X1 U466 ( .A1(n520), .A2(n412), .ZN(n413) );
  XNOR2_X1 U467 ( .A(n413), .B(KEYINPUT64), .ZN(n576) );
  XOR2_X1 U468 ( .A(G155GAT), .B(G106GAT), .Z(n415) );
  XNOR2_X1 U469 ( .A(G204GAT), .B(G78GAT), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U471 ( .A(n417), .B(n416), .Z(n419) );
  NAND2_X1 U472 ( .A1(G228GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U473 ( .A(n419), .B(n418), .ZN(n431) );
  XOR2_X1 U474 ( .A(KEYINPUT81), .B(KEYINPUT79), .Z(n421) );
  XNOR2_X1 U475 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n420) );
  XNOR2_X1 U476 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U477 ( .A(KEYINPUT78), .B(KEYINPUT23), .Z(n423) );
  XNOR2_X1 U478 ( .A(G22GAT), .B(G148GAT), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U480 ( .A(n425), .B(n424), .Z(n429) );
  XNOR2_X1 U481 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U483 ( .A(n431), .B(n430), .Z(n468) );
  NAND2_X1 U484 ( .A1(n576), .A2(n468), .ZN(n433) );
  XOR2_X1 U485 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n432) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n450) );
  XOR2_X1 U487 ( .A(G120GAT), .B(G71GAT), .Z(n435) );
  XNOR2_X1 U488 ( .A(G15GAT), .B(G127GAT), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n441) );
  XOR2_X1 U490 ( .A(KEYINPUT76), .B(KEYINPUT20), .Z(n439) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n449) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n447) );
  XOR2_X1 U495 ( .A(G183GAT), .B(G176GAT), .Z(n443) );
  XNOR2_X1 U496 ( .A(G43GAT), .B(G134GAT), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U498 ( .A(G190GAT), .B(G99GAT), .Z(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n449), .B(n448), .ZN(n463) );
  NOR2_X2 U502 ( .A1(n450), .A2(n463), .ZN(n452) );
  INV_X1 U503 ( .A(KEYINPUT119), .ZN(n451) );
  NAND2_X1 U504 ( .A1(n455), .A2(n348), .ZN(n454) );
  INV_X1 U505 ( .A(n455), .ZN(n456) );
  XNOR2_X1 U506 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n457) );
  XNOR2_X1 U507 ( .A(n457), .B(G183GAT), .ZN(n458) );
  XNOR2_X1 U508 ( .A(n459), .B(n458), .ZN(G1350GAT) );
  INV_X1 U509 ( .A(n577), .ZN(n536) );
  OR2_X1 U510 ( .A1(n582), .A2(n536), .ZN(n493) );
  NOR2_X1 U511 ( .A1(n348), .A2(n562), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n460), .B(KEYINPUT16), .ZN(n479) );
  INV_X1 U513 ( .A(n463), .ZN(n535) );
  INV_X1 U514 ( .A(n520), .ZN(n461) );
  XNOR2_X1 U515 ( .A(n464), .B(KEYINPUT27), .ZN(n471) );
  NOR2_X1 U516 ( .A1(n461), .A2(n471), .ZN(n552) );
  XNOR2_X1 U517 ( .A(n468), .B(KEYINPUT66), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT28), .ZN(n486) );
  NAND2_X1 U519 ( .A1(n552), .A2(n486), .ZN(n533) );
  NOR2_X1 U520 ( .A1(n535), .A2(n533), .ZN(n477) );
  NOR2_X1 U521 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U522 ( .A(KEYINPUT89), .B(n465), .ZN(n466) );
  NAND2_X1 U523 ( .A1(n466), .A2(n468), .ZN(n467) );
  XNOR2_X1 U524 ( .A(n467), .B(KEYINPUT25), .ZN(n473) );
  NOR2_X1 U525 ( .A1(n468), .A2(n535), .ZN(n469) );
  XNOR2_X1 U526 ( .A(n469), .B(KEYINPUT26), .ZN(n575) );
  INV_X1 U527 ( .A(n575), .ZN(n470) );
  NOR2_X1 U528 ( .A1(n471), .A2(n470), .ZN(n472) );
  NOR2_X1 U529 ( .A1(n473), .A2(n472), .ZN(n474) );
  NOR2_X1 U530 ( .A1(n475), .A2(n474), .ZN(n476) );
  NOR2_X1 U531 ( .A1(n477), .A2(n476), .ZN(n490) );
  INV_X1 U532 ( .A(n490), .ZN(n478) );
  NAND2_X1 U533 ( .A1(n479), .A2(n478), .ZN(n507) );
  NOR2_X1 U534 ( .A1(n493), .A2(n507), .ZN(n487) );
  NAND2_X1 U535 ( .A1(n520), .A2(n487), .ZN(n480) );
  XNOR2_X1 U536 ( .A(n480), .B(KEYINPUT34), .ZN(n481) );
  XNOR2_X1 U537 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  NAND2_X1 U538 ( .A1(n523), .A2(n487), .ZN(n482) );
  XNOR2_X1 U539 ( .A(n482), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT90), .B(KEYINPUT35), .Z(n484) );
  NAND2_X1 U541 ( .A1(n487), .A2(n535), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U543 ( .A(G15GAT), .B(n485), .ZN(G1326GAT) );
  XOR2_X1 U544 ( .A(G22GAT), .B(KEYINPUT91), .Z(n489) );
  INV_X1 U545 ( .A(n486), .ZN(n526) );
  NAND2_X1 U546 ( .A1(n487), .A2(n526), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(G1327GAT) );
  XOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT39), .Z(n497) );
  NOR2_X1 U549 ( .A1(n490), .A2(n591), .ZN(n491) );
  NAND2_X1 U550 ( .A1(n491), .A2(n562), .ZN(n492) );
  XOR2_X1 U551 ( .A(KEYINPUT37), .B(n492), .Z(n517) );
  NOR2_X1 U552 ( .A1(n517), .A2(n493), .ZN(n495) );
  XOR2_X1 U553 ( .A(KEYINPUT38), .B(KEYINPUT93), .Z(n494) );
  XNOR2_X1 U554 ( .A(n495), .B(n494), .ZN(n503) );
  NAND2_X1 U555 ( .A1(n503), .A2(n520), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(G1328GAT) );
  NAND2_X1 U557 ( .A1(n503), .A2(n523), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n498), .B(KEYINPUT94), .ZN(n499) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(n499), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT40), .B(KEYINPUT95), .Z(n501) );
  NAND2_X1 U561 ( .A1(n535), .A2(n503), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n502), .ZN(G1330GAT) );
  NAND2_X1 U564 ( .A1(n503), .A2(n526), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n504), .B(KEYINPUT96), .ZN(n505) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(n505), .ZN(G1331GAT) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n509) );
  XOR2_X1 U568 ( .A(KEYINPUT97), .B(n557), .Z(n572) );
  NAND2_X1 U569 ( .A1(n572), .A2(n536), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(KEYINPUT98), .ZN(n518) );
  NOR2_X1 U571 ( .A1(n518), .A2(n507), .ZN(n512) );
  NAND2_X1 U572 ( .A1(n512), .A2(n520), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n523), .A2(n512), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n510), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n512), .A2(n535), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT99), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U579 ( .A1(n512), .A2(n526), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(n516) );
  XOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT100), .Z(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(KEYINPUT102), .ZN(n522) );
  XOR2_X1 U584 ( .A(KEYINPUT101), .B(n519), .Z(n527) );
  NAND2_X1 U585 ( .A1(n527), .A2(n520), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n523), .A2(n527), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n524), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n527), .A2(n535), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n531) );
  NAND2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n529) );
  XOR2_X1 U593 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1339GAT) );
  NOR2_X1 U596 ( .A1(n532), .A2(n533), .ZN(n534) );
  NAND2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n544) );
  NOR2_X1 U598 ( .A1(n536), .A2(n544), .ZN(n537) );
  XOR2_X1 U599 ( .A(G113GAT), .B(n537), .Z(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT108), .Z(n539) );
  INV_X1 U601 ( .A(n544), .ZN(n549) );
  NAND2_X1 U602 ( .A1(n549), .A2(n572), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U604 ( .A(KEYINPUT49), .B(KEYINPUT109), .Z(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT112), .Z(n543) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(KEYINPUT111), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n547) );
  NOR2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U610 ( .A(n547), .B(n546), .Z(n548) );
  XNOR2_X1 U611 ( .A(KEYINPUT110), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U613 ( .A1(n549), .A2(n348), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n552), .A2(n575), .ZN(n553) );
  NOR2_X1 U616 ( .A1(n532), .A2(n553), .ZN(n565) );
  NAND2_X1 U617 ( .A1(n577), .A2(n565), .ZN(n554) );
  XNOR2_X1 U618 ( .A(n554), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT115), .B(KEYINPUT114), .Z(n556) );
  XNOR2_X1 U620 ( .A(KEYINPUT113), .B(KEYINPUT53), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(n561) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n559) );
  NAND2_X1 U623 ( .A1(n565), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  INV_X1 U626 ( .A(n562), .ZN(n587) );
  NAND2_X1 U627 ( .A1(n587), .A2(n565), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n563), .B(KEYINPUT116), .ZN(n564) );
  XNOR2_X1 U629 ( .A(G155GAT), .B(n564), .ZN(G1346GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n348), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U632 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n455), .A2(n577), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1348GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n570) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U638 ( .A(KEYINPUT56), .B(n571), .Z(n574) );
  NAND2_X1 U639 ( .A1(n455), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1349GAT) );
  XOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT125), .Z(n579) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n590) );
  INV_X1 U643 ( .A(n590), .ZN(n588) );
  NAND2_X1 U644 ( .A1(n588), .A2(n577), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n581) );
  XOR2_X1 U646 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n584) );
  NAND2_X1 U649 ( .A1(n588), .A2(n582), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n586) );
  XOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT126), .Z(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(G211GAT), .B(n589), .ZN(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(n592), .Z(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

