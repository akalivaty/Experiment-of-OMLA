//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n614, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT67), .Z(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT68), .ZN(G160));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n463), .B1(new_n477), .B2(new_n478), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI211_X1 g061(.A(G138), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n477), .A2(new_n478), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n489), .A2(new_n490), .A3(G138), .A4(new_n463), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n463), .A2(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT69), .A4(G2104), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n496), .A2(new_n500), .B1(new_n481), .B2(G126), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n492), .A2(new_n501), .A3(KEYINPUT70), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT70), .B1(new_n492), .B2(new_n501), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(G164));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  OR2_X1    g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT5), .B(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n505), .A2(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n513), .A2(new_n516), .ZN(G166));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n506), .A2(new_n507), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n521), .A2(G51), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  XOR2_X1   g101(.A(KEYINPUT5), .B(G543), .Z(new_n527));
  NAND2_X1  g102(.A1(new_n508), .A2(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n518), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n528), .A2(new_n529), .ZN(new_n532));
  OAI211_X1 g107(.A(KEYINPUT71), .B(new_n525), .C1(new_n532), .C2(new_n527), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(G168));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n535), .A2(new_n509), .B1(new_n511), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n515), .ZN(new_n539));
  OAI21_X1  g114(.A(KEYINPUT72), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n539), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n527), .A2(new_n519), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n542), .A2(G90), .B1(new_n521), .B2(G52), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n540), .A2(new_n545), .ZN(G171));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n547), .A2(new_n509), .B1(new_n511), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n515), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(new_n553));
  XOR2_X1   g128(.A(new_n553), .B(KEYINPUT73), .Z(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT75), .ZN(new_n557));
  XOR2_X1   g132(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n558));
  XNOR2_X1  g133(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(new_n521), .A2(G53), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n527), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G651), .B1(new_n542), .B2(G91), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n568));
  NAND2_X1  g143(.A1(G171), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n540), .A2(new_n545), .A3(KEYINPUT76), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n570), .A2(new_n572), .ZN(G301));
  INV_X1    g148(.A(G168), .ZN(G286));
  INV_X1    g149(.A(G166), .ZN(G303));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n576));
  INV_X1    g151(.A(G49), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n509), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n521), .A2(KEYINPUT77), .A3(G49), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n510), .A2(G74), .ZN(new_n581));
  AOI22_X1  g156(.A1(G651), .A2(new_n581), .B1(new_n542), .B2(G87), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(G288));
  AOI22_X1  g158(.A1(new_n542), .A2(G86), .B1(new_n521), .B2(G48), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n510), .A2(G61), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n515), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(KEYINPUT78), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n589));
  AOI211_X1 g164(.A(new_n589), .B(new_n515), .C1(new_n585), .C2(new_n586), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n584), .B1(new_n588), .B2(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OR3_X1    g167(.A1(new_n592), .A2(KEYINPUT79), .A3(new_n515), .ZN(new_n593));
  OAI21_X1  g168(.A(KEYINPUT79), .B1(new_n592), .B2(new_n515), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n542), .A2(G85), .B1(new_n521), .B2(G47), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(G290));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n511), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n542), .A2(KEYINPUT10), .A3(G92), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n527), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(new_n521), .B2(G54), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(G301), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G321));
  XOR2_X1   g184(.A(G321), .B(KEYINPUT80), .Z(G284));
  NOR2_X1   g185(.A1(G299), .A2(G868), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(G868), .B2(G168), .ZN(G280));
  XOR2_X1   g187(.A(G280), .B(KEYINPUT81), .Z(G297));
  INV_X1    g188(.A(new_n606), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g195(.A1(new_n476), .A2(G2105), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n489), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n479), .A2(G135), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n481), .A2(G123), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n463), .A2(G111), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n628), .B(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2096), .Z(new_n633));
  NAND3_X1  g208(.A1(new_n626), .A2(new_n627), .A3(new_n633), .ZN(G156));
  INV_X1    g209(.A(G14), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2430), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n640), .A2(new_n641), .ZN(new_n646));
  XOR2_X1   g221(.A(G2443), .B(G2446), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n648), .B1(new_n645), .B2(new_n646), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n638), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n653), .A2(new_n637), .A3(new_n649), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n635), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g234(.A(KEYINPUT83), .B1(new_n655), .B2(new_n657), .ZN(new_n660));
  AND3_X1   g235(.A1(new_n655), .A2(KEYINPUT83), .A3(new_n657), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G401));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  XNOR2_X1  g239(.A(G2072), .B(G2078), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT18), .Z(new_n668));
  AOI21_X1  g243(.A(new_n666), .B1(new_n665), .B2(KEYINPUT84), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(KEYINPUT84), .B2(new_n665), .ZN(new_n670));
  INV_X1    g245(.A(new_n664), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n665), .B(KEYINPUT17), .Z(new_n672));
  INV_X1    g247(.A(new_n666), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n670), .B(new_n671), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(new_n673), .A3(new_n664), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n668), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT87), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XOR2_X1   g256(.A(new_n680), .B(new_n681), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1956), .B(G2474), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT85), .ZN(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n685), .A2(new_n686), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n692), .A2(new_n689), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n692), .A2(new_n687), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(KEYINPUT86), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(KEYINPUT86), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n696), .A2(new_n689), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1991), .B(G1996), .Z(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n699), .A2(new_n700), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n683), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n703), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n705), .A2(new_n701), .A3(new_n682), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(G229));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G23), .ZN(new_n710));
  INV_X1    g285(.A(G288), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT33), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1976), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n709), .A2(G6), .ZN(new_n715));
  INV_X1    g290(.A(G305), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n709), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT32), .B(G1981), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n709), .A2(G22), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT88), .Z(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G303), .B2(G16), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G1971), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n714), .A2(new_n719), .A3(new_n720), .A4(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(KEYINPUT34), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(KEYINPUT34), .ZN(new_n727));
  MUX2_X1   g302(.A(G24), .B(G290), .S(G16), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G1986), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n728), .A2(G1986), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G25), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n479), .A2(G131), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n481), .A2(G119), .ZN(new_n734));
  OR2_X1    g309(.A1(G95), .A2(G2105), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n735), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n732), .B1(new_n738), .B2(new_n731), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT35), .B(G1991), .Z(new_n740));
  XOR2_X1   g315(.A(new_n739), .B(new_n740), .Z(new_n741));
  NOR3_X1   g316(.A1(new_n730), .A2(new_n741), .A3(KEYINPUT89), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n726), .A2(new_n727), .A3(new_n729), .A4(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT36), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n709), .A2(G4), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n614), .B2(new_n709), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1348), .ZN(new_n749));
  NOR2_X1   g324(.A1(G16), .A2(G19), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n552), .B2(G16), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G1341), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT30), .B(G28), .ZN(new_n753));
  OR2_X1    g328(.A1(KEYINPUT31), .A2(G11), .ZN(new_n754));
  NAND2_X1  g329(.A1(KEYINPUT31), .A2(G11), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n753), .A2(new_n731), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n752), .B(new_n756), .C1(new_n731), .C2(new_n632), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n751), .A2(G1341), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n731), .A2(G26), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT90), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT28), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n479), .A2(G140), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n481), .A2(G128), .ZN(new_n764));
  OR2_X1    g339(.A1(G104), .A2(G2105), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n765), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n762), .B1(new_n768), .B2(new_n731), .ZN(new_n769));
  INV_X1    g344(.A(G2067), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n731), .A2(G32), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n481), .A2(G129), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n621), .A2(G105), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G141), .B2(new_n479), .ZN(new_n776));
  NAND3_X1  g351(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT93), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT26), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n772), .B1(new_n781), .B2(new_n731), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT27), .B(G1996), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n759), .B(new_n771), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n731), .A2(G35), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G162), .B2(new_n731), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT29), .Z(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  AOI211_X1 g364(.A(new_n749), .B(new_n785), .C1(G2090), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n789), .A2(G2090), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n709), .A2(G21), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G168), .B2(new_n709), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT95), .B(G1966), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n709), .A2(G20), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT23), .Z(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G299), .B2(G16), .ZN(new_n798));
  INV_X1    g373(.A(G1956), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n791), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G34), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n802), .A2(KEYINPUT24), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(KEYINPUT24), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n731), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G160), .B2(new_n731), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT92), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n790), .B(new_n801), .C1(G2084), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n731), .A2(G33), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT91), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT25), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n489), .A2(G127), .ZN(new_n813));
  INV_X1    g388(.A(G115), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(new_n476), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n815), .A2(G2105), .B1(G139), .B2(new_n479), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n809), .B1(new_n818), .B2(new_n731), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(G2072), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n783), .A2(new_n784), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(G2072), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G2084), .B2(new_n807), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT94), .Z(new_n825));
  NOR2_X1   g400(.A1(G5), .A2(G16), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(G171), .B2(G16), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1961), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n731), .A2(G27), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(G164), .B2(new_n731), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G2078), .ZN(new_n831));
  NOR4_X1   g406(.A1(new_n808), .A2(new_n825), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n745), .A2(new_n746), .A3(new_n832), .ZN(G311));
  NAND3_X1  g408(.A1(new_n745), .A2(new_n746), .A3(new_n832), .ZN(G150));
  INV_X1    g409(.A(new_n552), .ZN(new_n835));
  INV_X1    g410(.A(G55), .ZN(new_n836));
  INV_X1    g411(.A(G93), .ZN(new_n837));
  OAI22_X1  g412(.A1(new_n836), .A2(new_n509), .B1(new_n511), .B2(new_n837), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n839), .A2(new_n515), .ZN(new_n840));
  OAI21_X1  g415(.A(KEYINPUT96), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n542), .A2(G93), .B1(new_n521), .B2(G55), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT96), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n842), .B(new_n843), .C1(new_n515), .C2(new_n839), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n835), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n838), .A2(new_n840), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n552), .A2(new_n846), .A3(new_n843), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n614), .A2(G559), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT39), .ZN(new_n852));
  AOI21_X1  g427(.A(G860), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n852), .B2(new_n851), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT97), .Z(new_n855));
  OAI21_X1  g430(.A(G860), .B1(new_n838), .B2(new_n840), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(G145));
  NOR2_X1   g433(.A1(new_n817), .A2(new_n780), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n479), .A2(G142), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n481), .A2(G130), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n463), .A2(G118), .ZN(new_n863));
  OAI21_X1  g438(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n861), .B(new_n862), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n623), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n817), .A2(new_n780), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n860), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n866), .B1(new_n870), .B2(new_n859), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n492), .A2(new_n501), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n767), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n737), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n869), .A3(new_n871), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(G160), .B(new_n632), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n485), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(G37), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT98), .ZN(new_n885));
  OR3_X1    g460(.A1(new_n879), .A2(new_n885), .A3(new_n881), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n885), .B1(new_n879), .B2(new_n881), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(KEYINPUT40), .Z(G395));
  NOR2_X1   g464(.A1(new_n846), .A2(G868), .ZN(new_n890));
  OR2_X1    g465(.A1(G166), .A2(KEYINPUT100), .ZN(new_n891));
  NAND2_X1  g466(.A1(G166), .A2(KEYINPUT100), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n716), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(G305), .A3(new_n892), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(G290), .B(G288), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n897), .A3(new_n895), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT42), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n848), .B(new_n617), .ZN(new_n903));
  NAND2_X1  g478(.A1(G299), .A2(new_n606), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n562), .A2(new_n601), .A3(new_n566), .A4(new_n605), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n905), .B1(new_n904), .B2(new_n906), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n903), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n904), .A2(new_n906), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n911), .B(KEYINPUT99), .Z(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n903), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n902), .B(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n890), .B1(new_n914), .B2(G868), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(G295));
  XNOR2_X1  g491(.A(new_n915), .B(KEYINPUT101), .ZN(G331));
  INV_X1    g492(.A(new_n911), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n845), .A2(new_n847), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n569), .A2(G168), .A3(new_n571), .ZN(new_n920));
  NAND2_X1  g495(.A1(G286), .A2(G171), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n919), .B1(new_n921), .B2(new_n920), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n918), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n920), .A2(new_n921), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n848), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n927), .B(new_n922), .C1(new_n907), .C2(new_n908), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n928), .A3(new_n901), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n925), .A2(new_n928), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n899), .A2(new_n900), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT102), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n901), .B1(new_n925), .B2(new_n928), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT102), .B1(new_n936), .B2(G37), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT43), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT103), .B1(new_n907), .B2(new_n908), .ZN(new_n939));
  OR2_X1    g514(.A1(new_n908), .A2(KEYINPUT103), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n927), .A2(new_n939), .A3(new_n940), .A4(new_n922), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n923), .A2(new_n924), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n932), .B(new_n941), .C1(new_n912), .C2(new_n942), .ZN(new_n943));
  AND4_X1   g518(.A1(KEYINPUT43), .A2(new_n943), .A3(new_n883), .A4(new_n929), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT44), .B1(new_n938), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  AND4_X1   g521(.A1(new_n946), .A2(new_n943), .A3(new_n883), .A4(new_n929), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n923), .A2(new_n924), .A3(new_n909), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n911), .B1(new_n927), .B2(new_n922), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n932), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(new_n934), .A3(new_n883), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n937), .A2(new_n951), .A3(new_n929), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n947), .B1(new_n952), .B2(KEYINPUT43), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n945), .B1(KEYINPUT44), .B2(new_n953), .ZN(G397));
  INV_X1    g529(.A(G1996), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n780), .B(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n767), .B(new_n770), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n738), .A2(new_n740), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n738), .A2(new_n740), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n956), .A2(new_n957), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(G1384), .B1(new_n492), .B2(new_n501), .ZN(new_n961));
  XNOR2_X1  g536(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G125), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n965), .B1(new_n477), .B2(new_n478), .ZN(new_n966));
  INV_X1    g541(.A(new_n467), .ZN(new_n967));
  OAI21_X1  g542(.A(G2105), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n470), .B1(new_n479), .B2(G137), .ZN(new_n969));
  XOR2_X1   g544(.A(KEYINPUT105), .B(G40), .Z(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT106), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n473), .A2(new_n974), .A3(new_n971), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n964), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(G290), .A2(G1986), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(G290), .A2(G1986), .ZN(new_n981));
  OR3_X1    g556(.A1(new_n980), .A2(KEYINPUT107), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n977), .B1(new_n980), .B2(KEYINPUT107), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n960), .A2(new_n978), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n975), .A2(new_n973), .B1(new_n961), .B2(KEYINPUT45), .ZN(new_n985));
  INV_X1    g560(.A(G2078), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT70), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n873), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n492), .A2(new_n501), .A3(KEYINPUT70), .ZN(new_n989));
  AOI21_X1  g564(.A(G1384), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n985), .B(new_n986), .C1(new_n990), .C2(new_n963), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT124), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT124), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n991), .A2(new_n995), .A3(new_n992), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n962), .A2(G1384), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n502), .B2(new_n503), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT116), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT116), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1001), .B(new_n998), .C1(new_n502), .C2(new_n503), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  INV_X1    g578(.A(G1384), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n873), .A2(new_n1004), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n1003), .A2(new_n1005), .B1(new_n973), .B2(new_n975), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1000), .A2(new_n986), .A3(new_n1002), .A4(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT123), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n974), .B1(new_n473), .B2(new_n971), .ZN(new_n1010));
  NOR4_X1   g585(.A1(new_n468), .A2(new_n472), .A3(KEYINPUT106), .A4(new_n970), .ZN(new_n1011));
  OAI22_X1  g586(.A1(new_n1010), .A2(new_n1011), .B1(new_n961), .B2(KEYINPUT45), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(KEYINPUT116), .B2(new_n999), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1013), .A2(KEYINPUT123), .A3(new_n986), .A4(new_n1002), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1009), .A2(new_n1014), .A3(KEYINPUT53), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1004), .B1(new_n502), .B2(new_n503), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT50), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n975), .A2(new_n973), .B1(new_n961), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1961), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n997), .A2(new_n1015), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n608), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT125), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1023), .A2(KEYINPUT125), .A3(new_n608), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT122), .ZN(new_n1029));
  AOI22_X1  g604(.A1(G286), .A2(G8), .B1(new_n1029), .B2(KEYINPUT51), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1031));
  INV_X1    g606(.A(G2084), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1000), .A2(new_n1002), .A3(new_n1006), .ZN(new_n1033));
  INV_X1    g608(.A(G1966), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1031), .A2(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G8), .ZN(new_n1036));
  OAI221_X1 g611(.A(new_n1030), .B1(new_n1029), .B2(KEYINPUT51), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1029), .A2(KEYINPUT51), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1036), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1030), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1038), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OR3_X1    g618(.A1(new_n1035), .A2(new_n1036), .A3(G168), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1037), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT62), .ZN(new_n1046));
  NAND3_X1  g621(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(G166), .B2(new_n1036), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1050), .B(KEYINPUT109), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1016), .A2(new_n962), .ZN(new_n1052));
  AOI21_X1  g627(.A(G1971), .B1(new_n1052), .B2(new_n985), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT108), .ZN(new_n1054));
  OAI22_X1  g629(.A1(new_n1053), .A2(new_n1054), .B1(new_n1020), .B2(G2090), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  OAI211_X1 g631(.A(G8), .B(new_n1051), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n584), .ZN(new_n1058));
  OAI21_X1  g633(.A(G1981), .B1(new_n1058), .B2(new_n587), .ZN(new_n1059));
  INV_X1    g634(.A(G1981), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n584), .B(new_n1060), .C1(new_n588), .C2(new_n590), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT49), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n976), .A2(new_n961), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1059), .A2(new_n1061), .A3(KEYINPUT49), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1064), .A2(G8), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(G8), .ZN(new_n1068));
  INV_X1    g643(.A(G1976), .ZN(new_n1069));
  NOR2_X1   g644(.A1(G288), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT52), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1070), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT110), .B(G1976), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(G288), .B2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1073), .A2(new_n1075), .A3(G8), .A4(new_n1065), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT111), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1072), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1057), .A2(new_n1080), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n1083));
  AOI22_X1  g658(.A1(KEYINPUT50), .A2(new_n1005), .B1(new_n973), .B2(new_n975), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1018), .B(new_n1004), .C1(new_n502), .C2(new_n503), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1084), .A2(KEYINPUT114), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT114), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1086), .A2(new_n1087), .A3(G2090), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1083), .B1(new_n1088), .B2(new_n1053), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1052), .A2(new_n985), .ZN(new_n1090));
  INV_X1    g665(.A(G1971), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1087), .A2(G2090), .ZN(new_n1093));
  OAI211_X1 g668(.A(KEYINPUT115), .B(new_n1092), .C1(new_n1093), .C2(new_n1086), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1089), .A2(new_n1094), .A3(G8), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1081), .B1(new_n1082), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT62), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1037), .A2(new_n1043), .A3(new_n1044), .A4(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1028), .A2(new_n1046), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1099));
  XOR2_X1   g674(.A(new_n1068), .B(KEYINPUT112), .Z(new_n1100));
  NAND2_X1  g675(.A1(new_n711), .A2(new_n1069), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1101), .B(KEYINPUT113), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1067), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1100), .B1(new_n1103), .B2(new_n1061), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1057), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(new_n1080), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n994), .A2(new_n996), .B1(new_n1021), .B2(new_n1020), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n1025), .B(G301), .C1(new_n1107), .C2(new_n1015), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT125), .B1(new_n1023), .B2(new_n608), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1022), .A2(KEYINPUT126), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT126), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n986), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n473), .B(new_n1114), .C1(new_n1005), .C2(new_n1003), .ZN(new_n1115));
  OAI22_X1  g690(.A1(new_n1111), .A2(new_n1113), .B1(new_n964), .B2(new_n1115), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n994), .A2(new_n996), .ZN(new_n1117));
  OR3_X1    g692(.A1(new_n1116), .A2(new_n1117), .A3(new_n608), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT54), .B1(new_n1110), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n799), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT56), .B(G2072), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1052), .A2(new_n985), .A3(new_n1122), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT57), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1125), .A2(KEYINPUT119), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(KEYINPUT119), .ZN(new_n1127));
  AND3_X1   g702(.A1(G299), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1127), .B1(G299), .B2(new_n1126), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1132));
  AOI21_X1  g707(.A(G1348), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1005), .B1(new_n975), .B2(new_n973), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n770), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(new_n606), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1131), .B1(new_n1132), .B2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(KEYINPUT60), .B(new_n1135), .C1(new_n1031), .C2(G1348), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT60), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(new_n1142), .A3(new_n614), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1124), .A2(new_n1144), .A3(new_n1145), .A4(new_n1130), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1130), .A2(new_n1144), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT61), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1143), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(KEYINPUT58), .B(G1341), .ZN(new_n1150));
  OAI22_X1  g725(.A1(new_n1090), .A2(G1996), .B1(new_n1134), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n835), .A2(KEYINPUT120), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT59), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1137), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1151), .A2(KEYINPUT59), .A3(new_n1152), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1139), .B1(new_n1149), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(G171), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1107), .A2(G301), .A3(new_n1015), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1160), .A2(KEYINPUT54), .A3(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1096), .A2(new_n1159), .A3(new_n1162), .A4(new_n1045), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1099), .B(new_n1106), .C1(new_n1119), .C2(new_n1163), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1035), .A2(new_n1036), .A3(G286), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT63), .B1(new_n1096), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(G8), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT117), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1082), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1092), .A2(KEYINPUT108), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1170), .B(new_n1171), .C1(G2090), .C2(new_n1020), .ZN(new_n1172));
  AOI21_X1  g747(.A(KEYINPUT117), .B1(new_n1172), .B2(G8), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1080), .B1(new_n1169), .B2(new_n1173), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1174), .A2(KEYINPUT118), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1057), .A2(new_n1165), .A3(KEYINPUT63), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1176), .B1(new_n1174), .B2(KEYINPUT118), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1166), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n984), .B1(new_n1164), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n981), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT48), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1180), .A2(new_n977), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(KEYINPUT48), .B1(new_n978), .B2(new_n981), .ZN(new_n1183));
  AOI211_X1 g758(.A(new_n1182), .B(new_n1183), .C1(new_n960), .C2(new_n978), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n977), .A2(G1996), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT46), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n977), .B1(new_n781), .B2(new_n957), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1188), .B(KEYINPUT47), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n956), .A2(new_n957), .ZN(new_n1190));
  OAI22_X1  g765(.A1(new_n1190), .A2(new_n959), .B1(G2067), .B2(new_n767), .ZN(new_n1191));
  AOI211_X1 g766(.A(new_n1184), .B(new_n1189), .C1(new_n978), .C2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1179), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g768(.A1(G227), .A2(new_n461), .ZN(new_n1195));
  AND3_X1   g769(.A1(new_n704), .A2(new_n706), .A3(new_n1195), .ZN(new_n1196));
  AND2_X1   g770(.A1(new_n886), .A2(new_n887), .ZN(new_n1197));
  OAI211_X1 g771(.A(new_n662), .B(new_n1196), .C1(new_n1197), .C2(new_n884), .ZN(new_n1198));
  OAI21_X1  g772(.A(KEYINPUT127), .B1(new_n953), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g773(.A1(new_n662), .A2(new_n1196), .ZN(new_n1200));
  NOR2_X1   g774(.A1(new_n1200), .A2(new_n888), .ZN(new_n1201));
  INV_X1    g775(.A(KEYINPUT127), .ZN(new_n1202));
  AOI21_X1  g776(.A(new_n946), .B1(new_n935), .B2(new_n937), .ZN(new_n1203));
  OAI211_X1 g777(.A(new_n1201), .B(new_n1202), .C1(new_n1203), .C2(new_n947), .ZN(new_n1204));
  AND2_X1   g778(.A1(new_n1199), .A2(new_n1204), .ZN(G308));
  NAND2_X1  g779(.A1(new_n1199), .A2(new_n1204), .ZN(G225));
endmodule


