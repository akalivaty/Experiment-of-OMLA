//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  INV_X1    g002(.A(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G141gat), .B(G148gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT75), .B(KEYINPUT2), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n203), .B(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n207), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n203), .B1(new_n206), .B2(KEYINPUT2), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT29), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT82), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  XOR2_X1   g018(.A(G197gat), .B(G204gat), .Z(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G211gat), .A2(G218gat), .ZN(new_n222));
  OR2_X1    g021(.A1(G211gat), .A2(G218gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT22), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n222), .B(new_n223), .C1(new_n220), .C2(new_n224), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n219), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n229), .A2(KEYINPUT29), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n213), .B1(new_n231), .B2(KEYINPUT3), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n202), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n229), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n227), .B(KEYINPUT81), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n226), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n214), .B1(new_n236), .B2(new_n216), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT77), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n213), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n209), .A2(new_n212), .A3(KEYINPUT77), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n202), .B(new_n234), .C1(new_n237), .C2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n233), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(KEYINPUT83), .A2(G22gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(G78gat), .B(G106gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT31), .B(G50gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  MUX2_X1   g048(.A(G22gat), .B(new_n246), .S(new_n249), .Z(new_n250));
  XNOR2_X1  g049(.A(new_n245), .B(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G8gat), .B(G36gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(G64gat), .B(G92gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G183gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT65), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G183gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n259), .A3(KEYINPUT27), .ZN(new_n260));
  NOR2_X1   g059(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(G190gat), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT67), .B1(new_n263), .B2(KEYINPUT28), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT28), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT65), .B(G183gat), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n261), .B1(new_n267), .B2(KEYINPUT27), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n265), .B(new_n266), .C1(new_n268), .C2(G190gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT27), .B(G183gat), .ZN(new_n270));
  INV_X1    g069(.A(G190gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(KEYINPUT28), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n264), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G169gat), .ZN(new_n274));
  INV_X1    g073(.A(G176gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n276), .A2(KEYINPUT26), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n277), .B1(G169gat), .B2(G176gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(KEYINPUT26), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n278), .A2(new_n279), .B1(G183gat), .B2(G190gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n274), .A2(new_n275), .A3(KEYINPUT23), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT23), .B1(new_n274), .B2(new_n275), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n282), .B1(new_n276), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT25), .ZN(new_n285));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT24), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n256), .A2(new_n271), .A3(KEYINPUT64), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT64), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n290), .B1(G183gat), .B2(G190gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n288), .A2(new_n289), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n284), .A2(new_n285), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n267), .A2(G190gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n288), .A2(new_n292), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT66), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n288), .A2(new_n292), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT66), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n298), .B(new_n299), .C1(G190gat), .C2(new_n267), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n297), .A2(new_n300), .A3(new_n284), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n294), .B1(new_n301), .B2(KEYINPUT25), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT29), .B1(new_n281), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G226gat), .ZN(new_n304));
  INV_X1    g103(.A(G233gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  AOI211_X1 g106(.A(new_n304), .B(new_n305), .C1(new_n281), .C2(new_n302), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n229), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n281), .A2(new_n302), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n306), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n311), .B(new_n228), .C1(new_n306), .C2(new_n303), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT87), .B(KEYINPUT37), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n309), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT88), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT88), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n309), .A2(new_n312), .A3(new_n316), .A4(new_n313), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n309), .A2(new_n312), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n315), .A2(new_n317), .B1(KEYINPUT37), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT38), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n255), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n315), .A2(new_n317), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT86), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n312), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n324), .B(KEYINPUT37), .C1(new_n318), .C2(KEYINPUT86), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n322), .A2(new_n320), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n318), .ZN(new_n328));
  INV_X1    g127(.A(new_n255), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n320), .ZN(new_n330));
  OAI22_X1  g129(.A1(new_n321), .A2(new_n327), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G120gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G113gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT69), .B(G113gat), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n333), .B1(new_n334), .B2(new_n332), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT1), .ZN(new_n336));
  XNOR2_X1  g135(.A(G127gat), .B(G134gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT70), .ZN(new_n339));
  INV_X1    g138(.A(new_n337), .ZN(new_n340));
  INV_X1    g139(.A(G113gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G120gat), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n333), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n340), .B(KEYINPUT68), .C1(new_n343), .C2(KEYINPUT1), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT68), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT1), .B1(new_n333), .B2(new_n342), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n345), .B1(new_n346), .B2(new_n337), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT70), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n335), .A2(new_n349), .A3(new_n336), .A4(new_n337), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n339), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n213), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(KEYINPUT4), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT4), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n348), .A3(new_n350), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n354), .B1(new_n355), .B2(new_n241), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n213), .A2(KEYINPUT3), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n215), .A3(new_n357), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n353), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n359), .A2(KEYINPUT79), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n353), .A2(new_n356), .A3(new_n358), .A4(new_n362), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n364), .B1(new_n365), .B2(new_n360), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G1gat), .B(G29gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(G85gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT0), .B(G57gat), .ZN(new_n370));
  XOR2_X1   g169(.A(new_n369), .B(new_n370), .Z(new_n371));
  XNOR2_X1  g170(.A(new_n355), .B(new_n213), .ZN(new_n372));
  INV_X1    g171(.A(new_n362), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n361), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n242), .A2(new_n351), .A3(KEYINPUT4), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n354), .B1(new_n355), .B2(new_n213), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n375), .A2(new_n362), .A3(new_n358), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n367), .A2(new_n371), .A3(new_n378), .ZN(new_n379));
  XOR2_X1   g178(.A(KEYINPUT80), .B(KEYINPUT6), .Z(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n363), .A2(new_n366), .B1(new_n374), .B2(new_n377), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n383), .A2(new_n371), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n383), .A2(new_n371), .A3(new_n381), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n252), .B1(new_n331), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT39), .B1(new_n372), .B2(new_n373), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT84), .ZN(new_n390));
  OR2_X1    g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OR2_X1    g190(.A1(new_n359), .A2(new_n362), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n390), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n394), .B(new_n371), .C1(KEYINPUT39), .C2(new_n392), .ZN(new_n395));
  NOR2_X1   g194(.A1(KEYINPUT85), .A2(KEYINPUT40), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT30), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n255), .B1(new_n318), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(new_n398), .B2(new_n318), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n328), .A2(KEYINPUT30), .A3(new_n255), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n367), .A2(new_n378), .ZN(new_n404));
  INV_X1    g203(.A(new_n371), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n395), .A2(new_n396), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n397), .A2(new_n403), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n402), .B1(new_n385), .B2(new_n386), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n388), .A2(new_n408), .B1(new_n409), .B2(new_n252), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT72), .ZN(new_n411));
  XNOR2_X1  g210(.A(G15gat), .B(G43gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(G71gat), .B(G99gat), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n412), .B(new_n413), .Z(new_n414));
  NAND2_X1  g213(.A1(G227gat), .A2(G233gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n310), .A2(new_n355), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n281), .A2(new_n351), .A3(new_n302), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT71), .B(KEYINPUT33), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n414), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT32), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n411), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n419), .ZN(new_n424));
  INV_X1    g223(.A(new_n414), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n415), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n281), .A2(new_n351), .A3(new_n302), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n351), .B1(new_n281), .B2(new_n302), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n425), .B1(new_n430), .B2(new_n424), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(KEYINPUT32), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(KEYINPUT72), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n423), .A2(new_n426), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n415), .A3(new_n417), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n435), .B(KEYINPUT34), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT73), .ZN(new_n438));
  INV_X1    g237(.A(new_n436), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n439), .A2(new_n423), .A3(new_n426), .A4(new_n433), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT36), .ZN(new_n442));
  INV_X1    g241(.A(new_n434), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(KEYINPUT73), .A3(new_n439), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT74), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n437), .A2(KEYINPUT36), .A3(new_n440), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n441), .A2(new_n444), .A3(KEYINPUT74), .A4(new_n442), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n251), .A2(new_n437), .A3(new_n440), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT35), .B1(new_n409), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT89), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g253(.A(KEYINPUT89), .B(KEYINPUT35), .C1(new_n409), .C2(new_n451), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n444), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT35), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n406), .A2(new_n379), .A3(new_n381), .ZN(new_n459));
  INV_X1    g258(.A(new_n386), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n459), .A2(new_n460), .B1(new_n401), .B2(new_n400), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n457), .A2(new_n458), .A3(new_n461), .A4(new_n251), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n410), .A2(new_n450), .B1(new_n456), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G99gat), .B(G106gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(KEYINPUT97), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(G99gat), .A2(G106gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT8), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT95), .B(G85gat), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(G92gat), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT96), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT96), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(G85gat), .A2(G92gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(KEYINPUT7), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n466), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n477), .ZN(new_n479));
  AOI211_X1 g278(.A(new_n479), .B(new_n465), .C1(new_n472), .C2(new_n474), .ZN(new_n480));
  XNOR2_X1  g279(.A(G71gat), .B(G78gat), .ZN(new_n481));
  XOR2_X1   g280(.A(G57gat), .B(G64gat), .Z(new_n482));
  INV_X1    g281(.A(KEYINPUT9), .ZN(new_n483));
  INV_X1    g282(.A(G71gat), .ZN(new_n484));
  INV_X1    g283(.A(G78gat), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n481), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n486), .A3(new_n481), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  OAI22_X1  g288(.A1(new_n478), .A2(new_n480), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n474), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n470), .A2(new_n473), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n477), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n465), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n489), .A2(new_n487), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n475), .A2(new_n477), .A3(new_n466), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT10), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n490), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n478), .A2(new_n480), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT94), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n489), .B2(new_n487), .ZN(new_n502));
  INV_X1    g301(.A(new_n487), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n503), .A2(KEYINPUT94), .A3(new_n488), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n500), .A2(KEYINPUT102), .A3(KEYINPUT10), .A4(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n494), .A2(new_n496), .A3(KEYINPUT10), .A4(new_n505), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT102), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n499), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G230gat), .A2(G233gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n490), .A2(new_n497), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(G230gat), .A3(G233gat), .ZN(new_n514));
  XOR2_X1   g313(.A(G176gat), .B(G204gat), .Z(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(G148gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT103), .B(G120gat), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n516), .B(new_n517), .Z(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n512), .A2(new_n514), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n511), .B(KEYINPUT104), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n510), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n519), .B1(new_n522), .B2(new_n514), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT92), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G1gat), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n529), .A2(KEYINPUT16), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(G8gat), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n528), .A2(new_n529), .ZN(new_n534));
  INV_X1    g333(.A(G8gat), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n534), .B(new_n535), .C1(new_n528), .C2(new_n531), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT17), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT14), .ZN(new_n539));
  INV_X1    g338(.A(G29gat), .ZN(new_n540));
  INV_X1    g339(.A(G36gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n542), .A2(new_n543), .B1(G29gat), .B2(G36gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT15), .ZN(new_n545));
  XOR2_X1   g344(.A(G43gat), .B(G50gat), .Z(new_n546));
  OR3_X1    g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n545), .ZN(new_n548));
  XNOR2_X1  g347(.A(G43gat), .B(G50gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT15), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n550), .A3(new_n544), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n547), .A2(KEYINPUT91), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT91), .B1(new_n547), .B2(new_n551), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n538), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n547), .A2(new_n551), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT17), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n537), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n552), .A2(new_n553), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n537), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NOR3_X1   g360(.A1(new_n557), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT93), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT18), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n537), .B(new_n558), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n560), .B(KEYINPUT13), .Z(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n554), .A2(new_n556), .ZN(new_n568));
  INV_X1    g367(.A(new_n537), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n537), .A2(new_n558), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(new_n571), .A3(new_n560), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT18), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(KEYINPUT93), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n564), .A2(new_n567), .A3(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(G169gat), .B(G197gat), .Z(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G113gat), .B(G141gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n580), .B(KEYINPUT12), .Z(new_n581));
  NAND2_X1  g380(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n581), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n564), .A2(new_n583), .A3(new_n574), .A4(new_n567), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NOR3_X1   g385(.A1(new_n463), .A2(new_n525), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G127gat), .B(G155gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(G211gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n495), .A2(KEYINPUT21), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n505), .A2(KEYINPUT21), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n569), .A2(new_n256), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n256), .B1(new_n569), .B2(new_n592), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n591), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n595), .ZN(new_n597));
  INV_X1    g396(.A(new_n591), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n593), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n596), .A2(new_n599), .A3(G231gat), .A4(G233gat), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n590), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n602), .A2(new_n603), .A3(new_n590), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n606), .B1(new_n605), .B2(new_n607), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT101), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n500), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT98), .B1(new_n478), .B2(new_n480), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(new_n568), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n558), .A2(new_n496), .A3(new_n494), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT99), .ZN(new_n617));
  AND2_X1   g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT41), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n617), .B1(new_n616), .B2(new_n619), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n615), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT100), .ZN(new_n623));
  XOR2_X1   g422(.A(G190gat), .B(G218gat), .Z(new_n624));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n625), .B(new_n615), .C1(new_n620), .C2(new_n621), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n624), .B1(new_n623), .B2(new_n626), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n611), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n624), .ZN(new_n630));
  INV_X1    g429(.A(new_n621), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n625), .B1(new_n633), .B2(new_n615), .ZN(new_n634));
  INV_X1    g433(.A(new_n626), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n630), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(KEYINPUT101), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n618), .A2(KEYINPUT41), .ZN(new_n639));
  XNOR2_X1  g438(.A(G134gat), .B(G162gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n629), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n611), .B(new_n641), .C1(new_n627), .C2(new_n628), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n610), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n587), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n387), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g448(.A1(new_n587), .A2(new_n646), .A3(new_n403), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT42), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT16), .B(G8gat), .ZN(new_n652));
  OR3_X1    g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n650), .B(KEYINPUT105), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n651), .B1(new_n654), .B2(G8gat), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(new_n652), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(G1325gat));
  AOI21_X1  g456(.A(G15gat), .B1(new_n647), .B2(new_n457), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n450), .A2(KEYINPUT106), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n447), .A2(new_n660), .A3(new_n448), .A4(new_n449), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n663), .A2(G15gat), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n658), .B1(new_n647), .B2(new_n664), .ZN(G1326gat));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n252), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n666), .A2(G22gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(G22gat), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n668), .B1(new_n667), .B2(new_n669), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(G1327gat));
  NOR2_X1   g471(.A1(new_n586), .A2(new_n525), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n610), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n328), .A2(new_n330), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n318), .A2(KEYINPUT37), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n322), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n329), .B1(new_n678), .B2(KEYINPUT38), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n676), .B1(new_n679), .B2(new_n326), .ZN(new_n680));
  INV_X1    g479(.A(new_n387), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n251), .B(new_n408), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n683), .B1(new_n461), .B2(new_n251), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n409), .A2(KEYINPUT108), .A3(new_n252), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n687), .B1(new_n659), .B2(new_n661), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n456), .A2(new_n462), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n675), .B(new_n645), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n643), .A2(new_n644), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT44), .B1(new_n463), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n674), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n693), .A2(new_n694), .A3(new_n387), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(new_n693), .B2(new_n387), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n695), .A2(new_n696), .A3(new_n540), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n463), .A2(new_n691), .A3(new_n674), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n698), .A2(new_n540), .A3(new_n387), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT45), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT110), .B1(new_n697), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n696), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n693), .A2(new_n694), .A3(new_n387), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(G29gat), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(new_n700), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n702), .A2(new_n707), .ZN(G1328gat));
  NAND3_X1  g507(.A1(new_n698), .A2(new_n541), .A3(new_n403), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT46), .Z(new_n710));
  NAND2_X1  g509(.A1(new_n690), .A2(new_n692), .ZN(new_n711));
  INV_X1    g510(.A(new_n674), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G36gat), .B1(new_n713), .B2(new_n402), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n710), .A2(new_n714), .ZN(G1329gat));
  AOI21_X1  g514(.A(G43gat), .B1(new_n698), .B2(new_n457), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n663), .A2(G43gat), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n716), .B1(new_n693), .B2(new_n717), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g518(.A(G50gat), .B1(new_n713), .B2(new_n251), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT111), .ZN(new_n721));
  INV_X1    g520(.A(G50gat), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n698), .A2(new_n722), .A3(new_n252), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n721), .A2(new_n724), .A3(KEYINPUT48), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n720), .B(new_n723), .C1(KEYINPUT111), .C2(new_n726), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n725), .A2(new_n727), .ZN(G1331gat));
  NOR2_X1   g527(.A1(new_n688), .A2(new_n689), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n524), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n610), .A2(new_n645), .A3(new_n585), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n681), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g533(.A1(new_n732), .A2(new_n402), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  AND2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n735), .B2(new_n736), .ZN(G1333gat));
  INV_X1    g538(.A(new_n457), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n484), .B1(new_n732), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n663), .A2(G71gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n732), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g543(.A1(new_n732), .A2(new_n251), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT112), .B(G78gat), .Z(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1335gat));
  NOR2_X1   g546(.A1(new_n608), .A2(new_n609), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n585), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n711), .A2(new_n525), .A3(new_n749), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT95), .B(G85gat), .Z(new_n751));
  NOR3_X1   g550(.A1(new_n750), .A2(new_n681), .A3(new_n751), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n645), .B(new_n749), .C1(new_n688), .C2(new_n689), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT51), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n524), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n387), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n752), .B1(new_n756), .B2(new_n751), .ZN(G1336gat));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n758), .A2(KEYINPUT52), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n758), .A2(KEYINPUT52), .ZN(new_n760));
  OAI21_X1  g559(.A(G92gat), .B1(new_n750), .B2(new_n402), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n753), .B(new_n762), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n402), .A2(G92gat), .A3(new_n524), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT113), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  AOI211_X1 g565(.A(new_n759), .B(new_n760), .C1(new_n761), .C2(new_n766), .ZN(new_n767));
  AND4_X1   g566(.A1(new_n758), .A2(new_n761), .A3(KEYINPUT52), .A4(new_n766), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(G1337gat));
  OR3_X1    g568(.A1(new_n750), .A2(KEYINPUT115), .A3(new_n662), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT115), .B1(new_n750), .B2(new_n662), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(G99gat), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(G99gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n773), .A3(new_n457), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(G1338gat));
  INV_X1    g574(.A(G106gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n755), .A2(new_n776), .A3(new_n252), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778));
  OAI21_X1  g577(.A(G106gat), .B1(new_n750), .B2(new_n251), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NOR4_X1   g579(.A1(new_n754), .A2(G106gat), .A3(new_n524), .A4(new_n251), .ZN(new_n781));
  INV_X1    g580(.A(new_n779), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT53), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(G1339gat));
  INV_X1    g583(.A(new_n521), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n499), .A2(new_n506), .A3(new_n509), .A4(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n512), .A2(KEYINPUT54), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n510), .A2(new_n788), .A3(new_n521), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n787), .A2(KEYINPUT55), .A3(new_n518), .A4(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n520), .B1(new_n790), .B2(KEYINPUT116), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n789), .A2(new_n518), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n787), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n792), .A2(new_n796), .A3(KEYINPUT55), .A4(new_n787), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n791), .A2(new_n585), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n565), .A2(new_n566), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n560), .B1(new_n570), .B2(new_n571), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n580), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n584), .B(new_n802), .C1(new_n523), .C2(new_n520), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n798), .A2(new_n799), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n799), .B1(new_n798), .B2(new_n803), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n804), .A2(new_n805), .A3(new_n645), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n795), .A3(new_n797), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n584), .A2(new_n802), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n645), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n610), .B1(new_n806), .B2(new_n811), .ZN(new_n812));
  AND4_X1   g611(.A1(new_n748), .A2(new_n691), .A3(new_n524), .A4(new_n586), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n681), .A2(new_n403), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n740), .A2(new_n252), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(G113gat), .B1(new_n819), .B2(new_n586), .ZN(new_n820));
  INV_X1    g619(.A(new_n451), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n586), .A2(new_n334), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n820), .B1(new_n822), .B2(new_n823), .ZN(G1340gat));
  OAI21_X1  g623(.A(G120gat), .B1(new_n819), .B2(new_n524), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n525), .A2(new_n332), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n822), .B2(new_n826), .ZN(G1341gat));
  INV_X1    g626(.A(G127gat), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n819), .A2(new_n828), .A3(new_n610), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n817), .A2(new_n748), .A3(new_n821), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n828), .B2(new_n830), .ZN(G1342gat));
  OR3_X1    g630(.A1(new_n822), .A2(G134gat), .A3(new_n691), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n832), .A2(KEYINPUT56), .ZN(new_n833));
  OAI21_X1  g632(.A(G134gat), .B1(new_n819), .B2(new_n691), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(KEYINPUT56), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(G1343gat));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(KEYINPUT121), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n837), .A2(KEYINPUT121), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n251), .B1(new_n812), .B2(new_n814), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT119), .B1(new_n840), .B2(KEYINPUT57), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n803), .A2(KEYINPUT120), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n803), .A2(KEYINPUT120), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n798), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n691), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n748), .B1(new_n845), .B2(new_n810), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n252), .B1(new_n846), .B2(new_n813), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n798), .A2(new_n803), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT117), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n798), .A2(new_n799), .A3(new_n803), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n691), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n748), .B1(new_n854), .B2(new_n810), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n813), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n850), .B(new_n848), .C1(new_n856), .C2(new_n251), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n849), .A3(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n662), .A2(new_n816), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT118), .ZN(new_n860));
  INV_X1    g659(.A(G141gat), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n586), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n858), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n840), .A2(new_n859), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n861), .B1(new_n864), .B2(new_n586), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n838), .B(new_n839), .C1(new_n863), .C2(new_n865), .ZN(new_n866));
  AND4_X1   g665(.A1(KEYINPUT121), .A2(new_n863), .A3(new_n837), .A4(new_n865), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(G1344gat));
  AND2_X1   g667(.A1(new_n860), .A2(new_n525), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n847), .A2(new_n848), .ZN(new_n870));
  OAI211_X1 g669(.A(KEYINPUT57), .B(new_n252), .C1(new_n855), .C2(new_n813), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n869), .A2(new_n875), .A3(new_n858), .ZN(new_n876));
  INV_X1    g675(.A(new_n864), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n875), .B1(new_n877), .B2(new_n525), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n874), .B(new_n876), .C1(G148gat), .C2(new_n878), .ZN(G1345gat));
  AOI21_X1  g678(.A(G155gat), .B1(new_n877), .B2(new_n748), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n858), .A2(new_n860), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n610), .A2(new_n204), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(G1346gat));
  AOI21_X1  g682(.A(G162gat), .B1(new_n877), .B2(new_n645), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n691), .A2(new_n205), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n881), .B2(new_n885), .ZN(G1347gat));
  NAND4_X1  g685(.A1(new_n815), .A2(new_n681), .A3(new_n403), .A4(new_n818), .ZN(new_n887));
  OAI21_X1  g686(.A(G169gat), .B1(new_n887), .B2(new_n586), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n815), .A2(new_n681), .A3(new_n403), .A4(new_n821), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n585), .A2(new_n274), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(G1348gat));
  NOR3_X1   g690(.A1(new_n887), .A2(new_n275), .A3(new_n524), .ZN(new_n892));
  INV_X1    g691(.A(new_n889), .ZN(new_n893));
  AOI21_X1  g692(.A(G176gat), .B1(new_n893), .B2(new_n525), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n894), .A2(KEYINPUT122), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(KEYINPUT122), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n892), .B1(new_n895), .B2(new_n896), .ZN(G1349gat));
  OAI21_X1  g696(.A(new_n267), .B1(new_n887), .B2(new_n610), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n899));
  AND4_X1   g698(.A1(new_n899), .A2(new_n893), .A3(new_n748), .A4(new_n270), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n889), .A2(new_n610), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n901), .B2(new_n270), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n898), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT60), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n905), .B(new_n898), .C1(new_n900), .C2(new_n902), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n887), .B2(new_n691), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(KEYINPUT61), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n893), .A2(new_n271), .A3(new_n645), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n908), .A2(new_n909), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(G1351gat));
  NOR3_X1   g715(.A1(new_n663), .A2(new_n387), .A3(new_n402), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n872), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(G197gat), .B1(new_n918), .B2(new_n586), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n840), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n586), .A2(G197gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(G1352gat));
  XNOR2_X1  g721(.A(KEYINPUT125), .B(G204gat), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n917), .A2(new_n525), .A3(new_n840), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT62), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n923), .B1(new_n918), .B2(new_n524), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n925), .A2(KEYINPUT62), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n928), .A2(KEYINPUT126), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n928), .A2(KEYINPUT126), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n926), .B(new_n927), .C1(new_n929), .C2(new_n930), .ZN(G1353gat));
  OR3_X1    g730(.A1(new_n920), .A2(G211gat), .A3(new_n610), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n872), .A2(new_n748), .A3(new_n917), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n872), .A2(KEYINPUT127), .A3(new_n748), .A4(new_n917), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n935), .A2(G211gat), .A3(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT63), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n932), .B1(new_n939), .B2(new_n940), .ZN(G1354gat));
  OAI21_X1  g740(.A(G218gat), .B1(new_n918), .B2(new_n691), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n691), .A2(G218gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n920), .B2(new_n943), .ZN(G1355gat));
endmodule


