//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G237), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G214), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(G237), .A2(G953), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(G143), .A3(G214), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(KEYINPUT81), .A2(KEYINPUT18), .A3(G131), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n198), .B(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G125), .B(G140), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  OR2_X1    g018(.A1(KEYINPUT72), .A2(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT72), .A2(G125), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(G140), .A3(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(G125), .A2(G140), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n204), .B1(new_n210), .B2(new_n203), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT82), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT82), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n213), .B(new_n204), .C1(new_n210), .C2(new_n203), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n201), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n197), .ZN(new_n216));
  AOI21_X1  g030(.A(G143), .B1(new_n196), .B2(G214), .ZN(new_n217));
  OAI21_X1  g031(.A(G131), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n219));
  INV_X1    g033(.A(G131), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n195), .A2(new_n220), .A3(new_n197), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT85), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n218), .A2(KEYINPUT85), .A3(new_n219), .A4(new_n221), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n198), .A2(KEYINPUT17), .A3(G131), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT16), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n228), .B1(new_n207), .B2(new_n209), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT72), .A2(G125), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT72), .A2(G125), .ZN(new_n231));
  NOR4_X1   g045(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT16), .A4(G140), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n203), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n230), .A2(new_n231), .ZN(new_n234));
  INV_X1    g048(.A(G140), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n228), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n208), .B1(new_n234), .B2(G140), .ZN(new_n237));
  OAI211_X1 g051(.A(G146), .B(new_n236), .C1(new_n237), .C2(new_n228), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT73), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n233), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  OAI211_X1 g054(.A(KEYINPUT73), .B(new_n203), .C1(new_n229), .C2(new_n232), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI211_X1 g056(.A(new_n190), .B(new_n215), .C1(new_n227), .C2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n215), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n218), .A2(new_n221), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n238), .A2(KEYINPUT74), .ZN(new_n246));
  INV_X1    g060(.A(new_n229), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT74), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n247), .A2(new_n248), .A3(G146), .A4(new_n236), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n207), .A2(KEYINPUT19), .A3(new_n209), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT19), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n202), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n203), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT83), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT83), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n250), .A2(new_n255), .A3(new_n203), .A4(new_n252), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n246), .A2(new_n249), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n245), .B1(new_n257), .B2(KEYINPUT84), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n246), .A2(new_n249), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n254), .A2(new_n256), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n259), .A2(KEYINPUT84), .A3(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n244), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n243), .B1(new_n262), .B2(new_n190), .ZN(new_n263));
  NOR2_X1   g077(.A1(G475), .A2(G902), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT20), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT20), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT84), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n232), .B1(new_n210), .B2(KEYINPUT16), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n248), .B1(new_n269), .B2(G146), .ZN(new_n270));
  NOR4_X1   g084(.A1(new_n229), .A2(new_n232), .A3(KEYINPUT74), .A4(new_n203), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n254), .A2(new_n256), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n268), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n257), .A2(KEYINPUT84), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n245), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n189), .B1(new_n276), .B2(new_n244), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n267), .B(new_n264), .C1(new_n277), .C2(new_n243), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n266), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT86), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n227), .A2(new_n242), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n280), .B(new_n190), .C1(new_n281), .C2(new_n215), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n215), .B1(new_n227), .B2(new_n242), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT86), .B1(new_n283), .B2(new_n189), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n243), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(G475), .B1(new_n285), .B2(G902), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n279), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT87), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT87), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n279), .A2(new_n289), .A3(new_n286), .ZN(new_n290));
  INV_X1    g104(.A(G128), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n291), .A2(G143), .ZN(new_n292));
  XOR2_X1   g106(.A(KEYINPUT66), .B(G128), .Z(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G143), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n292), .B1(new_n294), .B2(KEYINPUT13), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n194), .A2(KEYINPUT13), .A3(G128), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n296), .B(KEYINPUT88), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G134), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G134), .ZN(new_n300));
  INV_X1    g114(.A(new_n292), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT66), .B(G128), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n300), .B(new_n301), .C1(new_n302), .C2(new_n194), .ZN(new_n303));
  INV_X1    g117(.A(G122), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G116), .ZN(new_n305));
  INV_X1    g119(.A(G116), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G122), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n307), .A3(G107), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(new_n307), .ZN(new_n309));
  INV_X1    g123(.A(G107), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n303), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n299), .A2(KEYINPUT89), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT89), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n302), .A2(new_n194), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT13), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n301), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n300), .B1(new_n318), .B2(new_n297), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n315), .B1(new_n319), .B2(new_n312), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n310), .B1(new_n305), .B2(KEYINPUT14), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(new_n309), .ZN(new_n323));
  OAI21_X1  g137(.A(G134), .B1(new_n316), .B2(new_n292), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n303), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT90), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n323), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(KEYINPUT90), .A3(new_n303), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT9), .B(G234), .Z(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(G217), .A3(new_n192), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n321), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n332), .B1(new_n321), .B2(new_n329), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G478), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(KEYINPUT15), .ZN(new_n337));
  OR3_X1    g151(.A1(new_n335), .A2(G902), .A3(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n337), .B1(new_n335), .B2(G902), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n192), .A2(G952), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n341), .B1(G234), .B2(G237), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT21), .B(G898), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT91), .ZN(new_n345));
  INV_X1    g159(.A(G902), .ZN(new_n346));
  AOI211_X1 g160(.A(new_n346), .B(new_n192), .C1(G234), .C2(G237), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n343), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n340), .A2(new_n350), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n288), .A2(new_n290), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT2), .B(G113), .ZN(new_n353));
  INV_X1    g167(.A(G119), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G116), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n306), .A2(G119), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT68), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT68), .B1(new_n355), .B2(new_n356), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n353), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n355), .A2(new_n356), .ZN(new_n360));
  OR2_X1    g174(.A1(new_n360), .A2(new_n353), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT11), .B1(new_n300), .B2(G137), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT11), .ZN(new_n365));
  INV_X1    g179(.A(G137), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n366), .A3(G134), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n300), .A2(G137), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G131), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n220), .A3(new_n369), .ZN(new_n372));
  XNOR2_X1  g186(.A(G143), .B(G146), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(KEYINPUT0), .A2(G128), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT0), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(new_n291), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n374), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n373), .B1(new_n376), .B2(new_n291), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n371), .A2(new_n372), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n291), .A2(KEYINPUT1), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n203), .A2(G143), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n194), .A2(G146), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT65), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n383), .A2(KEYINPUT65), .A3(KEYINPUT1), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(new_n302), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n374), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT67), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(KEYINPUT67), .A3(new_n374), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n386), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT64), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n369), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n300), .B2(G137), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n369), .A2(new_n397), .ZN(new_n400));
  OAI21_X1  g214(.A(G131), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n372), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n363), .B(new_n381), .C1(new_n396), .C2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT28), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n391), .A2(KEYINPUT67), .A3(new_n374), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT67), .B1(new_n391), .B2(new_n374), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n385), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n402), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n363), .B1(new_n410), .B2(new_n381), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT69), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n403), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n410), .A2(KEYINPUT69), .A3(new_n363), .A4(new_n381), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n405), .B1(new_n415), .B2(new_n404), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n196), .A2(G210), .ZN(new_n417));
  INV_X1    g231(.A(G101), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n417), .B(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n420));
  XOR2_X1   g234(.A(new_n419), .B(new_n420), .Z(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT30), .B1(new_n410), .B2(new_n381), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT30), .ZN(new_n425));
  AOI211_X1 g239(.A(new_n425), .B(new_n380), .C1(new_n408), .C2(new_n409), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n427), .A2(new_n362), .B1(new_n413), .B2(new_n414), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT70), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT31), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n428), .A2(new_n429), .A3(new_n430), .A4(new_n421), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n381), .B1(new_n396), .B2(new_n402), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n425), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n410), .A2(KEYINPUT30), .A3(new_n381), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n362), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n413), .A2(new_n414), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n435), .A2(new_n436), .A3(new_n429), .A4(new_n421), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT31), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n423), .A2(new_n431), .A3(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(G472), .A2(G902), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT32), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(KEYINPUT32), .A3(new_n440), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n405), .B(new_n421), .C1(new_n415), .C2(new_n404), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n435), .A2(new_n436), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n422), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT29), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n445), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n421), .B1(new_n415), .B2(new_n404), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT71), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n403), .A2(new_n451), .A3(new_n404), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n451), .B1(new_n403), .B2(new_n404), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT29), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n346), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(G472), .B1(new_n449), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n443), .A2(new_n444), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G469), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n418), .A2(KEYINPUT77), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT77), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G101), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n310), .A3(G104), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n188), .A2(G107), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT3), .B1(new_n188), .B2(G107), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n462), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n310), .A2(G104), .ZN(new_n468));
  OAI211_X1 g282(.A(KEYINPUT78), .B(G101), .C1(new_n465), .C2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT78), .ZN(new_n470));
  XNOR2_X1  g284(.A(G104), .B(G107), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n470), .B1(new_n471), .B2(new_n418), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n467), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n408), .A2(KEYINPUT10), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n464), .B1(new_n466), .B2(new_n465), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(new_n467), .A3(KEYINPUT4), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n378), .A2(new_n379), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT4), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n475), .A2(new_n479), .A3(G101), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n291), .B1(new_n383), .B2(KEYINPUT1), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n385), .B1(new_n482), .B2(new_n373), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n483), .A2(new_n467), .A3(new_n472), .A4(new_n469), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT10), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n371), .A2(new_n372), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT79), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n474), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT80), .ZN(new_n491));
  XNOR2_X1  g305(.A(G110), .B(G140), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n192), .A2(G227), .ZN(new_n493));
  XOR2_X1   g307(.A(new_n492), .B(new_n493), .Z(new_n494));
  AND3_X1   g308(.A1(new_n490), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n467), .A2(new_n469), .A3(new_n472), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n385), .B(new_n496), .C1(new_n406), .C2(new_n407), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n484), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT12), .B1(new_n498), .B2(new_n488), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT12), .ZN(new_n500));
  INV_X1    g314(.A(new_n488), .ZN(new_n501));
  AOI211_X1 g315(.A(new_n500), .B(new_n501), .C1(new_n497), .C2(new_n484), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n491), .B1(new_n490), .B2(new_n494), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n495), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n474), .A2(new_n487), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n488), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n494), .B1(new_n507), .B2(new_n490), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n458), .B(new_n346), .C1(new_n505), .C2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n458), .A2(new_n346), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n494), .ZN(new_n512));
  INV_X1    g326(.A(new_n490), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n512), .B1(new_n503), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n507), .A2(new_n490), .A3(new_n494), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(G469), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n509), .A2(new_n511), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G221), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n330), .B2(new_n346), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(G214), .B1(G237), .B2(G902), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(G210), .B1(G237), .B2(G902), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT68), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n360), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT68), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(KEYINPUT5), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(G113), .B1(new_n355), .B2(KEYINPUT5), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n473), .A2(new_n361), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n362), .A2(new_n477), .A3(new_n480), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(G110), .B(G122), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(KEYINPUT6), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT6), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n534), .A2(new_n540), .A3(new_n536), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n192), .A2(G224), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n234), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n408), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n545), .B1(new_n378), .B2(new_n379), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n544), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  AOI211_X1 g363(.A(new_n543), .B(new_n547), .C1(new_n408), .C2(new_n545), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n542), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n531), .A2(new_n361), .A3(new_n496), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT5), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n361), .B1(new_n554), .B2(new_n529), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n473), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n535), .B(KEYINPUT8), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n553), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n548), .B1(new_n396), .B2(new_n234), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT7), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n544), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n538), .B(new_n558), .C1(new_n559), .C2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n547), .B1(new_n408), .B2(new_n545), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n563), .A2(new_n560), .A3(new_n544), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n346), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n524), .B1(new_n552), .B2(new_n565), .ZN(new_n566));
  AOI211_X1 g380(.A(new_n561), .B(new_n547), .C1(new_n408), .C2(new_n545), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n538), .A2(new_n558), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n559), .A2(KEYINPUT7), .A3(new_n543), .ZN(new_n570));
  AOI21_X1  g384(.A(G902), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n539), .B(new_n541), .C1(new_n549), .C2(new_n550), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n523), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n522), .B1(new_n566), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n517), .A2(new_n520), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT22), .B(G137), .ZN(new_n577));
  INV_X1    g391(.A(G234), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n518), .A2(new_n578), .A3(G953), .ZN(new_n579));
  XOR2_X1   g393(.A(new_n577), .B(new_n579), .Z(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n354), .A2(KEYINPUT23), .A3(G128), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n291), .A2(G119), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n293), .B2(G119), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n582), .B1(new_n584), .B2(KEYINPUT23), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT24), .B(G110), .Z(new_n586));
  OAI22_X1  g400(.A1(new_n585), .A2(G110), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n259), .A2(new_n587), .A3(new_n204), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT75), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n585), .A2(G110), .B1(new_n584), .B2(new_n586), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(new_n241), .A3(new_n240), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n588), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n589), .B1(new_n588), .B2(new_n591), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n581), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n588), .A2(new_n591), .A3(new_n580), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n346), .A3(new_n595), .ZN(new_n596));
  OR2_X1    g410(.A1(new_n596), .A2(KEYINPUT25), .ZN(new_n597));
  OAI21_X1  g411(.A(G217), .B1(new_n578), .B2(G902), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n596), .B2(KEYINPUT25), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT76), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n594), .A2(new_n595), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n598), .A2(new_n346), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n603), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n594), .A2(KEYINPUT76), .A3(new_n595), .A4(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n600), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n352), .A2(new_n457), .A3(new_n576), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT92), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(new_n462), .ZN(G3));
  NAND4_X1  g425(.A1(new_n571), .A2(KEYINPUT93), .A3(new_n523), .A4(new_n572), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n612), .A2(new_n521), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT93), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n566), .A2(new_n614), .A3(new_n573), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n613), .A2(new_n615), .A3(new_n349), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT96), .B(G478), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n335), .B2(G902), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT95), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT94), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n314), .A2(new_n320), .B1(new_n328), .B2(new_n327), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n620), .B1(new_n621), .B2(new_n332), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n622), .B(KEYINPUT33), .C1(new_n333), .C2(new_n334), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n321), .A2(new_n329), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n331), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n621), .A2(new_n332), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n625), .B(new_n626), .C1(new_n620), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n336), .A2(G902), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n619), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n630), .ZN(new_n632));
  AOI211_X1 g446(.A(KEYINPUT95), .B(new_n632), .C1(new_n623), .C2(new_n628), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n618), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n279), .A2(new_n289), .A3(new_n286), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n289), .B1(new_n279), .B2(new_n286), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n616), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(KEYINPUT97), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n288), .A2(new_n290), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT97), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n639), .A2(new_n640), .A3(new_n634), .A4(new_n616), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n517), .A2(new_n520), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n441), .ZN(new_n645));
  INV_X1    g459(.A(G472), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n439), .B2(new_n346), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n642), .A2(new_n608), .A3(new_n644), .A4(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT34), .B(G104), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT98), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n649), .B(new_n651), .ZN(G6));
  NOR2_X1   g466(.A1(new_n607), .A2(new_n350), .ZN(new_n653));
  INV_X1    g467(.A(new_n340), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n287), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n613), .A2(new_n615), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n656), .A2(new_n644), .A3(new_n658), .A4(new_n648), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT35), .B(G107), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  NOR3_X1   g475(.A1(new_n575), .A2(new_n645), .A3(new_n647), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n592), .A2(new_n593), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n581), .A2(KEYINPUT36), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n663), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n605), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n600), .A2(new_n667), .ZN(new_n668));
  AND4_X1   g482(.A1(new_n288), .A2(new_n668), .A3(new_n290), .A4(new_n351), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n662), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  INV_X1    g486(.A(G900), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n342), .B1(new_n347), .B2(new_n673), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n287), .A2(new_n654), .A3(new_n674), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n675), .A2(new_n668), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n676), .A2(new_n457), .A3(new_n644), .A4(new_n658), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XOR2_X1   g492(.A(new_n674), .B(KEYINPUT39), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n644), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n680), .B(KEYINPUT40), .Z(new_n681));
  NAND2_X1  g495(.A1(new_n446), .A2(new_n421), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n415), .A2(new_n422), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n682), .A2(new_n346), .A3(new_n683), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n443), .B(new_n444), .C1(new_n646), .C2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n654), .B1(new_n288), .B2(new_n290), .ZN(new_n686));
  AOI22_X1  g500(.A1(new_n597), .A2(new_n599), .B1(new_n605), .B2(new_n666), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n566), .A2(new_n573), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(new_n690));
  AND4_X1   g504(.A1(new_n521), .A2(new_n686), .A3(new_n687), .A4(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n681), .A2(new_n685), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G143), .ZN(G45));
  AND3_X1   g507(.A1(new_n439), .A2(KEYINPUT32), .A3(new_n440), .ZN(new_n694));
  AOI21_X1  g508(.A(KEYINPUT32), .B1(new_n439), .B2(new_n440), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n643), .B1(new_n696), .B2(new_n456), .ZN(new_n697));
  INV_X1    g511(.A(new_n674), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n634), .B(new_n698), .C1(new_n635), .C2(new_n636), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n687), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n697), .A2(new_n700), .A3(new_n658), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  INV_X1    g516(.A(KEYINPUT101), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n490), .A2(new_n494), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n498), .A2(new_n488), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n500), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n498), .A2(KEYINPUT12), .A3(new_n488), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n704), .A2(KEYINPUT80), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n495), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n508), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(G469), .B1(new_n710), .B2(G902), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT100), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n712), .A3(new_n509), .ZN(new_n713));
  OAI211_X1 g527(.A(KEYINPUT100), .B(G469), .C1(new_n710), .C2(G902), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n519), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n457), .A2(new_n608), .A3(new_n715), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n642), .A2(new_n703), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n703), .B1(new_n642), .B2(new_n716), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT102), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n719), .B(new_n721), .ZN(G15));
  AOI211_X1 g536(.A(new_n519), .B(new_n657), .C1(new_n713), .C2(new_n714), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(new_n457), .A3(new_n655), .A4(new_n653), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  NAND3_X1  g539(.A1(new_n723), .A2(new_n669), .A3(new_n457), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  XOR2_X1   g541(.A(KEYINPUT104), .B(G472), .Z(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n439), .B2(new_n346), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n411), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n404), .B1(new_n436), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n452), .A2(new_n453), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n422), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n431), .A3(new_n438), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n440), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT103), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(KEYINPUT103), .A3(new_n440), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n731), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n607), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n635), .A2(new_n636), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n743), .A2(new_n350), .A3(new_n654), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n742), .A2(KEYINPUT105), .A3(new_n744), .A4(new_n723), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT105), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n686), .A2(new_n349), .A3(new_n715), .A4(new_n658), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n608), .A2(new_n731), .A3(new_n739), .A4(new_n740), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G122), .ZN(G24));
  INV_X1    g565(.A(new_n699), .ZN(new_n752));
  INV_X1    g566(.A(new_n740), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT103), .B1(new_n736), .B2(new_n440), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n753), .A2(new_n730), .A3(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n752), .A2(new_n723), .A3(new_n755), .A4(new_n668), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G125), .ZN(G27));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n514), .A2(new_n758), .ZN(new_n759));
  OAI211_X1 g573(.A(KEYINPUT106), .B(new_n512), .C1(new_n503), .C2(new_n513), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n759), .A2(G469), .A3(new_n515), .A4(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n509), .A3(new_n511), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n566), .A2(new_n521), .A3(new_n573), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n520), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n699), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n443), .A2(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n444), .A2(new_n456), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n695), .A2(KEYINPUT107), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n765), .A2(new_n770), .A3(new_n608), .ZN(new_n771));
  INV_X1    g585(.A(new_n764), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n457), .A2(new_n608), .A3(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n699), .A2(KEYINPUT42), .ZN(new_n774));
  AOI22_X1  g588(.A1(new_n771), .A2(KEYINPUT42), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G131), .ZN(G33));
  AOI21_X1  g590(.A(new_n607), .B1(new_n696), .B2(new_n456), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(KEYINPUT108), .A3(new_n675), .A4(new_n772), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n457), .A2(new_n772), .A3(new_n608), .A4(new_n675), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT108), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G134), .ZN(G36));
  NAND2_X1  g597(.A1(new_n743), .A2(new_n634), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT43), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n743), .A2(KEYINPUT43), .A3(new_n634), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n648), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n789), .A3(new_n668), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  INV_X1    g607(.A(new_n763), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT45), .B1(new_n514), .B2(new_n515), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n458), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n759), .A2(KEYINPUT45), .A3(new_n515), .A4(new_n760), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n510), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n799), .A2(KEYINPUT46), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(KEYINPUT46), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n509), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n520), .A3(new_n679), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT109), .Z(new_n804));
  NAND2_X1  g618(.A1(new_n795), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g619(.A(KEYINPUT110), .B(G137), .Z(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(G39));
  NAND2_X1  g621(.A1(new_n802), .A2(new_n520), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n808), .A2(KEYINPUT47), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(KEYINPUT47), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n457), .A2(new_n699), .A3(new_n608), .A4(new_n794), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g627(.A(KEYINPUT111), .B(G140), .Z(new_n814));
  XNOR2_X1  g628(.A(new_n813), .B(new_n814), .ZN(G42));
  NOR2_X1   g629(.A1(G952), .A2(G953), .ZN(new_n816));
  XOR2_X1   g630(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n520), .A2(new_n687), .A3(new_n762), .A4(new_n698), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n685), .A2(new_n819), .A3(new_n658), .A4(new_n686), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n701), .A2(new_n677), .A3(new_n756), .A4(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n821), .A2(KEYINPUT52), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n288), .A2(new_n290), .A3(new_n340), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n662), .A3(new_n653), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n826), .A2(new_n609), .A3(new_n670), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n741), .A2(new_n699), .A3(new_n687), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n654), .A2(new_n763), .A3(new_n698), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n829), .A2(new_n287), .A3(new_n687), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n828), .A2(new_n772), .B1(new_n697), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n775), .A2(new_n827), .A3(new_n782), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n822), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n821), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n697), .B(new_n658), .C1(new_n700), .C2(new_n676), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(KEYINPUT114), .A3(new_n756), .A4(new_n820), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n835), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n724), .A2(new_n726), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n750), .B(new_n841), .C1(new_n717), .C2(new_n718), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n840), .B1(new_n749), .B2(new_n745), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n845), .B(KEYINPUT115), .C1(new_n717), .C2(new_n718), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n833), .A2(new_n839), .A3(new_n844), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT53), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n835), .A2(new_n838), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT52), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n842), .A2(new_n832), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .A4(new_n839), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n848), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n850), .A2(new_n851), .A3(new_n839), .ZN(new_n855));
  INV_X1    g669(.A(new_n842), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n775), .A2(new_n827), .A3(new_n782), .A4(new_n831), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n856), .A2(new_n839), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n822), .A2(KEYINPUT53), .ZN(new_n859));
  AOI22_X1  g673(.A1(KEYINPUT53), .A2(new_n855), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n818), .A2(new_n854), .B1(new_n860), .B2(KEYINPUT54), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n343), .B1(new_n786), .B2(new_n787), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n742), .A3(new_n763), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n520), .B1(new_n713), .B2(new_n714), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT118), .Z(new_n868));
  OAI211_X1 g682(.A(new_n865), .B(new_n866), .C1(new_n811), .C2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n690), .A2(new_n521), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n862), .A2(new_n715), .A3(new_n742), .A4(new_n870), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT50), .Z(new_n872));
  AND2_X1   g686(.A1(new_n715), .A2(new_n763), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n668), .A2(new_n862), .A3(new_n755), .A4(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n685), .A2(new_n607), .A3(new_n343), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n875), .A2(new_n873), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n639), .A2(new_n634), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n869), .A2(new_n872), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n823), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n341), .B1(new_n876), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n862), .A2(new_n658), .A3(new_n715), .A4(new_n742), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n770), .A2(new_n608), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n862), .A2(new_n886), .A3(new_n873), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT48), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n885), .A2(new_n888), .A3(KEYINPUT119), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n865), .B(new_n866), .C1(new_n811), .C2(new_n867), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n894), .A2(new_n872), .A3(KEYINPUT51), .A4(new_n878), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n881), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n816), .B1(new_n861), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n713), .A2(new_n714), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT49), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OR4_X1    g715(.A1(new_n607), .A2(new_n784), .A3(new_n519), .A4(new_n522), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT112), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(new_n903), .B2(new_n902), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT113), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  AOI211_X1 g722(.A(new_n690), .B(new_n685), .C1(new_n900), .C2(new_n899), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(KEYINPUT120), .B1(new_n898), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n855), .A2(KEYINPUT53), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n858), .A2(new_n859), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n914), .A2(new_n915), .A3(KEYINPUT54), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n817), .B1(new_n848), .B2(new_n853), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n896), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n913), .B(new_n910), .C1(new_n918), .C2(new_n816), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n912), .A2(new_n919), .ZN(G75));
  NOR2_X1   g734(.A1(new_n192), .A2(G952), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n848), .A2(G902), .A3(new_n853), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT56), .B1(new_n924), .B2(G210), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n542), .B(new_n551), .Z(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT55), .Z(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n922), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT121), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n923), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n848), .A2(KEYINPUT121), .A3(G902), .A4(new_n853), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n524), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n927), .B(KEYINPUT122), .Z(new_n935));
  NOR2_X1   g749(.A1(new_n935), .A2(KEYINPUT56), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n929), .B1(new_n934), .B2(new_n936), .ZN(G51));
  NOR2_X1   g751(.A1(new_n854), .A2(new_n818), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n938), .A2(new_n917), .ZN(new_n939));
  XNOR2_X1  g753(.A(KEYINPUT123), .B(KEYINPUT57), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n511), .B(new_n940), .ZN(new_n941));
  OAI22_X1  g755(.A1(new_n939), .A2(new_n941), .B1(new_n508), .B2(new_n505), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n933), .A2(new_n798), .A3(new_n797), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n921), .B1(new_n942), .B2(new_n943), .ZN(G54));
  NAND2_X1  g758(.A1(KEYINPUT58), .A2(G475), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n931), .B2(new_n932), .ZN(new_n946));
  INV_X1    g760(.A(new_n263), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n922), .B1(new_n946), .B2(new_n947), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(G60));
  XNOR2_X1  g764(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n336), .A2(new_n346), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n916), .B2(new_n917), .ZN(new_n955));
  INV_X1    g769(.A(new_n629), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n921), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n956), .A2(new_n953), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n938), .B2(new_n917), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT125), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n961), .B(new_n958), .C1(new_n938), .C2(new_n917), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n957), .A2(new_n960), .A3(new_n962), .ZN(G63));
  XNOR2_X1  g777(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n854), .ZN(new_n966));
  NAND2_X1  g780(.A1(G217), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT60), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n970), .A2(new_n602), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n966), .A2(new_n666), .A3(new_n969), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n922), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n965), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n970), .A2(new_n602), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n975), .A2(new_n922), .A3(new_n972), .A4(new_n964), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(G66));
  AOI21_X1  g791(.A(new_n192), .B1(new_n345), .B2(G224), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n856), .A2(new_n827), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n978), .B1(new_n979), .B2(new_n192), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n542), .B1(G898), .B2(new_n192), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n980), .B(new_n981), .Z(G69));
  AOI21_X1  g796(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n250), .A2(new_n252), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n427), .B(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT127), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n743), .A2(new_n654), .A3(new_n657), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n804), .A2(new_n886), .A3(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n837), .A2(new_n756), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n988), .A2(new_n775), .A3(new_n782), .A4(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  AOI22_X1  g805(.A1(new_n795), .A2(new_n804), .B1(new_n811), .B2(new_n812), .ZN(new_n992));
  AOI21_X1  g806(.A(G953), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n192), .A2(G900), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n986), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n805), .A2(new_n813), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n192), .B1(new_n996), .B2(new_n990), .ZN(new_n997));
  INV_X1    g811(.A(new_n994), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n997), .A2(KEYINPUT127), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n985), .B1(new_n995), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n985), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n692), .A2(new_n989), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT62), .Z(new_n1003));
  NOR2_X1   g817(.A1(new_n680), .A2(new_n794), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1004), .A2(new_n777), .A3(new_n825), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1003), .A2(new_n1005), .A3(new_n992), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1001), .B1(new_n1006), .B2(new_n192), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n983), .B1(new_n1000), .B2(new_n1007), .ZN(new_n1008));
  NOR3_X1   g822(.A1(new_n993), .A2(new_n986), .A3(new_n994), .ZN(new_n1009));
  AOI21_X1  g823(.A(KEYINPUT127), .B1(new_n997), .B2(new_n998), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1001), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n983), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1007), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1008), .A2(new_n1014), .ZN(G72));
  NAND2_X1  g829(.A1(G472), .A2(G902), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT63), .Z(new_n1017));
  OAI21_X1  g831(.A(new_n1017), .B1(new_n1006), .B2(new_n979), .ZN(new_n1018));
  INV_X1    g832(.A(new_n682), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n921), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n996), .A2(new_n979), .A3(new_n990), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1017), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n422), .B(new_n428), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n428), .A2(new_n421), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1022), .B1(new_n1025), .B2(new_n447), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1024), .B1(new_n860), .B2(new_n1026), .ZN(G57));
endmodule


