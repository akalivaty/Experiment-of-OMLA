//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1162, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  XOR2_X1   g019(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n463), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(G101), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT68), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n469), .A2(new_n465), .A3(G101), .A4(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n463), .A2(new_n465), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n466), .A2(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n465), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n465), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n482), .B1(G136), .B2(new_n486), .ZN(new_n487));
  XOR2_X1   g062(.A(new_n487), .B(KEYINPUT69), .Z(G162));
  NAND2_X1  g063(.A1(new_n478), .A2(G126), .ZN(new_n489));
  AND2_X1   g064(.A1(KEYINPUT70), .A2(G114), .ZN(new_n490));
  NOR2_X1   g065(.A1(KEYINPUT70), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2105), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n497), .A2(new_n465), .A3(G138), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n485), .A2(KEYINPUT71), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR3_X1   g076(.A1(new_n501), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n500), .B1(new_n463), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g079(.A(G138), .B(new_n465), .C1(new_n483), .C2(new_n484), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n496), .B1(new_n504), .B2(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT72), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT72), .A2(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  OAI211_X1 g092(.A(G88), .B(new_n512), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT72), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT72), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n524));
  OAI21_X1  g099(.A(KEYINPUT6), .B1(new_n519), .B2(new_n520), .ZN(new_n525));
  INV_X1    g100(.A(new_n517), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n509), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n524), .B1(new_n527), .B2(G50), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n527), .A2(new_n524), .A3(G50), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n523), .B1(new_n529), .B2(new_n530), .ZN(G166));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT74), .ZN(new_n533));
  XOR2_X1   g108(.A(new_n533), .B(KEYINPUT7), .Z(new_n534));
  AOI21_X1  g109(.A(new_n534), .B1(G51), .B2(new_n527), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n510), .A2(new_n511), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n536), .B1(new_n526), .B2(new_n525), .ZN(new_n537));
  AND2_X1   g112(.A1(G63), .A2(G651), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n537), .A2(G89), .B1(new_n512), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n535), .A2(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n536), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n521), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n544), .A2(new_n545), .B1(new_n527), .B2(G52), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n537), .A2(G90), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(G171));
  AOI22_X1  g124(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n521), .ZN(new_n551));
  XOR2_X1   g126(.A(new_n551), .B(KEYINPUT75), .Z(new_n552));
  AOI22_X1  g127(.A1(new_n537), .A2(G81), .B1(new_n527), .B2(G43), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT76), .Z(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(new_n537), .A2(G91), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n512), .A2(KEYINPUT77), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n510), .A2(new_n563), .A3(new_n511), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G651), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n561), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n527), .A2(G53), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(G299));
  XNOR2_X1  g147(.A(new_n548), .B(KEYINPUT78), .ZN(G301));
  NAND2_X1  g148(.A1(G75), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G62), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n536), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(new_n545), .ZN(new_n577));
  INV_X1    g152(.A(new_n530), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n518), .B(new_n577), .C1(new_n578), .C2(new_n528), .ZN(G303));
  NAND2_X1  g154(.A1(new_n537), .A2(G87), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n527), .A2(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(G48), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n525), .B2(new_n526), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n536), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n537), .A2(G86), .B1(new_n590), .B2(new_n545), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n537), .A2(G85), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  INV_X1    g169(.A(new_n527), .ZN(new_n595));
  XOR2_X1   g170(.A(KEYINPUT80), .B(G47), .Z(new_n596));
  OAI221_X1 g171(.A(new_n593), .B1(new_n521), .B2(new_n594), .C1(new_n595), .C2(new_n596), .ZN(G290));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n562), .B2(new_n564), .ZN(new_n599));
  AND2_X1   g174(.A1(G79), .A2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n527), .A2(G54), .ZN(new_n602));
  AND2_X1   g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n537), .A2(G92), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n537), .A2(KEYINPUT10), .A3(G92), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G301), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G284));
  AOI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G321));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(G299), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G168), .B2(new_n614), .ZN(G297));
  XOR2_X1   g191(.A(G297), .B(KEYINPUT81), .Z(G280));
  INV_X1    g192(.A(new_n609), .ZN(new_n618));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n552), .A2(new_n553), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(new_n614), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n609), .A2(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n614), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n486), .A2(G135), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT82), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT83), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(G111), .ZN(new_n631));
  AOI22_X1  g206(.A1(new_n628), .A2(new_n629), .B1(new_n631), .B2(G2105), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n630), .A2(new_n632), .B1(new_n478), .B2(G123), .ZN(new_n633));
  AND2_X1   g208(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n635), .A2(G2096), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n640), .A2(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(G2100), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n635), .A2(G2096), .ZN(new_n643));
  NAND4_X1  g218(.A1(new_n636), .A2(new_n641), .A3(new_n642), .A4(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(KEYINPUT14), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n656));
  XNOR2_X1  g231(.A(G2451), .B(G2454), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(G14), .B1(new_n655), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n660), .B1(new_n659), .B2(new_n655), .ZN(G401));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT85), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT17), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2084), .B(G2090), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n666), .B1(new_n663), .B2(new_n665), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n664), .B2(new_n665), .ZN(new_n669));
  INV_X1    g244(.A(new_n665), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n670), .A2(new_n666), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n663), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT18), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n667), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1956), .B(G2474), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT86), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT20), .Z(new_n685));
  OR2_X1    g260(.A1(new_n678), .A2(new_n680), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n686), .A2(new_n683), .A3(new_n681), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n685), .B(new_n687), .C1(new_n683), .C2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT87), .B(KEYINPUT88), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n692), .B(new_n695), .ZN(G229));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G21), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G168), .B2(new_n697), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n699), .A2(G1966), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT95), .ZN(new_n701));
  INV_X1    g276(.A(G1961), .ZN(new_n702));
  NOR2_X1   g277(.A1(G171), .A2(new_n697), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G5), .B2(new_n697), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n699), .A2(G1966), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT89), .B(G29), .Z(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(G27), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G164), .B2(new_n707), .ZN(new_n709));
  INV_X1    g284(.A(G2078), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n705), .B(new_n711), .C1(new_n702), .C2(new_n704), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n701), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n486), .A2(G141), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT93), .ZN(new_n715));
  AND3_X1   g290(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n716));
  NAND3_X1  g291(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT26), .ZN(new_n718));
  AOI211_X1 g293(.A(new_n716), .B(new_n718), .C1(G129), .C2(new_n478), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n722), .B2(G32), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT27), .B(G1996), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT94), .Z(new_n727));
  NOR2_X1   g302(.A1(G29), .A2(G33), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT25), .ZN(new_n730));
  NAND2_X1  g305(.A1(G115), .A2(G2104), .ZN(new_n731));
  INV_X1    g306(.A(G127), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n485), .B2(new_n732), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n733), .A2(G2105), .ZN(new_n734));
  AOI211_X1 g309(.A(new_n730), .B(new_n734), .C1(G139), .C2(new_n486), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n728), .B1(new_n735), .B2(G29), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT92), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G2072), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT31), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(G11), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(G11), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT30), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n742), .A2(G28), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n722), .B1(new_n742), .B2(G28), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n740), .B(new_n741), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT24), .B(G34), .ZN(new_n746));
  AOI22_X1  g321(.A1(G160), .A2(G29), .B1(new_n706), .B2(new_n746), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n747), .A2(G2084), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n745), .B(new_n748), .C1(new_n634), .C2(new_n707), .ZN(new_n749));
  OAI221_X1 g324(.A(new_n749), .B1(G2084), .B2(new_n747), .C1(new_n724), .C2(new_n725), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n738), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n713), .A2(new_n727), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT96), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n697), .A2(G20), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT23), .Z(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G299), .B2(G16), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1956), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n707), .A2(G35), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G162), .B2(new_n707), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT29), .Z(new_n760));
  INV_X1    g335(.A(G2090), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT97), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n760), .A2(new_n761), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n697), .A2(G19), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n554), .B2(new_n697), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1341), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n697), .A2(G4), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n618), .B2(new_n697), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1348), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n706), .A2(G26), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT28), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n486), .A2(G140), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n478), .A2(G128), .ZN(new_n776));
  OR2_X1    g351(.A1(G104), .A2(G2105), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n777), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n774), .B1(new_n780), .B2(new_n722), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2067), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n769), .A2(new_n772), .A3(new_n782), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n764), .A2(new_n765), .A3(new_n766), .A4(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n753), .A2(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G6), .B(G305), .S(G16), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT32), .ZN(new_n787));
  INV_X1    g362(.A(G1981), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n697), .A2(G23), .ZN(new_n790));
  INV_X1    g365(.A(G288), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(new_n697), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT33), .B(G1976), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n697), .A2(G22), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G166), .B2(new_n697), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n796), .A2(G1971), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n796), .A2(G1971), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n794), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n789), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(KEYINPUT34), .ZN(new_n801));
  MUX2_X1   g376(.A(G24), .B(G290), .S(G16), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G1986), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n707), .A2(G25), .ZN(new_n804));
  OAI21_X1  g379(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G107), .B2(new_n465), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT90), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n486), .A2(G131), .B1(G119), .B2(new_n478), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n804), .B1(new_n810), .B2(new_n707), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT35), .B(G1991), .Z(new_n812));
  XOR2_X1   g387(.A(new_n811), .B(new_n812), .Z(new_n813));
  NOR2_X1   g388(.A1(new_n802), .A2(G1986), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n813), .A2(KEYINPUT91), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n801), .A2(new_n803), .A3(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT36), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n800), .A2(KEYINPUT34), .ZN(new_n818));
  OR3_X1    g393(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n817), .B1(new_n816), .B2(new_n818), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n785), .A2(new_n819), .A3(new_n820), .ZN(G150));
  INV_X1    g396(.A(G150), .ZN(G311));
  AOI22_X1  g397(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(new_n521), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n537), .A2(G93), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n527), .A2(G55), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G860), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT100), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT37), .ZN(new_n830));
  INV_X1    g405(.A(new_n827), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n554), .A2(KEYINPUT99), .A3(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n831), .A2(KEYINPUT99), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(KEYINPUT99), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n833), .A2(new_n621), .A3(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n618), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n842));
  INV_X1    g417(.A(G860), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n841), .B2(KEYINPUT39), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n830), .B1(new_n842), .B2(new_n844), .ZN(G145));
  XNOR2_X1  g420(.A(G162), .B(G160), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n635), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT71), .B1(new_n485), .B2(new_n498), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n463), .A2(new_n500), .A3(new_n502), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n506), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AOI22_X1  g425(.A1(G126), .A2(new_n478), .B1(new_n492), .B2(new_n494), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n779), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n721), .B(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n735), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n478), .A2(G130), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n465), .A2(G118), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n858));
  INV_X1    g433(.A(G142), .ZN(new_n859));
  OAI221_X1 g434(.A(new_n856), .B1(new_n857), .B2(new_n858), .C1(new_n859), .C2(new_n472), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT101), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n638), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n810), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT102), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n855), .A2(new_n863), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT103), .Z(new_n867));
  OAI21_X1  g442(.A(new_n847), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n864), .B(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n847), .B1(new_n855), .B2(new_n863), .ZN(new_n871));
  AOI21_X1  g446(.A(G37), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g449(.A1(new_n827), .A2(new_n614), .ZN(new_n875));
  XNOR2_X1  g450(.A(G166), .B(G305), .ZN(new_n876));
  XNOR2_X1  g451(.A(G290), .B(G288), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT42), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT106), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n878), .B(KEYINPUT105), .Z(new_n882));
  OAI21_X1  g457(.A(new_n881), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n836), .B(new_n623), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n618), .A2(G299), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n609), .A2(new_n571), .A3(new_n569), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n886), .B(KEYINPUT104), .Z(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n885), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(new_n618), .B2(G299), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n891), .A2(new_n892), .B1(new_n886), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n889), .B1(new_n894), .B2(new_n884), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n883), .B(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n875), .B1(new_n896), .B2(new_n614), .ZN(G295));
  OAI21_X1  g472(.A(new_n875), .B1(new_n896), .B2(new_n614), .ZN(G331));
  INV_X1    g473(.A(new_n882), .ZN(new_n899));
  NAND2_X1  g474(.A1(G286), .A2(new_n548), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(G286), .B2(G301), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n836), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n901), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n832), .A2(new_n835), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n888), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n890), .A2(new_n893), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(KEYINPUT41), .B2(new_n887), .ZN(new_n909));
  INV_X1    g484(.A(new_n906), .ZN(new_n910));
  AOI22_X1  g485(.A1(KEYINPUT107), .A2(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n907), .A2(KEYINPUT107), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n899), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(G37), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n907), .B1(new_n894), .B2(new_n906), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n914), .B1(new_n915), .B2(new_n882), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n913), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n887), .B1(new_n902), .B2(new_n905), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n891), .A2(new_n892), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n893), .A2(new_n886), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n919), .B1(new_n922), .B2(new_n910), .ZN(new_n923));
  AOI21_X1  g498(.A(G37), .B1(new_n923), .B2(new_n899), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n915), .A2(new_n882), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT43), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT44), .B1(new_n918), .B2(new_n926), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n913), .A2(new_n916), .A3(KEYINPUT43), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n917), .B1(new_n924), .B2(new_n925), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n927), .B1(new_n930), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n932));
  INV_X1    g507(.A(G1384), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n932), .B1(new_n852), .B2(new_n933), .ZN(new_n934));
  AOI211_X1 g509(.A(KEYINPUT109), .B(G1384), .C1(new_n850), .C2(new_n851), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT50), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n486), .A2(G137), .B1(new_n468), .B2(new_n470), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n937), .B(G40), .C1(new_n465), .C2(new_n464), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT50), .ZN(new_n939));
  AOI21_X1  g514(.A(G1384), .B1(new_n850), .B2(new_n851), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(G1956), .B1(new_n936), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n852), .A2(new_n933), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n938), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n940), .A2(KEYINPUT45), .ZN(new_n946));
  XOR2_X1   g521(.A(KEYINPUT56), .B(G2072), .Z(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT115), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n942), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g525(.A(new_n570), .B(KEYINPUT9), .Z(new_n951));
  OAI21_X1  g526(.A(KEYINPUT57), .B1(new_n951), .B2(new_n568), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT57), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n569), .A2(new_n953), .A3(new_n571), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n950), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT109), .B1(G164), .B2(G1384), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n940), .A2(new_n932), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n939), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G40), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n466), .A2(new_n474), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(new_n940), .B2(new_n939), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(G1348), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n958), .A2(new_n962), .A3(new_n959), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n966), .A2(G2067), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(new_n609), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT116), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n955), .B(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n950), .ZN(new_n972));
  AOI22_X1  g547(.A1(new_n957), .A2(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n944), .B1(G164), .B2(G1384), .ZN(new_n974));
  INV_X1    g549(.A(G1996), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n974), .A2(new_n975), .A3(new_n946), .A4(new_n962), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT117), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n945), .A2(KEYINPUT117), .A3(new_n975), .A4(new_n946), .ZN(new_n979));
  XOR2_X1   g554(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(G1341), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n966), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n978), .A2(new_n979), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n554), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT59), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT60), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(new_n965), .B2(new_n967), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n603), .A2(KEYINPUT120), .A3(new_n608), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n989), .A2(KEYINPUT60), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n934), .A2(new_n935), .ZN(new_n991));
  INV_X1    g566(.A(G2067), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(new_n992), .A3(new_n962), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n963), .B1(new_n991), .B2(new_n939), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n990), .B(new_n993), .C1(new_n994), .C2(G1348), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT120), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n609), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n988), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT61), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(KEYINPUT119), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(new_n950), .B2(new_n956), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1000), .ZN(new_n1002));
  NOR4_X1   g577(.A1(new_n942), .A2(new_n955), .A3(new_n949), .A4(new_n1002), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n986), .B(new_n998), .C1(new_n1001), .C2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n972), .A2(new_n999), .A3(new_n955), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n968), .A2(new_n996), .A3(KEYINPUT60), .A4(new_n609), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n983), .A2(KEYINPUT59), .A3(new_n554), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n973), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n960), .A2(new_n761), .A3(new_n964), .ZN(new_n1010));
  INV_X1    g585(.A(G1971), .ZN(new_n1011));
  INV_X1    g586(.A(new_n946), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n962), .B1(new_n940), .B2(KEYINPUT45), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT110), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n1017));
  INV_X1    g592(.A(G8), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(G166), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1019), .A2(new_n1020), .A3(KEYINPUT111), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT111), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1010), .A2(new_n1024), .A3(new_n1014), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1016), .A2(G8), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT49), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n537), .A2(G86), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n590), .A2(new_n545), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n525), .A2(new_n526), .ZN(new_n1031));
  INV_X1    g606(.A(new_n584), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n586), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI211_X1 g608(.A(KEYINPUT79), .B(new_n584), .C1(new_n525), .C2(new_n526), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1030), .A2(new_n1035), .A3(G1981), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n788), .B1(new_n587), .B2(new_n591), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1027), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(G1981), .B1(new_n1030), .B2(new_n1035), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n587), .A2(new_n591), .A3(new_n788), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(new_n1040), .A3(KEYINPUT49), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n966), .A2(G8), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT113), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1018), .B1(new_n991), .B2(new_n962), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1045), .A2(new_n1046), .A3(new_n1041), .A4(new_n1038), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n791), .A2(G1976), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT52), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G1976), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT112), .B1(G288), .B2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1043), .A2(new_n1051), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1044), .A2(new_n1047), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n936), .A2(new_n761), .A3(new_n941), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1056), .A2(new_n1014), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1055), .B1(new_n1057), .B2(new_n1018), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1026), .A2(new_n1053), .A3(new_n1054), .A4(new_n1058), .ZN(new_n1059));
  XOR2_X1   g634(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n1060));
  INV_X1    g635(.A(KEYINPUT123), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n945), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1013), .A2(KEYINPUT123), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(G2078), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n946), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n945), .A2(new_n710), .A3(new_n946), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1064), .A2(new_n1067), .B1(new_n1068), .B2(new_n1065), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n960), .A2(new_n964), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(new_n702), .ZN(new_n1072));
  AOI211_X1 g647(.A(KEYINPUT122), .B(G1961), .C1(new_n960), .C2(new_n964), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1069), .B(G301), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(new_n702), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1068), .A2(new_n1065), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n938), .B1(KEYINPUT45), .B2(new_n940), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1077), .B(new_n1066), .C1(new_n991), .C2(KEYINPUT45), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n611), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1060), .B1(new_n1074), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1059), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1077), .B1(new_n991), .B2(KEYINPUT45), .ZN(new_n1083));
  INV_X1    g658(.A(G1966), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G2084), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n960), .A2(new_n1086), .A3(new_n964), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(G168), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G8), .ZN(new_n1089));
  AOI21_X1  g664(.A(G168), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT51), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT51), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(new_n1092), .A3(G8), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1069), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G171), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1075), .A2(G301), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1096), .A2(KEYINPUT54), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1091), .A2(new_n1093), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1009), .A2(new_n1082), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT114), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1025), .A2(G8), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1024), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1016), .A2(KEYINPUT114), .A3(G8), .A4(new_n1025), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1103), .A2(new_n1104), .A3(new_n1055), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1106));
  AOI211_X1 g681(.A(new_n1018), .B(G286), .C1(new_n1085), .C2(new_n1087), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT63), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1110), .A2(new_n1050), .A3(new_n791), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1043), .B1(new_n1111), .B2(new_n1040), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT63), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1107), .A2(new_n1058), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1026), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1112), .B1(new_n1106), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1099), .A2(new_n1109), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT124), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1099), .A2(KEYINPUT124), .A3(new_n1109), .A4(new_n1116), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1059), .A2(new_n1080), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1119), .A2(new_n1120), .A3(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n779), .B(new_n992), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(KEYINPUT108), .ZN(new_n1129));
  AOI211_X1 g704(.A(new_n938), .B(new_n974), .C1(new_n1129), .C2(new_n721), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1129), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1130), .B1(G1996), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n974), .A2(new_n938), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n975), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n721), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n810), .B(new_n812), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n1133), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1132), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(G290), .B(G1986), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1139), .B1(new_n1133), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1127), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1130), .B1(KEYINPUT46), .B2(new_n1135), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT46), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT125), .B1(new_n1134), .B2(new_n1144), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1134), .A2(KEYINPUT125), .A3(new_n1144), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1143), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT47), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1148), .A2(KEYINPUT126), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(KEYINPUT126), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n810), .A2(new_n812), .ZN(new_n1152));
  OAI22_X1  g727(.A1(new_n1151), .A2(new_n1152), .B1(G2067), .B2(new_n779), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1139), .ZN(new_n1154));
  NOR2_X1   g729(.A1(G290), .A2(G1986), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1133), .A2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT48), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1153), .A2(new_n1133), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1149), .A2(new_n1150), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1142), .A2(new_n1159), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g735(.A1(G227), .A2(new_n461), .ZN(new_n1162));
  XOR2_X1   g736(.A(new_n1162), .B(KEYINPUT127), .Z(new_n1163));
  NOR3_X1   g737(.A1(G229), .A2(new_n1163), .A3(G401), .ZN(new_n1164));
  OAI211_X1 g738(.A(new_n1164), .B(new_n873), .C1(new_n928), .C2(new_n929), .ZN(G225));
  INV_X1    g739(.A(G225), .ZN(G308));
endmodule


