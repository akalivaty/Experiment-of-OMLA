//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1215, new_n1216, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT64), .Z(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n210), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT65), .Z(new_n228));
  INV_X1    g0028(.A(KEYINPUT1), .ZN(new_n229));
  AND2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n228), .A2(new_n229), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR3_X1   g0033(.A1(new_n232), .A2(new_n208), .A3(new_n233), .ZN(new_n234));
  NOR4_X1   g0034(.A1(new_n214), .A2(new_n230), .A3(new_n231), .A4(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT66), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n233), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n255), .B1(new_n207), .B2(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G13), .ZN(new_n259));
  NOR3_X1   g0059(.A1(new_n259), .A2(new_n208), .A3(G1), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n258), .B1(new_n260), .B2(new_n253), .ZN(new_n261));
  AND3_X1   g0061(.A1(KEYINPUT74), .A2(G58), .A3(G68), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT74), .B1(G58), .B2(G68), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G58), .A2(G68), .ZN(new_n264));
  NOR3_X1   g0064(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G159), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  OAI22_X1  g0068(.A1(new_n265), .A2(new_n208), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT16), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT73), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT7), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n275));
  INV_X1    g0075(.A(G33), .ZN(new_n276));
  NOR3_X1   g0076(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n273), .B(new_n208), .C1(new_n277), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G68), .ZN(new_n281));
  OR2_X1    g0081(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n282));
  NAND2_X1  g0082(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G33), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(G20), .B1(new_n284), .B2(new_n278), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(new_n273), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n272), .B1(new_n281), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n274), .A2(new_n275), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n279), .B1(new_n288), .B2(G33), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT7), .B1(new_n289), .B2(G20), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n290), .A2(KEYINPUT73), .A3(G68), .A4(new_n280), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n271), .B1(new_n287), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT3), .B(G33), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n273), .B1(new_n293), .B2(G20), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n282), .A2(new_n283), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n295), .B1(new_n296), .B2(new_n276), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n208), .A2(KEYINPUT7), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n294), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n269), .B1(new_n299), .B2(G68), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n255), .B1(new_n300), .B2(KEYINPUT16), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n261), .B1(new_n292), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n303));
  INV_X1    g0103(.A(G274), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n305), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n306), .B1(G232), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(G223), .A2(G1698), .ZN(new_n310));
  INV_X1    g0110(.A(G226), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n310), .B1(new_n311), .B2(G1698), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n289), .A2(new_n312), .B1(G33), .B2(G87), .ZN(new_n313));
  INV_X1    g0113(.A(new_n303), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n309), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G200), .ZN(new_n316));
  INV_X1    g0116(.A(G190), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(new_n315), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n302), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n319), .B(KEYINPUT17), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n302), .A2(KEYINPUT75), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT75), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n322), .B(new_n261), .C1(new_n292), .C2(new_n301), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n315), .A2(G169), .ZN(new_n324));
  INV_X1    g0124(.A(G179), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(new_n315), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n321), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT18), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n328), .A2(KEYINPUT76), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(KEYINPUT76), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n327), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n330), .B1(new_n327), .B2(new_n329), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n331), .A2(new_n332), .A3(KEYINPUT77), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT77), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n321), .A2(new_n323), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n335), .A2(KEYINPUT76), .A3(new_n328), .A4(new_n326), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n327), .A2(new_n329), .A3(new_n330), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n320), .B1(new_n333), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G150), .ZN(new_n340));
  OAI22_X1  g0140(.A1(new_n340), .A2(new_n268), .B1(new_n201), .B2(new_n208), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n208), .A2(G33), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n341), .B1(new_n253), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n255), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G50), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n260), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n257), .B2(new_n347), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G1698), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n293), .A2(G222), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n293), .A2(G1698), .ZN(new_n353));
  INV_X1    g0153(.A(G223), .ZN(new_n354));
  OAI221_X1 g0154(.A(new_n352), .B1(new_n202), .B2(new_n293), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n303), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n306), .B1(G226), .B2(new_n308), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n350), .A2(KEYINPUT9), .B1(G200), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n358), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G190), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n359), .B(new_n361), .C1(KEYINPUT9), .C2(new_n350), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT10), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n362), .B(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G169), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n350), .B1(new_n365), .B2(new_n358), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n360), .A2(new_n325), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n267), .A2(G50), .B1(G20), .B2(new_n216), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n202), .B2(new_n342), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n371), .A2(new_n255), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n372), .A2(KEYINPUT11), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(KEYINPUT11), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n259), .A2(G1), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G20), .ZN(new_n376));
  OR3_X1    g0176(.A1(new_n376), .A2(KEYINPUT12), .A3(G68), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT12), .B1(new_n376), .B2(G68), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n377), .A2(new_n378), .B1(G68), .B2(new_n256), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n373), .A2(new_n374), .A3(new_n379), .ZN(new_n380));
  XOR2_X1   g0180(.A(new_n380), .B(KEYINPUT70), .Z(new_n381));
  INV_X1    g0181(.A(KEYINPUT13), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G97), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n293), .A2(new_n351), .ZN(new_n384));
  OAI221_X1 g0184(.A(new_n383), .B1(new_n384), .B2(new_n311), .C1(new_n223), .C2(new_n353), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n303), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n306), .B1(G238), .B2(new_n308), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n382), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(new_n382), .A3(new_n387), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(G179), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(KEYINPUT69), .A2(G169), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n389), .B2(new_n390), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT14), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n392), .ZN(new_n396));
  INV_X1    g0196(.A(new_n390), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n394), .B(new_n396), .C1(new_n397), .C2(new_n388), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n381), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n389), .A2(new_n390), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G200), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n402), .B(new_n380), .C1(new_n401), .C2(new_n317), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT71), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n293), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G107), .ZN(new_n408));
  OAI221_X1 g0208(.A(new_n408), .B1(new_n384), .B2(new_n223), .C1(new_n217), .C2(new_n353), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n303), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n306), .B1(G244), .B2(new_n308), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n365), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n251), .A2(new_n268), .B1(new_n208), .B2(new_n202), .ZN(new_n414));
  XNOR2_X1  g0214(.A(KEYINPUT15), .B(G87), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n342), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n255), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT67), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n376), .A2(G77), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(G77), .B2(new_n256), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n413), .A2(new_n421), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n422), .A2(KEYINPUT68), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n410), .A2(new_n325), .A3(new_n411), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(KEYINPUT68), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n421), .B1(G200), .B2(new_n412), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n317), .B2(new_n412), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n369), .A2(new_n406), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n400), .A2(KEYINPUT71), .A3(new_n403), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n339), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT84), .ZN(new_n434));
  INV_X1    g0234(.A(G41), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n207), .B(G45), .C1(new_n435), .C2(KEYINPUT5), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT79), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(KEYINPUT5), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n436), .B2(KEYINPUT79), .ZN(new_n440));
  OAI211_X1 g0240(.A(G270), .B(new_n314), .C1(new_n438), .C2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n303), .A2(new_n304), .ZN(new_n442));
  INV_X1    g0242(.A(G45), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(G1), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT79), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n444), .B(new_n445), .C1(KEYINPUT5), .C2(new_n435), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n442), .A2(new_n437), .A3(new_n439), .A4(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n434), .B1(new_n441), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n441), .A2(new_n434), .A3(new_n447), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n284), .A2(new_n278), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G264), .A2(G1698), .ZN(new_n452));
  INV_X1    g0252(.A(G303), .ZN(new_n453));
  OAI22_X1  g0253(.A1(new_n451), .A2(new_n452), .B1(new_n453), .B2(new_n293), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT85), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n225), .A2(G1698), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n289), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n456), .B1(new_n289), .B2(new_n457), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n455), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n449), .A2(new_n450), .B1(new_n461), .B2(new_n303), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G283), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n463), .B(new_n208), .C1(G33), .C2(new_n224), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(new_n255), .C1(new_n208), .C2(G116), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT20), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT86), .B1(new_n465), .B2(new_n466), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n345), .B(new_n376), .C1(G1), .C2(new_n276), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G116), .ZN(new_n471));
  INV_X1    g0271(.A(G116), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n376), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n467), .A2(new_n468), .ZN(new_n476));
  OAI21_X1  g0276(.A(G169), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT21), .B1(new_n462), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n450), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n289), .A2(new_n457), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT85), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n454), .B1(new_n481), .B2(new_n458), .ZN(new_n482));
  OAI22_X1  g0282(.A1(new_n479), .A2(new_n448), .B1(new_n482), .B2(new_n314), .ZN(new_n483));
  INV_X1    g0283(.A(new_n476), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n467), .A2(new_n468), .B1(new_n471), .B2(new_n473), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n365), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT21), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n483), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n325), .B1(new_n484), .B2(new_n485), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n478), .A2(new_n488), .B1(new_n462), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n484), .A2(new_n485), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(new_n483), .B2(G200), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n317), .B2(new_n483), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT80), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n293), .A2(KEYINPUT4), .A3(G244), .A4(new_n351), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n293), .A2(G250), .A3(G1698), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n496), .A2(new_n463), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n351), .A2(G244), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n451), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n314), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n314), .B1(new_n438), .B2(new_n440), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n447), .B1(new_n503), .B2(new_n225), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(G200), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n495), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(KEYINPUT80), .B(G200), .C1(new_n502), .C2(new_n504), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n299), .A2(G107), .ZN(new_n510));
  INV_X1    g0310(.A(G107), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(KEYINPUT6), .A3(G97), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n224), .A2(new_n511), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(new_n204), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n512), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n515), .A2(G20), .B1(G77), .B2(new_n267), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n255), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n260), .A2(new_n224), .ZN(new_n519));
  XNOR2_X1  g0319(.A(new_n519), .B(KEYINPUT78), .ZN(new_n520));
  INV_X1    g0320(.A(new_n470), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(G97), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n502), .A2(new_n504), .A3(new_n317), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n509), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n505), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n527), .A2(new_n365), .B1(new_n518), .B2(new_n522), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n505), .A2(new_n325), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n444), .A2(new_n304), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n219), .B1(new_n443), .B2(G1), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n314), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  MUX2_X1   g0334(.A(G238), .B(G244), .S(G1698), .Z(new_n535));
  NAND2_X1  g0335(.A1(new_n289), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n276), .A2(new_n472), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n534), .B1(new_n539), .B2(new_n303), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT81), .B1(new_n540), .B2(new_n325), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n537), .B1(new_n289), .B2(new_n535), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n533), .B1(new_n542), .B2(new_n314), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT81), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n543), .A2(new_n544), .A3(G179), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n415), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(new_n376), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT19), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n208), .B1(new_n383), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT82), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(KEYINPUT82), .B(new_n208), .C1(new_n383), .C2(new_n549), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n552), .B(new_n553), .C1(G87), .C2(new_n205), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n549), .B1(new_n342), .B2(new_n224), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n289), .A2(new_n208), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n554), .B(new_n555), .C1(new_n556), .C2(new_n216), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n548), .B1(new_n557), .B2(new_n255), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n521), .A2(new_n547), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n558), .A2(new_n559), .B1(new_n365), .B2(new_n543), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n543), .A2(G200), .ZN(new_n561));
  OAI211_X1 g0361(.A(G190), .B(new_n533), .C1(new_n542), .C2(new_n314), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n557), .A2(new_n255), .ZN(new_n564));
  INV_X1    g0364(.A(new_n548), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n521), .A2(KEYINPUT83), .A3(G87), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT83), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n470), .B2(new_n218), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n564), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n546), .A2(new_n560), .B1(new_n563), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n526), .A2(new_n530), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT22), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n208), .A2(G87), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n573), .B1(new_n407), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT23), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n208), .B2(G107), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n511), .A2(KEYINPUT23), .A3(G20), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n577), .A2(new_n578), .B1(new_n537), .B2(new_n208), .ZN(new_n579));
  NAND2_X1  g0379(.A1(KEYINPUT22), .A2(G87), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n575), .B(new_n579), .C1(new_n556), .C2(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n581), .A2(KEYINPUT24), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n581), .A2(KEYINPUT24), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n255), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT25), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n376), .B2(G107), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n260), .A2(KEYINPUT25), .A3(new_n511), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n521), .A2(G107), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(G264), .B(new_n314), .C1(new_n438), .C2(new_n440), .ZN(new_n590));
  NOR2_X1   g0390(.A1(G250), .A2(G1698), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n225), .B2(G1698), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n289), .A2(new_n592), .B1(G33), .B2(G294), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n590), .B1(new_n593), .B2(new_n314), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT87), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n590), .B(KEYINPUT87), .C1(new_n593), .C2(new_n314), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n596), .A2(G179), .A3(new_n447), .A4(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n447), .ZN(new_n599));
  OAI21_X1  g0399(.A(G169), .B1(new_n594), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n589), .A2(new_n601), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n594), .A2(G190), .A3(new_n599), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n596), .A2(new_n447), .A3(new_n597), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n603), .B1(new_n604), .B2(new_n506), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n602), .B1(new_n589), .B2(new_n605), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n494), .A2(new_n572), .A3(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n433), .A2(new_n607), .ZN(G372));
  INV_X1    g0408(.A(new_n368), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n302), .A2(new_n326), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n610), .B(KEYINPUT18), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n403), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n400), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n611), .B1(new_n614), .B2(new_n320), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n609), .B1(new_n615), .B2(new_n364), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n433), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n509), .A2(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n560), .B1(G179), .B2(new_n543), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n570), .A2(new_n563), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n605), .A2(new_n589), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n619), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n478), .A2(new_n488), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n462), .A2(G179), .A3(new_n491), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n602), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT88), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT88), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n490), .A2(new_n630), .A3(new_n602), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n624), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n571), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT26), .B1(new_n633), .B2(new_n530), .ZN(new_n634));
  INV_X1    g0434(.A(new_n530), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n622), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(new_n637), .A3(new_n620), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n617), .B1(new_n618), .B2(new_n639), .ZN(G369));
  INV_X1    g0440(.A(new_n606), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n375), .A2(new_n208), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(G213), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n589), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n641), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n628), .A2(new_n647), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n491), .A2(new_n647), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n490), .A2(new_n493), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n490), .B2(new_n653), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(G330), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n490), .A2(new_n647), .ZN(new_n659));
  INV_X1    g0459(.A(new_n647), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n659), .A2(new_n641), .B1(new_n628), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n658), .A2(new_n661), .ZN(G399));
  INV_X1    g0462(.A(new_n211), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(G41), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G1), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n232), .B2(new_n665), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT28), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n619), .A2(new_n622), .A3(new_n623), .ZN(new_n670));
  INV_X1    g0470(.A(new_n631), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n630), .B1(new_n490), .B2(new_n602), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n634), .A2(new_n637), .A3(new_n620), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n647), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n635), .A2(new_n636), .A3(new_n571), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n620), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n636), .B1(new_n622), .B2(new_n635), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n670), .B1(new_n627), .B2(new_n628), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n660), .ZN(new_n682));
  MUX2_X1   g0482(.A(new_n675), .B(new_n682), .S(KEYINPUT29), .Z(new_n683));
  NOR2_X1   g0483(.A1(new_n543), .A2(new_n325), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n505), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n596), .A2(new_n597), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n685), .A2(new_n686), .A3(KEYINPUT30), .A4(new_n462), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n505), .A2(new_n684), .A3(new_n596), .A4(new_n597), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n689), .B2(new_n483), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n505), .A2(G179), .A3(new_n540), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n691), .A2(new_n483), .A3(new_n604), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n687), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n647), .ZN(new_n694));
  XNOR2_X1  g0494(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT31), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(new_n694), .ZN(new_n698));
  AOI21_X1  g0498(.A(KEYINPUT90), .B1(new_n607), .B2(new_n660), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n619), .A2(new_n623), .A3(new_n602), .A4(new_n571), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT90), .ZN(new_n701));
  NOR4_X1   g0501(.A1(new_n700), .A2(new_n494), .A3(new_n701), .A4(new_n647), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n698), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n683), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n669), .B1(new_n705), .B2(G1), .ZN(G364));
  NOR2_X1   g0506(.A1(new_n259), .A2(G20), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n207), .B1(new_n707), .B2(G45), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n664), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n655), .B2(G330), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(G330), .B2(new_n655), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n663), .A2(new_n407), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G355), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(G116), .B2(new_n211), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n663), .A2(new_n289), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n232), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n717), .B1(new_n443), .B2(new_n718), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n246), .A2(new_n443), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n715), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G13), .A2(G33), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n233), .B1(G20), .B2(new_n365), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n710), .B1(new_n721), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n325), .A2(G200), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n208), .A2(G190), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n293), .B1(new_n732), .B2(G311), .ZN(new_n733));
  INV_X1    g0533(.A(G322), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n208), .A2(new_n317), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n729), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n733), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n735), .A2(new_n325), .A3(G200), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n738), .A2(KEYINPUT94), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(KEYINPUT94), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n737), .B1(new_n742), .B2(G303), .ZN(new_n743));
  NAND3_X1  g0543(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G190), .ZN(new_n745));
  INV_X1    g0545(.A(G317), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n746), .A2(KEYINPUT33), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(KEYINPUT33), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n317), .A2(G179), .A3(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n208), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n744), .A2(new_n317), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n752), .A2(G294), .B1(G326), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n743), .A2(new_n749), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n730), .A2(new_n325), .A3(new_n506), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT95), .Z(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G329), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n730), .A2(new_n325), .A3(G200), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT92), .Z(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G283), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n758), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n751), .B(KEYINPUT93), .Z(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G97), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n760), .A2(G107), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n293), .B1(new_n738), .B2(new_n218), .ZN(new_n767));
  INV_X1    g0567(.A(new_n736), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n767), .B1(G58), .B2(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n745), .A2(G68), .B1(new_n753), .B2(G50), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n765), .A2(new_n766), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  OR3_X1    g0571(.A1(new_n756), .A2(KEYINPUT32), .A3(new_n266), .ZN(new_n772));
  OAI21_X1  g0572(.A(KEYINPUT32), .B1(new_n756), .B2(new_n266), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n732), .A2(KEYINPUT91), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n732), .A2(KEYINPUT91), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n772), .B(new_n773), .C1(new_n777), .C2(new_n202), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n755), .A2(new_n763), .B1(new_n771), .B2(new_n778), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n779), .A2(KEYINPUT96), .ZN(new_n780));
  INV_X1    g0580(.A(new_n725), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(new_n779), .B2(KEYINPUT96), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n728), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n724), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n783), .B1(new_n655), .B2(new_n784), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n712), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(G396));
  NAND2_X1  g0587(.A1(new_n421), .A2(new_n647), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n612), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n426), .A2(new_n428), .A3(new_n788), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n675), .B(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n710), .B1(new_n794), .B2(new_n704), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT99), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n794), .A2(new_n704), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n725), .A2(new_n722), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT97), .Z(new_n802));
  OAI21_X1  g0602(.A(new_n710), .B1(new_n802), .B2(G77), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n792), .A2(new_n723), .ZN(new_n804));
  INV_X1    g0604(.A(G294), .ZN(new_n805));
  INV_X1    g0605(.A(new_n753), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n407), .B1(new_n736), .B2(new_n805), .C1(new_n453), .C2(new_n806), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n777), .A2(new_n472), .B1(new_n741), .B2(new_n511), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n807), .B(new_n808), .C1(G283), .C2(new_n745), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n760), .A2(G87), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n757), .A2(G311), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n809), .A2(new_n765), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(KEYINPUT98), .B(G143), .Z(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n814), .A2(new_n768), .B1(G137), .B2(new_n753), .ZN(new_n815));
  INV_X1    g0615(.A(new_n745), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n815), .B1(new_n340), .B2(new_n816), .C1(new_n777), .C2(new_n266), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT34), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n289), .B1(new_n222), .B2(new_n751), .C1(new_n741), .C2(new_n347), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G132), .B2(new_n757), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n817), .A2(new_n818), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n760), .A2(G68), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n812), .B1(new_n819), .B2(new_n824), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n803), .B(new_n804), .C1(new_n725), .C2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n800), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G384));
  OR2_X1    g0628(.A1(new_n515), .A2(KEYINPUT35), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n515), .A2(KEYINPUT35), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n233), .A2(new_n208), .A3(new_n472), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT36), .Z(new_n833));
  OR4_X1    g0633(.A1(new_n202), .A2(new_n262), .A3(new_n263), .A4(new_n232), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n347), .A2(G68), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n207), .B(G13), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n381), .A2(new_n647), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n400), .A2(new_n403), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n404), .A2(new_n381), .A3(new_n647), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n793), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(KEYINPUT102), .B1(new_n694), .B2(new_n697), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT102), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n693), .A2(new_n843), .A3(KEYINPUT31), .A4(new_n647), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n842), .A2(new_n844), .B1(new_n694), .B2(new_n695), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n699), .B2(new_n702), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n292), .A2(new_n345), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n269), .B1(new_n287), .B2(new_n291), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n849), .B1(KEYINPUT16), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n851), .A2(new_n261), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n852), .A2(new_n645), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n339), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n319), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n856), .A2(new_n327), .ZN(new_n857));
  INV_X1    g0657(.A(new_n645), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n335), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n326), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n319), .B1(new_n852), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(KEYINPUT37), .B1(new_n862), .B2(new_n853), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT38), .B1(new_n854), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT17), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n319), .B(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT77), .B1(new_n331), .B2(new_n332), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n336), .A2(new_n334), .A3(new_n337), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n853), .ZN(new_n871));
  OAI211_X1 g0671(.A(KEYINPUT38), .B(new_n864), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n848), .B1(new_n865), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT40), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n611), .B1(new_n320), .B2(KEYINPUT100), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT100), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n867), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n859), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n319), .A2(new_n610), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n855), .B1(new_n859), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n859), .B2(new_n857), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n876), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n872), .A2(new_n885), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n841), .A2(new_n846), .A3(KEYINPUT40), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n874), .A2(new_n875), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n888), .B(KEYINPUT103), .Z(new_n889));
  AND2_X1   g0689(.A1(new_n433), .A2(new_n846), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n891), .A2(G330), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n864), .B1(new_n870), .B2(new_n871), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n876), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n872), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n404), .B(new_n838), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n660), .B(new_n792), .C1(new_n632), .C2(new_n638), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n426), .A2(new_n647), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n897), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n896), .A2(new_n901), .B1(new_n611), .B2(new_n645), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n886), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n895), .A2(KEYINPUT39), .A3(new_n872), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n400), .A2(new_n647), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n902), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT101), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n902), .B(KEYINPUT101), .C1(new_n906), .C2(new_n908), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n616), .B1(new_n683), .B2(new_n433), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n913), .B(new_n914), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n893), .A2(new_n915), .B1(new_n207), .B2(new_n707), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n893), .A2(new_n915), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n837), .B1(new_n916), .B2(new_n917), .ZN(G367));
  NAND2_X1  g0718(.A1(new_n523), .A2(new_n647), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n619), .A2(KEYINPUT105), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n530), .B2(new_n660), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT105), .B1(new_n619), .B2(new_n919), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n659), .A2(new_n641), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT42), .Z(new_n926));
  XNOR2_X1  g0726(.A(new_n923), .B(KEYINPUT106), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n530), .B1(new_n927), .B2(new_n602), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n926), .B1(new_n660), .B2(new_n928), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n570), .A2(new_n660), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n622), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n620), .B2(new_n930), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(KEYINPUT104), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n932), .A2(KEYINPUT104), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT43), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n929), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n929), .B2(new_n937), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n927), .A2(new_n658), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n939), .B(new_n940), .Z(new_n941));
  XOR2_X1   g0741(.A(new_n664), .B(KEYINPUT41), .Z(new_n942));
  NAND2_X1  g0742(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n943));
  INV_X1    g0743(.A(new_n923), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n943), .B1(new_n944), .B2(new_n661), .ZN(new_n945));
  NOR2_X1   g0745(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT109), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n945), .B(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n944), .A2(new_n661), .ZN(new_n949));
  XOR2_X1   g0749(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(new_n658), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n924), .B1(new_n651), .B2(new_n659), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(new_n656), .Z(new_n955));
  NAND3_X1  g0755(.A1(new_n953), .A2(new_n705), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n942), .B1(new_n956), .B2(new_n705), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n941), .B1(new_n957), .B2(new_n709), .ZN(new_n958));
  INV_X1    g0758(.A(new_n710), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n726), .B1(new_n211), .B2(new_n415), .C1(new_n717), .C2(new_n242), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT110), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n961), .B2(new_n960), .ZN(new_n963));
  INV_X1    g0763(.A(new_n777), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(G50), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n806), .A2(new_n813), .B1(new_n816), .B2(new_n266), .ZN(new_n966));
  INV_X1    g0766(.A(G137), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n756), .A2(new_n967), .B1(new_n759), .B2(new_n202), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n764), .A2(G68), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n293), .B1(new_n738), .B2(new_n222), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(G150), .B2(new_n768), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n965), .A2(new_n969), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n964), .A2(G283), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n289), .B1(G303), .B2(new_n768), .ZN(new_n975));
  INV_X1    g0775(.A(new_n738), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT46), .B1(new_n976), .B2(G116), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(G311), .B2(new_n753), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n742), .A2(KEYINPUT46), .A3(G116), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n974), .A2(new_n975), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n756), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n981), .A2(G317), .B1(G294), .B2(new_n745), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n982), .B1(new_n224), .B2(new_n759), .C1(new_n511), .C2(new_n751), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n973), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT47), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n963), .B1(new_n985), .B2(new_n725), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n932), .B2(new_n784), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n958), .A2(new_n987), .ZN(G387));
  NAND2_X1  g0788(.A1(new_n955), .A2(new_n709), .ZN(new_n989));
  INV_X1    g0789(.A(new_n666), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n713), .A2(new_n990), .B1(new_n511), .B2(new_n663), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n239), .A2(new_n443), .ZN(new_n992));
  INV_X1    g0792(.A(new_n251), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n347), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT50), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n666), .B(new_n443), .C1(new_n216), .C2(new_n202), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n716), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n991), .B1(new_n992), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n959), .B1(new_n998), .B2(new_n726), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n768), .A2(G317), .B1(G311), .B2(new_n745), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n734), .B2(new_n806), .C1(new_n777), .C2(new_n453), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT48), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G283), .A2(new_n752), .B1(new_n976), .B2(G294), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1007), .A2(KEYINPUT49), .ZN(new_n1008));
  INV_X1    g0808(.A(G326), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n451), .B1(new_n472), .B2(new_n759), .C1(new_n1009), .C2(new_n756), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n1007), .B2(KEYINPUT49), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n976), .A2(G77), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n347), .B2(new_n736), .C1(new_n216), .C2(new_n731), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n253), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1014), .A2(new_n816), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n756), .A2(new_n340), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n289), .B1(new_n806), .B2(new_n266), .ZN(new_n1017));
  NOR4_X1   g0817(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n764), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1019), .A2(new_n415), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G97), .B2(new_n760), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1008), .A2(new_n1011), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n999), .B1(new_n651), .B2(new_n784), .C1(new_n781), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n705), .A2(new_n955), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n664), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n705), .A2(new_n955), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n989), .B(new_n1023), .C1(new_n1025), .C2(new_n1026), .ZN(G393));
  INV_X1    g0827(.A(new_n953), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n1024), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n956), .A2(new_n664), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n953), .A2(new_n709), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n927), .A2(new_n724), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n768), .A2(G311), .B1(G317), .B2(new_n753), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT52), .Z(new_n1034));
  OAI22_X1  g0834(.A1(new_n751), .A2(new_n472), .B1(new_n756), .B2(new_n734), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G303), .B2(new_n745), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n407), .B1(new_n731), .B2(new_n805), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G283), .B2(new_n976), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1034), .A2(new_n766), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n964), .A2(new_n993), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n756), .A2(new_n813), .B1(new_n816), .B2(new_n347), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n451), .B(new_n1041), .C1(G68), .C2(new_n976), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n764), .A2(G77), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1040), .A2(new_n1042), .A3(new_n810), .A4(new_n1043), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n768), .A2(G159), .B1(G150), .B2(new_n753), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT51), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1039), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n725), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n726), .B1(new_n224), .B2(new_n211), .C1(new_n717), .C2(new_n249), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1032), .A2(new_n710), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1030), .A2(new_n1031), .A3(new_n1050), .ZN(G390));
  OAI21_X1  g0851(.A(KEYINPUT111), .B1(new_n901), .B2(new_n907), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT111), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n899), .B1(new_n675), .B2(new_n792), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1053), .B(new_n908), .C1(new_n1054), .C2(new_n897), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n906), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n900), .B1(new_n682), .B2(new_n793), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n840), .A2(new_n839), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n907), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n886), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n792), .A2(G330), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n703), .A2(new_n1058), .A3(new_n1061), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n846), .A2(new_n1061), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1062), .B1(new_n1064), .B2(KEYINPUT112), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  AND3_X1   g0866(.A1(new_n1056), .A2(new_n1060), .A3(new_n1066), .ZN(new_n1067));
  AND3_X1   g0867(.A1(new_n846), .A2(new_n1058), .A3(new_n1061), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1056), .A2(new_n1060), .B1(KEYINPUT112), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1054), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1058), .B1(new_n703), .B2(new_n1061), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1071), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(KEYINPUT114), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT114), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1075), .B(new_n1071), .C1(new_n1068), .C2(new_n1072), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1062), .A2(new_n1057), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n430), .A2(new_n432), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1081), .A2(new_n846), .A3(G330), .A4(new_n870), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT113), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1082), .B(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n914), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1080), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n665), .B1(new_n1070), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1085), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n723), .B1(new_n904), .B2(new_n905), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n757), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1043), .B(new_n823), .C1(new_n805), .C2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n816), .A2(new_n511), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n407), .B1(new_n736), .B2(new_n472), .C1(new_n762), .C2(new_n806), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n777), .A2(new_n224), .B1(new_n741), .B2(new_n218), .ZN(new_n1097));
  NOR4_X1   g0897(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(G128), .ZN(new_n1099));
  INV_X1    g0899(.A(G132), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n806), .A2(new_n1099), .B1(new_n736), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n745), .A2(G137), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(KEYINPUT54), .B(G143), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1102), .B1(new_n777), .B2(new_n1103), .C1(new_n1019), .C2(new_n266), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT115), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT53), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n738), .B2(new_n340), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n976), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1101), .B(new_n1105), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n293), .B1(new_n759), .B2(new_n347), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n757), .B2(G125), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT116), .Z(new_n1112));
  AOI21_X1  g0912(.A(new_n1098), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n710), .B1(new_n253), .B2(new_n802), .C1(new_n1113), .C2(new_n781), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1070), .A2(new_n708), .B1(new_n1092), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1091), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(G378));
  NAND2_X1  g0917(.A1(new_n1090), .A2(new_n1086), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n887), .A2(new_n886), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n847), .B1(new_n895), .B2(new_n872), .ZN(new_n1120));
  OAI211_X1 g0920(.A(G330), .B(new_n1119), .C1(new_n1120), .C2(KEYINPUT40), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n350), .A2(new_n645), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n369), .B(new_n1122), .Z(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1123), .B(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT119), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1121), .A2(KEYINPUT119), .A3(new_n1125), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n911), .A2(new_n912), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1125), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n888), .A2(KEYINPUT120), .A3(G330), .A4(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT120), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1130), .A2(new_n1131), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1131), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1138));
  OAI211_X1 g0938(.A(KEYINPUT57), .B(new_n1118), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(KEYINPUT121), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1118), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT57), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1121), .A2(KEYINPUT119), .A3(new_n1125), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT119), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n913), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1130), .A2(new_n1131), .A3(new_n1136), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT121), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1150), .A2(new_n1151), .A3(KEYINPUT57), .A4(new_n1118), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1140), .A2(new_n1143), .A3(new_n1152), .A4(new_n664), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1125), .A2(new_n722), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n710), .B1(new_n802), .B2(G50), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(G33), .A2(G41), .ZN(new_n1156));
  AOI211_X1 g0956(.A(G50), .B(new_n1156), .C1(new_n451), .C2(new_n435), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1012), .B1(new_n222), .B2(new_n759), .C1(new_n511), .C2(new_n736), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n806), .A2(new_n472), .ZN(new_n1159));
  NOR4_X1   g0959(.A1(new_n1158), .A2(G41), .A3(new_n289), .A4(new_n1159), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n732), .A2(new_n547), .B1(G97), .B2(new_n745), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT117), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n757), .A2(G283), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1160), .A2(new_n970), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT58), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1157), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n738), .A2(new_n1103), .B1(new_n736), .B2(new_n1099), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G137), .B2(new_n732), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n745), .A2(G132), .B1(new_n753), .B2(G125), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(new_n1019), .C2(new_n340), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT118), .Z(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(KEYINPUT59), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n981), .A2(G124), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n759), .A2(new_n266), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n1156), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1171), .A2(KEYINPUT59), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1166), .B1(new_n1165), .B2(new_n1164), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1155), .B1(new_n1177), .B2(new_n725), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1150), .A2(new_n709), .B1(new_n1154), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1153), .A2(new_n1179), .ZN(G375));
  NOR2_X1   g0980(.A1(new_n1080), .A2(new_n1086), .ZN(new_n1181));
  OR3_X1    g0981(.A1(new_n1181), .A2(new_n1089), .A3(new_n942), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n897), .A2(new_n722), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n710), .B1(new_n802), .B2(G68), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n1019), .A2(new_n415), .B1(new_n761), .B2(new_n202), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n407), .B1(new_n736), .B2(new_n762), .C1(new_n805), .C2(new_n806), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G116), .B2(new_n745), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n224), .B2(new_n741), .C1(new_n511), .C2(new_n777), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1185), .B(new_n1188), .C1(G303), .C2(new_n757), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1189), .A2(KEYINPUT122), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(KEYINPUT122), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n764), .A2(G50), .B1(new_n757), .B2(G128), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n289), .B1(new_n967), .B2(new_n736), .C1(new_n340), .C2(new_n731), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n742), .B2(G159), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n816), .A2(new_n1103), .B1(new_n759), .B2(new_n222), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G132), .B2(new_n753), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1192), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1190), .A2(new_n1191), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1184), .B1(new_n1198), .B2(new_n725), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1080), .A2(new_n709), .B1(new_n1183), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1182), .A2(new_n1200), .ZN(G381));
  INV_X1    g1001(.A(G390), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n958), .A2(new_n1202), .A3(new_n987), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1204), .A2(new_n1200), .A3(new_n1182), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT123), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1153), .A2(new_n1116), .A3(new_n1179), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT124), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1212), .A2(new_n1213), .ZN(G407));
  INV_X1    g1014(.A(G213), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n1209), .B2(new_n646), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1212), .B2(new_n1213), .ZN(G409));
  INV_X1    g1017(.A(KEYINPUT61), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1215), .A2(G343), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1153), .A2(G378), .A3(new_n1179), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1179), .B1(new_n942), .B2(new_n1141), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1116), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1219), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1219), .A2(G2897), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1087), .A2(KEYINPUT60), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n665), .B1(new_n1226), .B2(new_n1181), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1181), .B2(new_n1226), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1228), .A2(G384), .A3(new_n1200), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(G384), .B1(new_n1228), .B2(new_n1200), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1225), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1228), .A2(new_n1200), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n827), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(new_n1229), .A3(new_n1224), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1218), .B1(new_n1223), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT127), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  OAI211_X1 g1039(.A(KEYINPUT127), .B(new_n1218), .C1(new_n1223), .C2(new_n1236), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1223), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT62), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT62), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1223), .A2(new_n1244), .A3(new_n1241), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1239), .A2(new_n1240), .A3(new_n1243), .A4(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(G387), .A2(G390), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1203), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(G393), .B(new_n786), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT126), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1247), .B(new_n1203), .C1(KEYINPUT126), .C2(new_n1249), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1246), .A2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1253), .B(new_n1218), .C1(new_n1223), .C2(new_n1236), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1242), .A2(KEYINPUT125), .A3(KEYINPUT63), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT63), .B1(new_n1242), .B2(KEYINPUT125), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1257), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1255), .A2(new_n1260), .ZN(G405));
  XNOR2_X1  g1061(.A(G375), .B(G378), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1241), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1264), .A2(new_n1254), .A3(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1254), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(G402));
endmodule


