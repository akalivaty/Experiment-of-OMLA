//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1251, new_n1252, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  OAI21_X1  g0006(.A(G50), .B1(G58), .B2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G50), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G116), .ZN(new_n221));
  INV_X1    g0021(.A(G270), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n217), .B1(new_n223), .B2(KEYINPUT64), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT65), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n224), .B(new_n226), .C1(KEYINPUT64), .C2(new_n223), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(new_n203), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n206), .B(new_n212), .C1(new_n228), .C2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(new_n214), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n247), .B1(G41), .B2(G45), .ZN(new_n248));
  INV_X1    g0048(.A(G274), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n209), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n248), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n250), .B1(new_n255), .B2(G226), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT67), .ZN(new_n259));
  NOR3_X1   g0059(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  AOI21_X1  g0064(.A(KEYINPUT67), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G222), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G77), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n268), .B1(new_n269), .B2(new_n266), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n259), .B1(new_n257), .B2(new_n258), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n263), .A2(KEYINPUT67), .A3(new_n264), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(new_n272), .A3(G1698), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT68), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n270), .B1(G223), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n256), .B1(new_n275), .B2(new_n253), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G200), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT9), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G50), .A2(G58), .ZN(new_n280));
  INV_X1    g0080(.A(G68), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n210), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n282), .B(KEYINPUT69), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n210), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(G150), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n284), .A2(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n209), .B1(new_n203), .B2(new_n262), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G13), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n294), .A2(new_n210), .A3(G1), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(new_n291), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n247), .A2(G20), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G50), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n294), .A2(G1), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G20), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n297), .A2(new_n299), .B1(G50), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n279), .B1(new_n293), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n302), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n304), .B(KEYINPUT9), .C1(new_n292), .C2(new_n290), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G190), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n276), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT10), .B1(new_n278), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n276), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G190), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n311), .A2(new_n312), .A3(new_n277), .A4(new_n306), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n250), .B1(new_n255), .B2(G244), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n271), .A2(new_n272), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G107), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n266), .A2(G232), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n318), .B1(new_n319), .B2(G1698), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(G238), .B2(new_n274), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n315), .B(new_n316), .C1(new_n321), .C2(new_n253), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n297), .A2(KEYINPUT71), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT71), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n296), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(G77), .A3(new_n298), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n295), .A2(new_n269), .ZN(new_n328));
  XOR2_X1   g0128(.A(KEYINPUT15), .B(G87), .Z(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n330), .A2(new_n285), .B1(new_n210), .B2(new_n269), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n284), .A2(new_n288), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n291), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n327), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n316), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n274), .A2(G238), .ZN(new_n336));
  INV_X1    g0136(.A(new_n320), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n335), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n322), .B(new_n334), .C1(new_n340), .C2(G169), .ZN(new_n341));
  OAI211_X1 g0141(.A(G190), .B(new_n316), .C1(new_n321), .C2(new_n253), .ZN(new_n342));
  INV_X1    g0142(.A(new_n334), .ZN(new_n343));
  INV_X1    g0143(.A(G200), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n342), .B(new_n343), .C1(new_n340), .C2(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT72), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n284), .B1(new_n247), .B2(G20), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(new_n296), .B1(new_n295), .B2(new_n284), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT7), .B1(new_n317), .B2(new_n210), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n264), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT76), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n257), .A2(new_n258), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT76), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n354), .A2(new_n355), .A3(KEYINPUT7), .A4(new_n210), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(G68), .B1(new_n351), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n213), .A2(new_n281), .ZN(new_n359));
  NOR2_X1   g0159(.A1(G58), .A2(G68), .ZN(new_n360));
  OAI21_X1  g0160(.A(G20), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n287), .A2(G159), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT16), .B1(new_n358), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT7), .B1(new_n354), .B2(new_n210), .ZN(new_n366));
  INV_X1    g0166(.A(new_n352), .ZN(new_n367));
  OAI21_X1  g0167(.A(G68), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(KEYINPUT16), .A3(new_n364), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n291), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n350), .B1(new_n365), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT18), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n220), .A2(G1698), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n373), .B1(G223), .B2(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G87), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n253), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n250), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n254), .B2(new_n214), .ZN(new_n378));
  OAI21_X1  g0178(.A(G169), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n376), .A2(new_n378), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(new_n380), .B2(new_n315), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n371), .A2(new_n372), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n372), .B1(new_n371), .B2(new_n381), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT16), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n210), .B1(new_n260), .B2(new_n265), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT7), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g0188(.A(new_n352), .B(new_n355), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n281), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n385), .B1(new_n390), .B2(new_n363), .ZN(new_n391));
  INV_X1    g0191(.A(new_n370), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n344), .B1(new_n376), .B2(new_n378), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n380), .B2(G190), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n393), .A2(KEYINPUT17), .A3(new_n350), .A4(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n395), .B(new_n350), .C1(new_n365), .C2(new_n370), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n314), .A2(new_n348), .A3(new_n384), .A4(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G238), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n377), .B1(new_n254), .B2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n271), .A2(new_n272), .A3(G232), .A4(G1698), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n271), .A2(new_n272), .A3(G226), .A4(new_n267), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G97), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n403), .B1(new_n407), .B2(new_n339), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT13), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI211_X1 g0210(.A(KEYINPUT13), .B(new_n403), .C1(new_n407), .C2(new_n339), .ZN(new_n411));
  OAI21_X1  g0211(.A(G169), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT14), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n407), .A2(new_n339), .ZN(new_n415));
  INV_X1    g0215(.A(new_n403), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT13), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n408), .A2(new_n409), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(KEYINPUT14), .A3(G169), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT73), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n417), .A2(new_n422), .A3(KEYINPUT13), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT73), .B1(new_n408), .B2(new_n409), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n423), .A2(new_n424), .A3(new_n419), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n414), .A2(new_n421), .B1(new_n425), .B2(G179), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT75), .ZN(new_n427));
  AOI211_X1 g0227(.A(G68), .B(new_n301), .C1(new_n427), .C2(KEYINPUT12), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(KEYINPUT12), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n428), .B(new_n429), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n288), .A2(new_n219), .B1(new_n210), .B2(G68), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n285), .A2(new_n269), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n291), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  XOR2_X1   g0233(.A(KEYINPUT74), .B(KEYINPUT11), .Z(new_n434));
  XNOR2_X1  g0234(.A(new_n433), .B(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n326), .A2(G68), .A3(new_n298), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n426), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n420), .A2(G200), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n423), .A2(new_n424), .A3(G190), .A4(new_n419), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(new_n438), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n310), .A2(new_n315), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n293), .A2(new_n302), .ZN(new_n446));
  INV_X1    g0246(.A(G169), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n446), .B1(new_n276), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(KEYINPUT70), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT70), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n451), .B1(new_n445), .B2(new_n448), .ZN(new_n452));
  OAI22_X1  g0252(.A1(new_n450), .A2(new_n452), .B1(new_n346), .B2(new_n347), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n401), .A2(new_n444), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n262), .A2(G1), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT78), .ZN(new_n457));
  AND4_X1   g0257(.A1(G116), .A2(new_n323), .A3(new_n325), .A4(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n300), .A2(G20), .A3(new_n221), .ZN(new_n459));
  AOI21_X1  g0259(.A(G20), .B1(G33), .B2(G283), .ZN(new_n460));
  INV_X1    g0260(.A(G97), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n460), .B1(G33), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n462), .B(new_n291), .C1(new_n210), .C2(G116), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT20), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n463), .A2(new_n464), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n459), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n458), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g0269(.A(KEYINPUT5), .B(G41), .ZN(new_n470));
  INV_X1    g0270(.A(G45), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G1), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n253), .A2(new_n470), .A3(G274), .A4(new_n472), .ZN(new_n473));
  AND2_X1   g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  NOR2_X1   g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n253), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n473), .B1(new_n477), .B2(new_n222), .ZN(new_n478));
  OAI21_X1  g0278(.A(G303), .B1(new_n260), .B2(new_n265), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n263), .A2(new_n264), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n216), .A2(new_n267), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(G257), .B(new_n267), .C1(new_n257), .C2(new_n258), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT81), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n480), .A2(KEYINPUT81), .A3(G257), .A4(new_n267), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n479), .A2(new_n482), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n478), .B1(new_n487), .B2(new_n339), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(new_n447), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT21), .B1(new_n469), .B2(new_n489), .ZN(new_n490));
  AOI211_X1 g0290(.A(new_n315), .B(new_n478), .C1(new_n487), .C2(new_n339), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(new_n489), .B2(KEYINPUT21), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT82), .B1(new_n492), .B2(new_n468), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n487), .A2(new_n339), .ZN(new_n494));
  INV_X1    g0294(.A(new_n478), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(KEYINPUT21), .A3(G169), .ZN(new_n497));
  INV_X1    g0297(.A(new_n491), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT82), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(new_n500), .A3(new_n469), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n490), .B1(new_n493), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G87), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n503), .A2(KEYINPUT22), .A3(G20), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n271), .A2(new_n272), .A3(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n210), .B(G87), .C1(new_n257), .C2(new_n258), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n506), .A2(KEYINPUT83), .A3(KEYINPUT22), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT83), .B1(new_n506), .B2(KEYINPUT22), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT24), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT23), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n210), .B2(G107), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n215), .A2(KEYINPUT23), .A3(G20), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G116), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n512), .A2(new_n513), .B1(new_n515), .B2(new_n210), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n509), .A2(new_n510), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n510), .B1(new_n509), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n291), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n457), .A2(new_n296), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n520), .A2(new_n215), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n295), .A2(KEYINPUT25), .A3(new_n215), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT84), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT25), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n301), .B2(G107), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g0326(.A1(new_n523), .A2(new_n525), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n521), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n519), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(G250), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n267), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(G257), .B2(new_n267), .ZN(new_n532));
  INV_X1    g0332(.A(G294), .ZN(new_n533));
  OAI22_X1  g0333(.A1(new_n532), .A2(new_n354), .B1(new_n262), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n470), .A2(new_n472), .B1(new_n251), .B2(new_n252), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n534), .A2(new_n339), .B1(new_n535), .B2(G264), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n473), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(G179), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n447), .B2(new_n537), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n529), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n502), .A2(new_n540), .ZN(new_n541));
  MUX2_X1   g0341(.A(new_n301), .B(new_n520), .S(G97), .Z(new_n542));
  NAND2_X1  g0342(.A1(new_n287), .A2(G77), .ZN(new_n543));
  XNOR2_X1  g0343(.A(new_n543), .B(KEYINPUT77), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT6), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n545), .A2(new_n461), .A3(G107), .ZN(new_n546));
  XNOR2_X1  g0346(.A(G97), .B(G107), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n544), .B1(new_n210), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(G20), .B1(new_n271), .B2(new_n272), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n353), .B(new_n356), .C1(new_n550), .C2(KEYINPUT7), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n549), .B1(new_n551), .B2(G107), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n542), .B1(new_n552), .B2(new_n292), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n476), .A2(G257), .A3(new_n253), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n473), .ZN(new_n555));
  OAI211_X1 g0355(.A(G244), .B(new_n267), .C1(new_n257), .C2(new_n258), .ZN(new_n556));
  XNOR2_X1  g0356(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n556), .A2(new_n557), .B1(G33), .B2(G283), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n271), .A2(new_n272), .A3(G250), .A4(G1698), .ZN(new_n559));
  AND2_X1   g0359(.A1(KEYINPUT4), .A2(G244), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n271), .A2(new_n272), .A3(new_n267), .A4(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n555), .B1(new_n562), .B2(new_n339), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n315), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n339), .ZN(new_n565));
  INV_X1    g0365(.A(new_n555), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n447), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n553), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n215), .B1(new_n388), .B2(new_n389), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n291), .B1(new_n570), .B2(new_n549), .ZN(new_n571));
  AOI21_X1  g0371(.A(G200), .B1(new_n565), .B2(new_n566), .ZN(new_n572));
  AOI211_X1 g0372(.A(G190), .B(new_n555), .C1(new_n562), .C2(new_n339), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n571), .B(new_n542), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n488), .A2(G190), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n485), .A2(new_n486), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n317), .A2(G303), .B1(new_n480), .B2(new_n481), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n253), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(G200), .B1(new_n578), .B2(new_n478), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n468), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n569), .A2(new_n574), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n537), .A2(new_n344), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(G190), .B2(new_n537), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n519), .A2(new_n528), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n247), .A2(G45), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G250), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n339), .A2(new_n586), .B1(new_n249), .B2(new_n585), .ZN(new_n587));
  OAI211_X1 g0387(.A(G244), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n588));
  OAI211_X1 g0388(.A(G238), .B(new_n267), .C1(new_n257), .C2(new_n258), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n589), .A3(new_n514), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n307), .B(new_n587), .C1(new_n339), .C2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n329), .A2(new_n301), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT19), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n210), .B1(new_n406), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n503), .A2(new_n461), .A3(new_n215), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n210), .B(G68), .C1(new_n257), .C2(new_n258), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n593), .B1(new_n285), .B2(new_n461), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n592), .B1(new_n599), .B2(new_n291), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n457), .A2(G87), .A3(new_n296), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n587), .B1(new_n590), .B2(new_n339), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n600), .B(new_n601), .C1(new_n602), .C2(new_n344), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT80), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n591), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n590), .A2(new_n339), .ZN(new_n606));
  INV_X1    g0406(.A(new_n587), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(G200), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n609), .A2(KEYINPUT80), .A3(new_n600), .A4(new_n601), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n447), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n457), .A2(new_n296), .A3(new_n329), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n600), .A2(new_n612), .B1(new_n602), .B2(new_n315), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n605), .A2(new_n610), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n584), .A2(new_n614), .ZN(new_n615));
  NOR4_X1   g0415(.A1(new_n455), .A2(new_n541), .A3(new_n581), .A4(new_n615), .ZN(G372));
  NOR2_X1   g0416(.A1(new_n450), .A2(new_n452), .ZN(new_n617));
  INV_X1    g0417(.A(new_n341), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n618), .A2(new_n443), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n400), .B1(new_n619), .B2(new_n439), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT86), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n382), .B2(new_n383), .ZN(new_n622));
  INV_X1    g0422(.A(new_n350), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(new_n391), .B2(new_n392), .ZN(new_n624));
  INV_X1    g0424(.A(new_n381), .ZN(new_n625));
  OAI21_X1  g0425(.A(KEYINPUT18), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n371), .A2(new_n372), .A3(new_n381), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(KEYINPUT86), .A3(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n620), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n617), .B1(new_n630), .B2(new_n314), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n569), .A2(new_n574), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n609), .A2(KEYINPUT85), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n600), .A2(new_n601), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n591), .A2(new_n634), .ZN(new_n635));
  OR3_X1    g0435(.A1(new_n602), .A2(KEYINPUT85), .A3(new_n344), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n613), .A2(new_n611), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n632), .A2(new_n584), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n490), .B1(new_n469), .B2(new_n499), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n641), .B1(new_n540), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n639), .A2(new_n569), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n605), .A2(new_n610), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n638), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n648), .A2(new_n569), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n646), .B(new_n638), .C1(new_n649), .C2(new_n645), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n631), .B1(new_n455), .B2(new_n651), .ZN(G369));
  INV_X1    g0452(.A(G330), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n300), .A2(new_n210), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  INV_X1    g0456(.A(G213), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n468), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT87), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n502), .A2(new_n580), .A3(new_n661), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n642), .A2(new_n661), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n653), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n659), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n540), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n529), .A2(new_n666), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n584), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n669), .B2(new_n540), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n665), .A2(KEYINPUT88), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT88), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n664), .B2(new_n670), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n502), .A2(new_n666), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n667), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n675), .A2(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n204), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n595), .A2(G116), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G1), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n207), .B2(new_n683), .ZN(new_n686));
  XOR2_X1   g0486(.A(new_n686), .B(KEYINPUT28), .Z(new_n687));
  INV_X1    g0487(.A(new_n641), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n541), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n638), .B1(new_n644), .B2(new_n645), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n690), .B1(new_n645), .B2(new_n649), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n666), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT29), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n659), .B1(new_n643), .B2(new_n650), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT29), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n615), .A2(new_n581), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n502), .A2(new_n698), .A3(new_n540), .A4(new_n659), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n536), .A2(new_n602), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n488), .A2(new_n700), .A3(G179), .A4(new_n563), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n491), .A2(KEYINPUT30), .A3(new_n563), .A4(new_n700), .ZN(new_n704));
  AOI21_X1  g0504(.A(G179), .B1(new_n536), .B2(new_n473), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n496), .A2(new_n567), .A3(new_n608), .A4(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n666), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT31), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT31), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n707), .A2(new_n710), .A3(new_n666), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n699), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n697), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n687), .B1(new_n715), .B2(new_n247), .ZN(new_n716));
  XOR2_X1   g0516(.A(new_n716), .B(KEYINPUT89), .Z(G364));
  NOR2_X1   g0517(.A1(new_n294), .A2(G20), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n247), .B1(new_n718), .B2(G45), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n682), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n662), .A2(new_n663), .A3(new_n653), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n665), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n662), .A2(new_n663), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n317), .A2(new_n681), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G355), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(G116), .B2(new_n204), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n242), .A2(G45), .ZN(new_n732));
  AOI211_X1 g0532(.A(new_n480), .B(new_n681), .C1(new_n471), .C2(new_n208), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n209), .B1(G20), .B2(new_n447), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n727), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n721), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n735), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n210), .A2(new_n307), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n344), .A2(G179), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G303), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n210), .A2(G190), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n741), .ZN(new_n745));
  INV_X1    g0545(.A(G283), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n742), .A2(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G179), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G190), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n266), .B(new_n747), .C1(G294), .C2(new_n750), .ZN(new_n751));
  XOR2_X1   g0551(.A(KEYINPUT33), .B(G317), .Z(new_n752));
  NOR2_X1   g0552(.A1(new_n315), .A2(new_n344), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n744), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n315), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n740), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G322), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n752), .A2(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT90), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n755), .A2(new_n744), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  INV_X1    g0562(.A(G326), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n740), .A2(new_n753), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n761), .A2(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n744), .A2(new_n748), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n765), .B1(G329), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n751), .A2(new_n759), .A3(new_n768), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n761), .A2(new_n269), .B1(new_n219), .B2(new_n764), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n317), .ZN(new_n771));
  INV_X1    g0571(.A(G159), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n766), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT32), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n750), .A2(G97), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n213), .A2(new_n756), .B1(new_n754), .B2(new_n281), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n742), .A2(new_n503), .B1(new_n745), .B2(new_n215), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n771), .A2(new_n774), .A3(new_n775), .A4(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n739), .B1(new_n769), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n738), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n728), .A2(new_n781), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n724), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(G396));
  NOR2_X1   g0584(.A1(new_n735), .A2(new_n725), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT91), .Z(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n722), .B1(new_n787), .B2(new_n269), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n764), .A2(new_n743), .B1(new_n756), .B2(new_n533), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n761), .A2(new_n221), .B1(new_n215), .B2(new_n742), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT92), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n754), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n753), .A2(new_n744), .A3(KEYINPUT92), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n789), .B(new_n790), .C1(G283), .C2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n745), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G87), .A2(new_n796), .B1(new_n767), .B2(G311), .ZN(new_n797));
  AND4_X1   g0597(.A1(new_n317), .A2(new_n795), .A3(new_n775), .A4(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G137), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n764), .A2(new_n799), .B1(new_n754), .B2(new_n286), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT93), .ZN(new_n801));
  INV_X1    g0601(.A(G143), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n801), .B1(new_n802), .B2(new_n756), .C1(new_n772), .C2(new_n761), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT34), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n480), .B1(new_n742), .B2(new_n219), .ZN(new_n805));
  INV_X1    g0605(.A(G132), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n745), .A2(new_n281), .B1(new_n766), .B2(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n805), .B(new_n807), .C1(G58), .C2(new_n750), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n798), .B1(new_n804), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n334), .A2(new_n666), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n341), .A2(new_n345), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(KEYINPUT94), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n618), .A2(new_n666), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT94), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n341), .A2(new_n345), .A3(new_n814), .A4(new_n810), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n788), .B1(new_n739), .B2(new_n809), .C1(new_n816), .C2(new_n726), .ZN(new_n817));
  INV_X1    g0617(.A(new_n714), .ZN(new_n818));
  INV_X1    g0618(.A(new_n816), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n694), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n812), .A2(new_n815), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n821), .B(new_n659), .C1(new_n643), .C2(new_n650), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n818), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n823), .A2(KEYINPUT95), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(KEYINPUT95), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT96), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n818), .B1(new_n820), .B2(new_n822), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n824), .B(new_n825), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n826), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n722), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n817), .B1(new_n828), .B2(new_n830), .ZN(G384));
  INV_X1    g0631(.A(new_n548), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n832), .A2(KEYINPUT35), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(KEYINPUT35), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n833), .A2(G116), .A3(new_n211), .A4(new_n834), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT36), .Z(new_n836));
  OAI211_X1 g0636(.A(new_n208), .B(G77), .C1(new_n213), .C2(new_n281), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n219), .A2(G68), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n247), .B(G13), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n440), .A2(new_n666), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT98), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT97), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n626), .A2(new_n627), .A3(new_n399), .A4(new_n396), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n387), .B1(new_n480), .B2(G20), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n281), .B1(new_n845), .B2(new_n352), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n385), .B1(new_n846), .B2(new_n363), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n847), .A2(new_n291), .A3(new_n369), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n848), .A2(new_n623), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n658), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n371), .A2(new_n381), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n371), .A2(new_n658), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT37), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n852), .A2(new_n853), .A3(new_n854), .A4(new_n397), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n848), .A2(new_n623), .B1(new_n381), .B2(new_n658), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n397), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT37), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n844), .A2(new_n851), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n843), .B1(new_n859), .B2(KEYINPUT38), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n850), .B1(new_n384), .B2(new_n400), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n855), .A2(new_n858), .ZN(new_n863));
  OAI211_X1 g0663(.A(KEYINPUT97), .B(new_n861), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n844), .A2(new_n851), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n855), .A2(new_n858), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n865), .A2(KEYINPUT38), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n860), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n842), .B1(new_n868), .B2(KEYINPUT39), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n622), .A2(new_n628), .A3(new_n400), .ZN(new_n870));
  INV_X1    g0670(.A(new_n853), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n852), .A2(new_n853), .A3(new_n397), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n855), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n861), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT99), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n867), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n859), .A2(KEYINPUT99), .A3(KEYINPUT38), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n877), .A2(new_n878), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n869), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT100), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n868), .A2(new_n842), .A3(KEYINPUT39), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n884), .B1(new_n883), .B2(new_n885), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n841), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n629), .A2(new_n658), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n438), .A2(new_n659), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n443), .B(new_n891), .C1(new_n426), .C2(new_n438), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n421), .A2(new_n414), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n425), .A2(G179), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n341), .A2(new_n666), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n897), .B1(new_n822), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n889), .B1(new_n900), .B2(new_n868), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n888), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n454), .A2(new_n693), .A3(new_n696), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n903), .A2(new_n631), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n902), .B(new_n904), .Z(new_n905));
  AND3_X1   g0705(.A1(new_n713), .A2(new_n816), .A3(new_n896), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT40), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n868), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n713), .A2(new_n816), .A3(new_n896), .ZN(new_n909));
  AND4_X1   g0709(.A1(KEYINPUT99), .A2(new_n865), .A3(KEYINPUT38), .A4(new_n866), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT99), .B1(new_n859), .B2(KEYINPUT38), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n909), .B1(new_n912), .B2(new_n877), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n908), .B1(new_n913), .B2(new_n907), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(new_n454), .A3(new_n713), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(G330), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n914), .B1(new_n454), .B2(new_n713), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n905), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n247), .B2(new_n718), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n905), .A2(new_n918), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n840), .B1(new_n920), .B2(new_n921), .ZN(G367));
  AOI21_X1  g0722(.A(new_n737), .B1(new_n681), .B2(new_n329), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n681), .A2(new_n480), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n237), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n722), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(KEYINPUT104), .Z(new_n927));
  AOI21_X1  g0727(.A(new_n480), .B1(new_n767), .B2(G317), .ZN(new_n928));
  OAI221_X1 g0728(.A(new_n928), .B1(new_n461), .B2(new_n745), .C1(new_n746), .C2(new_n761), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(G294), .B2(new_n794), .ZN(new_n930));
  INV_X1    g0730(.A(new_n742), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(KEYINPUT46), .A3(G116), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT46), .B1(new_n931), .B2(G116), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(G107), .B2(new_n750), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n764), .A2(new_n762), .B1(new_n756), .B2(new_n743), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT105), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n930), .A2(new_n932), .A3(new_n934), .A4(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n794), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n938), .A2(new_n772), .B1(new_n219), .B2(new_n761), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT106), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n796), .A2(G77), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n941), .B(new_n266), .C1(new_n286), .C2(new_n756), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(G68), .B2(new_n750), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n931), .A2(G58), .ZN(new_n944));
  INV_X1    g0744(.A(new_n764), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n945), .A2(G143), .B1(new_n767), .B2(G137), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n940), .A2(new_n943), .A3(new_n944), .A4(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n939), .A2(KEYINPUT106), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n937), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT47), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n735), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n949), .A2(new_n950), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n666), .A2(new_n634), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n640), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n638), .B2(new_n954), .ZN(new_n956));
  INV_X1    g0756(.A(new_n727), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n927), .B1(new_n952), .B2(new_n953), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT107), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT102), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n553), .A2(new_n666), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n568), .A2(new_n564), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT101), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n632), .A2(new_n961), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n963), .A2(KEYINPUT101), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n677), .B2(new_n678), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT44), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n677), .A2(new_n678), .A3(new_n969), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT45), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n675), .A2(new_n971), .A3(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n675), .B1(new_n971), .B2(new_n974), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n715), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n670), .A2(new_n676), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n677), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n664), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n665), .A2(new_n980), .A3(new_n677), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n960), .B1(new_n978), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n977), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n975), .ZN(new_n988));
  INV_X1    g0788(.A(new_n985), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n988), .A2(KEYINPUT102), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n715), .B1(new_n986), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n682), .B(KEYINPUT41), .Z(new_n992));
  OAI21_X1  g0792(.A(new_n719), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n969), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(new_n677), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT42), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n569), .B1(new_n994), .B2(new_n540), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n659), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n675), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1005), .A2(new_n994), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1007));
  AND3_X1   g0807(.A1(new_n1004), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1006), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n993), .A2(KEYINPUT103), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(KEYINPUT103), .B1(new_n993), .B2(new_n1010), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n959), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1014), .A2(KEYINPUT108), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(KEYINPUT108), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(G387));
  INV_X1    g0817(.A(new_n750), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n1018), .A2(new_n746), .B1(new_n742), .B2(new_n533), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n756), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1020), .A2(G317), .B1(new_n760), .B2(G303), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n757), .B2(new_n764), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G311), .B2(new_n794), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1019), .B1(new_n1023), .B2(KEYINPUT48), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT110), .Z(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(KEYINPUT48), .B2(new_n1023), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n354), .B1(new_n766), .B2(new_n763), .C1(new_n221), .C2(new_n745), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n767), .A2(G150), .B1(new_n760), .B2(G68), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n219), .B2(new_n756), .C1(new_n284), .C2(new_n754), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n354), .B1(new_n796), .B2(G97), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n269), .B2(new_n742), .C1(new_n772), .C2(new_n764), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1018), .A2(new_n330), .ZN(new_n1035));
  NOR3_X1   g0835(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n735), .B1(new_n1030), .B2(new_n1036), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n234), .A2(new_n471), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n684), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1038), .A2(new_n924), .B1(new_n1039), .B2(new_n729), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n684), .B(new_n471), .C1(new_n281), .C2(new_n269), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT50), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n284), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1042), .B1(new_n1043), .B2(new_n219), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n284), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n1041), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n1040), .A2(new_n1046), .B1(G107), .B2(new_n204), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n722), .B1(new_n1047), .B2(new_n736), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT109), .Z(new_n1049));
  NAND2_X1  g0849(.A1(new_n1037), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n671), .B2(new_n727), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n720), .B2(new_n984), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n715), .A2(new_n982), .A3(new_n983), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n985), .A2(new_n682), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1054), .ZN(G393));
  OAI21_X1  g0855(.A(new_n682), .B1(new_n988), .B2(new_n989), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n986), .B2(new_n990), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n988), .A2(new_n720), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n737), .B1(G97), .B2(new_n681), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n245), .A2(new_n924), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n722), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n742), .A2(new_n281), .B1(new_n766), .B2(new_n802), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n354), .B(new_n1063), .C1(G87), .C2(new_n796), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT112), .Z(new_n1065));
  OAI22_X1  g0865(.A1(new_n764), .A2(new_n286), .B1(new_n756), .B2(new_n772), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1043), .A2(new_n760), .B1(new_n750), .B2(G77), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(new_n219), .C2(new_n938), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G317), .A2(new_n945), .B1(new_n1020), .B2(G311), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT52), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n742), .A2(new_n746), .B1(new_n745), .B2(new_n215), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n761), .A2(new_n533), .B1(new_n766), .B2(new_n757), .ZN(new_n1074));
  NOR4_X1   g0874(.A1(new_n1072), .A2(new_n266), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n794), .A2(G303), .B1(G116), .B2(new_n750), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT113), .Z(new_n1077));
  AOI22_X1  g0877(.A1(new_n1065), .A2(new_n1070), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1062), .B1(new_n739), .B2(new_n1078), .C1(new_n969), .C2(new_n957), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1059), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1058), .A2(new_n1081), .ZN(G390));
  NAND3_X1  g0882(.A1(new_n713), .A2(new_n816), .A3(G330), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n896), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n900), .A2(new_n841), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n886), .A2(new_n887), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n841), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n870), .A2(new_n871), .B1(new_n855), .B2(new_n874), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n880), .B(new_n881), .C1(KEYINPUT38), .C2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n898), .B1(new_n692), .B2(new_n821), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1089), .B(new_n1091), .C1(new_n1092), .C2(new_n897), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1086), .B1(new_n1088), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n883), .A2(new_n885), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(KEYINPUT100), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1085), .B(new_n1093), .C1(new_n1099), .C2(new_n1087), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1095), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n454), .A2(new_n818), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n903), .A2(new_n631), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1083), .A2(new_n897), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1085), .A2(KEYINPUT114), .A3(new_n1092), .A4(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1085), .A2(new_n1092), .A3(new_n1104), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT114), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1085), .A2(new_n1104), .B1(new_n822), .B2(new_n899), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1103), .B(new_n1105), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1101), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1110), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1095), .A2(new_n1100), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1111), .A2(new_n682), .A3(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1099), .A2(new_n726), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n742), .A2(new_n286), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT53), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n266), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G132), .A2(new_n1020), .B1(new_n767), .B2(G125), .ZN(new_n1119));
  INV_X1    g0919(.A(G128), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1119), .B1(new_n219), .B2(new_n745), .C1(new_n1120), .C2(new_n764), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1118), .B(new_n1121), .C1(new_n1117), .C2(new_n1116), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT54), .B(G143), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n761), .A2(new_n1123), .B1(new_n1018), .B2(new_n772), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n794), .B2(G137), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT115), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n794), .A2(G107), .B1(G97), .B2(new_n760), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT116), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n745), .A2(new_n281), .B1(new_n766), .B2(new_n533), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n764), .A2(new_n746), .B1(new_n756), .B2(new_n221), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1129), .B(new_n1130), .C1(G77), .C2(new_n750), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n317), .B1(new_n503), .B2(new_n742), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1132), .A2(KEYINPUT117), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(KEYINPUT117), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1131), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1122), .A2(new_n1126), .B1(new_n1128), .B2(new_n1135), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n721), .B1(new_n1043), .B2(new_n786), .C1(new_n1136), .C2(new_n739), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1115), .A2(new_n1137), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1095), .A2(new_n1100), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n720), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1114), .A2(new_n1140), .ZN(G378));
  NAND2_X1  g0941(.A1(new_n314), .A2(new_n449), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n658), .B1(new_n293), .B2(new_n302), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n314), .A2(new_n449), .A3(new_n1143), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n907), .B1(new_n1091), .B2(new_n906), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n906), .A2(new_n868), .A3(new_n907), .ZN(new_n1154));
  OAI211_X1 g0954(.A(G330), .B(new_n1152), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1152), .B1(new_n914), .B2(G330), .ZN(new_n1157));
  OAI21_X1  g0957(.A(KEYINPUT122), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1158), .A2(new_n888), .A3(new_n901), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT122), .ZN(new_n1160));
  OAI21_X1  g0960(.A(G330), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1152), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1160), .B1(new_n1163), .B2(new_n1155), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1089), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n901), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1159), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n720), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1162), .A2(new_n725), .ZN(new_n1170));
  INV_X1    g0970(.A(G125), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n764), .A2(new_n1171), .B1(new_n754), .B2(new_n806), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n760), .A2(G137), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1173), .B1(new_n1120), .B2(new_n756), .C1(new_n742), .C2(new_n1123), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1172), .B(new_n1174), .C1(G150), .C2(new_n750), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G159), .A2(new_n796), .B1(new_n767), .B2(G124), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(G33), .A2(G41), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT118), .Z(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT120), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1178), .A2(new_n1179), .A3(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G116), .A2(new_n945), .B1(new_n931), .B2(G77), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n750), .A2(G68), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n480), .A2(G41), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n796), .A2(G58), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n461), .A2(new_n754), .B1(new_n756), .B2(new_n215), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n761), .A2(new_n330), .B1(new_n766), .B2(new_n746), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(KEYINPUT58), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT58), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1182), .A2(new_n219), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1195), .B(new_n1196), .C1(new_n1189), .C2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n735), .B1(new_n1186), .B2(new_n1198), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT121), .Z(new_n1200));
  AOI211_X1 g1000(.A(new_n722), .B(new_n1200), .C1(new_n219), .C2(new_n785), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1170), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1169), .A2(KEYINPUT123), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT123), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n719), .B1(new_n1159), .B2(new_n1167), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1202), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1203), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1113), .A2(new_n1103), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT57), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n902), .B1(new_n1157), .B2(new_n1156), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n888), .A2(new_n901), .A3(new_n1163), .A4(new_n1155), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1210), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1209), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n682), .ZN(new_n1215));
  AOI21_X1  g1015(.A(KEYINPUT57), .B1(new_n1209), .B2(new_n1168), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1208), .B1(new_n1215), .B2(new_n1216), .ZN(G375));
  OAI21_X1  g1017(.A(new_n1105), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1218), .A2(new_n719), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n721), .B1(new_n786), .B2(G68), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n931), .A2(G159), .B1(new_n760), .B2(G150), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n806), .B2(new_n764), .C1(new_n938), .C2(new_n1123), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G137), .A2(new_n1020), .B1(new_n767), .B2(G128), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n750), .A2(G50), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1223), .A2(new_n480), .A3(new_n1190), .A4(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1035), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1020), .A2(G283), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1226), .A2(new_n317), .A3(new_n941), .A4(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n945), .A2(G294), .B1(new_n760), .B2(G107), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(G97), .A2(new_n931), .B1(new_n767), .B2(G303), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(new_n938), .C2(new_n221), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n1222), .A2(new_n1225), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1220), .B1(new_n1232), .B2(new_n735), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n896), .B2(new_n726), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1219), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1103), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1218), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n992), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n1238), .A3(new_n1110), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1235), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(G381));
  NAND3_X1  g1041(.A1(new_n1052), .A2(new_n783), .A3(new_n1054), .ZN(new_n1242));
  OR4_X1    g1042(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n1101), .A2(new_n719), .B1(new_n1115), .B2(new_n1137), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n683), .B1(new_n1101), .B2(new_n1110), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1245), .B1(new_n1113), .B2(new_n1246), .ZN(new_n1247));
  OR2_X1    g1047(.A1(G375), .A2(KEYINPUT124), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(G375), .A2(KEYINPUT124), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1244), .A2(new_n1247), .A3(new_n1248), .A4(new_n1249), .ZN(G407));
  NOR2_X1   g1050(.A1(new_n657), .A2(G343), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1248), .A2(new_n1247), .A3(new_n1249), .A4(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(G407), .A2(G213), .A3(new_n1252), .ZN(G409));
  OAI211_X1 g1053(.A(new_n1208), .B(G378), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n1209), .A2(new_n1238), .A3(new_n1168), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1202), .B1(new_n1256), .B2(new_n719), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1247), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1251), .B1(new_n1254), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1110), .A2(KEYINPUT60), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1237), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1218), .A2(KEYINPUT60), .A3(new_n1236), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(new_n682), .A3(new_n1262), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1263), .A2(G384), .A3(new_n1235), .ZN(new_n1264));
  AOI21_X1  g1064(.A(G384), .B1(new_n1263), .B2(new_n1235), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT125), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1251), .A2(G2897), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1266), .A2(new_n1267), .A3(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1268), .B1(new_n1271), .B2(KEYINPUT125), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(KEYINPUT125), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1270), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(KEYINPUT63), .B1(new_n1259), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1259), .A2(new_n1271), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1259), .A2(KEYINPUT63), .A3(new_n1271), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT103), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT102), .B1(new_n988), .B2(new_n989), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n978), .A2(new_n960), .A3(new_n985), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n979), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n720), .B1(new_n1282), .B2(new_n1238), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1010), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1279), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1011), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G393), .A2(G396), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1242), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1288), .B1(new_n1057), .B2(new_n1080), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT108), .B1(new_n1287), .B2(new_n1242), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1289), .B1(G390), .B2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1286), .A2(new_n959), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1291), .B1(new_n1286), .B2(new_n959), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1293), .A2(new_n1294), .A3(KEYINPUT61), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1277), .A2(new_n1278), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT62), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1259), .A2(new_n1297), .A3(new_n1271), .ZN(new_n1298));
  XOR2_X1   g1098(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n1259), .B2(new_n1274), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1297), .B1(new_n1259), .B2(new_n1271), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1298), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1296), .B1(new_n1302), .B2(new_n1303), .ZN(G405));
  NAND2_X1  g1104(.A1(new_n1266), .A2(KEYINPUT127), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1306), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1291), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1014), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1309), .A2(new_n1292), .A3(new_n1305), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1307), .A2(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1254), .B1(KEYINPUT127), .B2(new_n1266), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1312), .B1(G375), .B2(new_n1247), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1311), .B(new_n1313), .ZN(G402));
endmodule


