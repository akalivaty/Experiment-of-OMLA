//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n574, new_n576, new_n577, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n647, new_n648, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(KEYINPUT64), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(new_n453), .B2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(KEYINPUT64), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(KEYINPUT66), .A3(G125), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT65), .B(G2105), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n467), .A2(KEYINPUT67), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n475), .A2(new_n477), .B1(G101), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(KEYINPUT67), .B(G2104), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT68), .B1(new_n484), .B2(new_n465), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n481), .A2(new_n486), .A3(KEYINPUT3), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n465), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(KEYINPUT69), .B1(new_n465), .B2(G2104), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n476), .A2(G137), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n488), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n483), .A2(new_n494), .ZN(G160));
  AOI21_X1  g070(.A(new_n491), .B1(new_n485), .B2(new_n487), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(new_n477), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n497), .B(KEYINPUT70), .ZN(new_n498));
  INV_X1    g073(.A(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n498), .A2(G124), .B1(G136), .B2(new_n501), .ZN(new_n502));
  OAI221_X1 g077(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n476), .C2(G112), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(new_n504), .B(KEYINPUT71), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G162));
  AND3_X1   g081(.A1(new_n499), .A2(G102), .A3(G2104), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n476), .A2(new_n473), .A3(G138), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n476), .A2(G138), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n488), .A2(KEYINPUT4), .A3(new_n492), .A4(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT72), .A2(G114), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT72), .A2(G114), .ZN(new_n514));
  NOR3_X1   g089(.A1(new_n513), .A2(new_n514), .A3(new_n467), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(new_n496), .B2(G126), .ZN(new_n516));
  OAI211_X1 g091(.A(new_n510), .B(new_n512), .C1(new_n516), .C2(new_n499), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(G164));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n520), .B2(G651), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(KEYINPUT73), .A3(KEYINPUT6), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n521), .A2(new_n523), .B1(new_n520), .B2(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT5), .B(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G88), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n521), .A2(new_n523), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n520), .A2(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G50), .ZN(new_n534));
  NAND2_X1  g109(.A1(G75), .A2(G543), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n532), .A2(KEYINPUT5), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT5), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G62), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n535), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G651), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(KEYINPUT74), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n541), .A2(new_n544), .A3(G651), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n528), .A2(new_n534), .A3(new_n543), .A4(new_n545), .ZN(G303));
  INV_X1    g121(.A(G303), .ZN(G166));
  NAND3_X1  g122(.A1(new_n524), .A2(G51), .A3(G543), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n524), .A2(G89), .A3(new_n525), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n550));
  NAND3_X1  g125(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT7), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n548), .A2(new_n549), .A3(new_n550), .A4(new_n552), .ZN(G286));
  INV_X1    g128(.A(G286), .ZN(G168));
  NAND2_X1  g129(.A1(G77), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G64), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n539), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n524), .A2(G52), .A3(G543), .ZN(new_n559));
  INV_X1    g134(.A(G90), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n558), .B(new_n559), .C1(new_n560), .C2(new_n526), .ZN(G301));
  INV_X1    g136(.A(G301), .ZN(G171));
  AOI22_X1  g137(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n563), .A2(new_n522), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n529), .A2(G43), .A3(G543), .A4(new_n530), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n529), .A2(G81), .A3(new_n530), .A4(new_n525), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT75), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n567), .B1(new_n565), .B2(new_n566), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n564), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G860), .ZN(G153));
  AND3_X1   g148(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G36), .ZN(G176));
  NAND2_X1  g150(.A1(G1), .A2(G3), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT8), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n574), .A2(new_n577), .ZN(G188));
  NOR2_X1   g153(.A1(new_n537), .A2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n532), .A2(KEYINPUT5), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT76), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n536), .A2(new_n538), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(G65), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(G78), .A2(G543), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n522), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AND3_X1   g161(.A1(new_n524), .A2(G91), .A3(new_n525), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n529), .A2(G53), .A3(G543), .A4(new_n530), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT9), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n524), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n588), .A2(new_n594), .ZN(G299));
  NAND4_X1  g170(.A1(new_n529), .A2(G87), .A3(new_n530), .A4(new_n525), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT77), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(KEYINPUT78), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n524), .A2(G49), .A3(G543), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT78), .ZN(new_n602));
  OAI211_X1 g177(.A(new_n602), .B(G651), .C1(new_n525), .C2(G74), .ZN(new_n603));
  AND3_X1   g178(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n598), .A2(new_n604), .ZN(G288));
  NAND2_X1  g180(.A1(new_n533), .A2(G48), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n527), .A2(G86), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n525), .A2(G61), .ZN(new_n608));
  NAND2_X1  g183(.A1(G73), .A2(G543), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n522), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT79), .ZN(new_n611));
  AND2_X1   g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n606), .B(new_n607), .C1(new_n612), .C2(new_n613), .ZN(G305));
  INV_X1    g189(.A(G60), .ZN(new_n615));
  INV_X1    g190(.A(G72), .ZN(new_n616));
  OAI22_X1  g191(.A1(new_n539), .A2(new_n615), .B1(new_n616), .B2(new_n532), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT80), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI221_X1 g194(.A(KEYINPUT80), .B1(new_n616), .B2(new_n532), .C1(new_n539), .C2(new_n615), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n619), .A2(G651), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(KEYINPUT81), .ZN(new_n622));
  AOI22_X1  g197(.A1(G85), .A2(new_n527), .B1(new_n533), .B2(G47), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n624));
  NAND4_X1  g199(.A1(new_n619), .A2(new_n624), .A3(new_n620), .A4(G651), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n622), .A2(new_n623), .A3(new_n625), .ZN(G290));
  NAND2_X1  g201(.A1(G301), .A2(G868), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n524), .A2(G92), .A3(new_n525), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT10), .ZN(new_n629));
  AND3_X1   g204(.A1(new_n536), .A2(new_n538), .A3(new_n582), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n582), .B1(new_n536), .B2(new_n538), .ZN(new_n631));
  INV_X1    g206(.A(G66), .ZN(new_n632));
  NOR3_X1   g207(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(G79), .A2(G543), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(G651), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n637));
  AND3_X1   g212(.A1(new_n524), .A2(G54), .A3(G543), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n581), .A2(G66), .A3(new_n583), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n522), .B1(new_n641), .B2(new_n634), .ZN(new_n642));
  OAI21_X1  g217(.A(KEYINPUT82), .B1(new_n642), .B2(new_n638), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n629), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n627), .B1(new_n644), .B2(G868), .ZN(G284));
  OAI21_X1  g220(.A(new_n627), .B1(new_n644), .B2(G868), .ZN(G321));
  NAND2_X1  g221(.A1(G286), .A2(G868), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n593), .A2(new_n586), .A3(new_n587), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n647), .B1(new_n648), .B2(G868), .ZN(G297));
  OAI21_X1  g224(.A(new_n647), .B1(new_n648), .B2(G868), .ZN(G280));
  INV_X1    g225(.A(new_n629), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n637), .B1(new_n636), .B2(new_n639), .ZN(new_n652));
  NOR3_X1   g227(.A1(new_n642), .A2(KEYINPUT82), .A3(new_n638), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n654), .A2(G559), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(G860), .B2(new_n644), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT83), .ZN(G148));
  OAI21_X1  g232(.A(G868), .B1(new_n654), .B2(G559), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(G868), .B2(new_n572), .ZN(G323));
  XNOR2_X1  g234(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g235(.A1(new_n498), .A2(G123), .B1(G135), .B2(new_n501), .ZN(new_n661));
  OAI221_X1 g236(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n476), .C2(G111), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(G2096), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n482), .A2(new_n473), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT13), .B(G2100), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n664), .A2(new_n669), .ZN(G156));
  XNOR2_X1  g245(.A(G2427), .B(G2438), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2430), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT15), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n673), .A2(G2435), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(G2435), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(KEYINPUT14), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1341), .B(G1348), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT16), .B(G2443), .Z(new_n679));
  XNOR2_X1  g254(.A(G2451), .B(G2454), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT85), .B(G2446), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n684), .A2(G14), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT86), .ZN(G401));
  XOR2_X1   g262(.A(G2072), .B(G2078), .Z(new_n688));
  XOR2_X1   g263(.A(G2067), .B(G2678), .Z(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G2084), .B(G2090), .Z(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n688), .B1(new_n692), .B2(KEYINPUT18), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G2096), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(G2100), .Z(new_n695));
  AND2_X1   g270(.A1(new_n692), .A2(KEYINPUT17), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n690), .A2(new_n691), .ZN(new_n697));
  AOI21_X1  g272(.A(KEYINPUT18), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n695), .B(new_n698), .ZN(G227));
  XOR2_X1   g274(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n700));
  XNOR2_X1  g275(.A(G1961), .B(G1966), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT87), .ZN(new_n702));
  XOR2_X1   g277(.A(G1956), .B(G2474), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1971), .B(G1976), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT19), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n700), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n702), .A2(new_n703), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n704), .A2(new_n706), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n704), .A2(new_n700), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(new_n708), .ZN(new_n711));
  OAI221_X1 g286(.A(new_n707), .B1(new_n708), .B2(new_n709), .C1(new_n711), .C2(new_n706), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1986), .ZN(new_n713));
  XOR2_X1   g288(.A(G1991), .B(G1996), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT89), .B(G1981), .Z(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n715), .B(new_n718), .ZN(G229));
  NOR2_X1   g294(.A1(G16), .A2(G23), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n598), .A2(new_n604), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(G16), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT33), .B(G1976), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT91), .B(KEYINPUT92), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G22), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G166), .B2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(G1971), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  MUX2_X1   g306(.A(G6), .B(G305), .S(G16), .Z(new_n732));
  XOR2_X1   g307(.A(KEYINPUT32), .B(G1981), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n726), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT34), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OR2_X1    g312(.A1(G25), .A2(G29), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n498), .A2(G119), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n501), .A2(G131), .ZN(new_n740));
  OAI221_X1 g315(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n476), .C2(G107), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G29), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n738), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n744), .A2(KEYINPUT90), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(KEYINPUT90), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT35), .B(G1991), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n745), .A2(new_n748), .A3(new_n746), .ZN(new_n750));
  MUX2_X1   g325(.A(G24), .B(G290), .S(G16), .Z(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(G1986), .Z(new_n752));
  AND3_X1   g327(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT36), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n737), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n756));
  OAI21_X1  g331(.A(KEYINPUT36), .B1(new_n756), .B2(new_n736), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n743), .A2(G26), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n498), .A2(G128), .B1(G140), .B2(new_n501), .ZN(new_n760));
  OAI221_X1 g335(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n476), .C2(G116), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n760), .A2(KEYINPUT94), .A3(new_n761), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n759), .B1(new_n766), .B2(G29), .ZN(new_n767));
  MUX2_X1   g342(.A(new_n759), .B(new_n767), .S(KEYINPUT28), .Z(new_n768));
  INV_X1    g343(.A(G2067), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT31), .B(G11), .Z(new_n771));
  INV_X1    g346(.A(KEYINPUT24), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n743), .B1(new_n772), .B2(G34), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT97), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n772), .A2(G34), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n773), .A2(new_n774), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G160), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(new_n743), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(G2084), .Z(new_n781));
  INV_X1    g356(.A(new_n663), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n781), .B1(G29), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n727), .A2(G21), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G168), .B2(new_n727), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G1966), .Z(new_n786));
  NAND3_X1  g361(.A1(new_n727), .A2(KEYINPUT23), .A3(G20), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT23), .ZN(new_n788));
  INV_X1    g363(.A(G20), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(G16), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n787), .B(new_n790), .C1(new_n648), .C2(new_n727), .ZN(new_n791));
  INV_X1    g366(.A(G1956), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(G171), .A2(G16), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G5), .B2(G16), .ZN(new_n795));
  INV_X1    g370(.A(G1961), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT99), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n783), .A2(new_n786), .A3(new_n793), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n743), .A2(G32), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n498), .A2(G129), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n482), .A2(G105), .ZN(new_n802));
  NAND3_X1  g377(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT26), .Z(new_n804));
  INV_X1    g379(.A(G141), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n802), .B(new_n804), .C1(new_n500), .C2(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n800), .B1(new_n807), .B2(new_n743), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT27), .B(G1996), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n727), .A2(G19), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n572), .B2(new_n727), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1341), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT98), .B(KEYINPUT30), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G28), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n813), .B1(new_n743), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT95), .B1(G29), .B2(G33), .ZN(new_n817));
  OR3_X1    g392(.A1(KEYINPUT95), .A2(G29), .A3(G33), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT96), .B(KEYINPUT25), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n822));
  INV_X1    g397(.A(G139), .ZN(new_n823));
  OAI221_X1 g398(.A(new_n821), .B1(new_n476), .B2(new_n822), .C1(new_n500), .C2(new_n823), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n817), .B(new_n818), .C1(new_n824), .C2(new_n743), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G2072), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n727), .A2(G4), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n644), .B2(new_n727), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT93), .B(G1348), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n816), .A2(new_n826), .A3(new_n830), .ZN(new_n831));
  OR3_X1    g406(.A1(new_n799), .A2(new_n810), .A3(new_n831), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n770), .A2(new_n771), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n743), .A2(G27), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G164), .B2(new_n743), .ZN(new_n835));
  INV_X1    g410(.A(G2078), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n795), .A2(new_n796), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n758), .A2(new_n833), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(G29), .A2(G35), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G162), .B2(G29), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT29), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(G2090), .Z(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n839), .A2(new_n844), .ZN(G311));
  AND2_X1   g420(.A1(new_n758), .A2(new_n833), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n846), .A2(new_n837), .A3(new_n838), .A4(new_n843), .ZN(G150));
  NAND2_X1  g422(.A1(new_n527), .A2(G93), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n533), .A2(G55), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(new_n522), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(G860), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n571), .A2(KEYINPUT101), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT101), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n857), .B(new_n564), .C1(new_n569), .C2(new_n570), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n571), .A2(KEYINPUT101), .A3(new_n852), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT39), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n644), .A2(G559), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n854), .B1(new_n866), .B2(G860), .ZN(G145));
  XNOR2_X1  g442(.A(new_n807), .B(new_n824), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n764), .A2(new_n517), .A3(new_n765), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n517), .B1(new_n764), .B2(new_n765), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n870), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n868), .B1(new_n874), .B2(new_n871), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n877));
  OR3_X1    g452(.A1(new_n476), .A2(new_n877), .A3(G118), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n476), .B2(G118), .ZN(new_n879));
  OR2_X1    g454(.A1(G106), .A2(G2105), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n878), .A2(new_n879), .A3(G2104), .A4(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G142), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n881), .B1(new_n500), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(new_n498), .B2(G130), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n742), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n742), .A2(new_n884), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n885), .A2(new_n886), .A3(new_n667), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n667), .B1(new_n885), .B2(new_n886), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n876), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n873), .A2(new_n889), .A3(new_n875), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n505), .A2(new_n663), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n505), .A2(new_n663), .ZN(new_n897));
  AOI21_X1  g472(.A(G160), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n897), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n899), .A2(new_n779), .A3(new_n895), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n894), .B(new_n901), .C1(new_n892), .C2(new_n891), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n898), .A2(new_n900), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n891), .A3(new_n893), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g482(.A(new_n861), .B(new_n655), .Z(new_n908));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n648), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(G299), .A2(KEYINPUT104), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n654), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n644), .A2(new_n909), .A3(new_n648), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n908), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n912), .A2(new_n917), .A3(new_n913), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n917), .B1(new_n912), .B2(new_n913), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n916), .B1(new_n920), .B2(new_n908), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n921), .A2(KEYINPUT42), .ZN(new_n922));
  NAND2_X1  g497(.A1(G290), .A2(new_n721), .ZN(new_n923));
  NAND4_X1  g498(.A1(G288), .A2(new_n623), .A3(new_n622), .A4(new_n625), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT105), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(G305), .B(G303), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n923), .A2(KEYINPUT105), .A3(new_n924), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n928), .A2(new_n925), .ZN(new_n929));
  INV_X1    g504(.A(new_n926), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n921), .A2(KEYINPUT42), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n922), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n922), .B2(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(G868), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(G868), .B2(new_n856), .ZN(G295));
  OAI21_X1  g511(.A(new_n935), .B1(G868), .B2(new_n856), .ZN(G331));
  XNOR2_X1  g512(.A(G301), .B(G286), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n859), .A2(new_n939), .A3(new_n860), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n939), .B1(new_n859), .B2(new_n860), .ZN(new_n942));
  OAI22_X1  g517(.A1(new_n918), .A2(new_n919), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n858), .A2(new_n856), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n565), .A2(new_n566), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT75), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n568), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n857), .B1(new_n947), .B2(new_n564), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n860), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n938), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n915), .A2(new_n940), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n931), .A2(new_n943), .A3(new_n952), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n941), .A2(new_n914), .A3(new_n942), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n918), .A2(KEYINPUT108), .B1(new_n940), .B2(new_n951), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n910), .B1(new_n654), .B2(new_n911), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n909), .B1(new_n588), .B2(new_n594), .ZN(new_n957));
  NOR4_X1   g532(.A1(new_n593), .A2(new_n586), .A3(KEYINPUT104), .A4(new_n587), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n644), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT41), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n912), .A2(new_n917), .A3(new_n913), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n954), .B1(new_n955), .B2(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n903), .B(new_n953), .C1(new_n964), .C2(new_n931), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n943), .A2(new_n967), .A3(new_n952), .ZN(new_n968));
  INV_X1    g543(.A(new_n931), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n967), .B1(new_n943), .B2(new_n952), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n903), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT107), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n960), .A2(new_n962), .B1(new_n940), .B2(new_n951), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT106), .B1(new_n974), .B2(new_n954), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n975), .A2(new_n969), .A3(new_n968), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(new_n977), .A3(new_n903), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n973), .A2(new_n953), .A3(new_n978), .ZN(new_n979));
  OAI211_X1 g554(.A(KEYINPUT44), .B(new_n966), .C1(new_n979), .C2(KEYINPUT43), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT109), .B1(new_n965), .B2(KEYINPUT43), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT108), .ZN(new_n983));
  OAI22_X1  g558(.A1(new_n941), .A2(new_n942), .B1(new_n962), .B2(new_n961), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n952), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(G37), .B1(new_n985), .B2(new_n969), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n986), .A2(new_n987), .A3(new_n988), .A4(new_n953), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n982), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n976), .A2(new_n977), .A3(new_n903), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n977), .B1(new_n976), .B2(new_n903), .ZN(new_n993));
  INV_X1    g568(.A(new_n953), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n991), .B1(new_n995), .B2(new_n988), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n981), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n990), .B1(new_n979), .B2(KEYINPUT43), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n999), .A2(KEYINPUT110), .A3(KEYINPUT44), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n980), .B1(new_n998), .B2(new_n1000), .ZN(G397));
  INV_X1    g576(.A(G1384), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n484), .A2(KEYINPUT68), .A3(new_n465), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n486), .B1(new_n481), .B2(KEYINPUT3), .ZN(new_n1004));
  OAI211_X1 g579(.A(G126), .B(new_n492), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n515), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n499), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n512), .A2(new_n510), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT45), .B(new_n1002), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT45), .B1(new_n517), .B2(new_n1002), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT115), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1002), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n475), .A2(new_n477), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n482), .A2(G101), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1017), .A2(new_n494), .A3(G40), .A4(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n483), .A2(KEYINPUT111), .A3(G40), .A4(new_n494), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1015), .A2(new_n1016), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(KEYINPUT56), .B(G2072), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1012), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n648), .B(KEYINPUT57), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1013), .A2(KEYINPUT50), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n517), .A2(new_n1029), .A3(new_n1002), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n792), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1025), .A2(new_n1026), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1025), .A2(new_n1032), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1026), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1031), .A2(new_n829), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1007), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n512), .A2(new_n510), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1384), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1028), .A2(new_n1041), .A3(new_n769), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n654), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1033), .B1(new_n1037), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1036), .A2(new_n1033), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT61), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1036), .A2(KEYINPUT61), .A3(new_n1033), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1038), .A2(KEYINPUT60), .A3(new_n1042), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(KEYINPUT122), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(KEYINPUT122), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n644), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(KEYINPUT122), .A3(new_n654), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1050), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT60), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1047), .B(new_n1048), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1012), .A2(new_n1023), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1057), .B1(new_n1058), .B2(G1996), .ZN(new_n1059));
  XOR2_X1   g634(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n1060));
  XNOR2_X1  g635(.A(new_n1060), .B(G1341), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n1062), .B2(new_n1013), .ZN(new_n1063));
  INV_X1    g638(.A(G1996), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1012), .A2(new_n1023), .A3(KEYINPUT120), .A4(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1059), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n572), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(KEYINPUT59), .A3(new_n572), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1044), .B1(new_n1056), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G8), .ZN(new_n1073));
  NOR2_X1   g648(.A1(G168), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1062), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1076));
  OAI22_X1  g651(.A1(new_n1076), .A2(G1966), .B1(G2084), .B2(new_n1031), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  OAI211_X1 g653(.A(KEYINPUT51), .B(new_n1075), .C1(new_n1078), .C2(new_n1073), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1080), .B(G8), .C1(new_n1077), .C2(G286), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1078), .A2(KEYINPUT123), .A3(new_n1075), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n1077), .B2(new_n1074), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1079), .B(new_n1081), .C1(new_n1082), .C2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1012), .A2(new_n1023), .A3(new_n836), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1031), .A2(new_n796), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1019), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1093), .A2(KEYINPUT124), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1088), .A2(G2078), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(KEYINPUT124), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1092), .A2(new_n1094), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  AND4_X1   g672(.A1(G301), .A2(new_n1089), .A3(new_n1091), .A4(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1090), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1076), .A2(new_n1095), .ZN(new_n1100));
  AOI21_X1  g675(.A(G301), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1086), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1089), .A2(new_n1091), .A3(new_n1097), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(G171), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT125), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1099), .A2(G301), .A3(new_n1100), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1104), .A2(new_n1105), .A3(KEYINPUT54), .A4(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1073), .B1(new_n1028), .B2(new_n1041), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n607), .A2(new_n606), .ZN(new_n1109));
  OAI21_X1  g684(.A(G1981), .B1(new_n1109), .B2(new_n610), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(G305), .B2(G1981), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT49), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(KEYINPUT117), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1108), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1112), .B1(new_n1111), .B2(KEYINPUT117), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n721), .A2(G1976), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(KEYINPUT116), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1108), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1119), .B1(new_n1108), .B2(new_n1117), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OR3_X1    g697(.A1(new_n721), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1116), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(G303), .A2(G8), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(KEYINPUT55), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1031), .A2(G2090), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(new_n1058), .B2(new_n730), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1128), .B2(new_n1073), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1126), .ZN(new_n1130));
  AOI21_X1  g705(.A(G1971), .B1(new_n1012), .B2(new_n1023), .ZN(new_n1131));
  OAI211_X1 g706(.A(G8), .B(new_n1130), .C1(new_n1131), .C2(new_n1127), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1124), .A2(new_n1129), .A3(new_n1132), .ZN(new_n1133));
  AND4_X1   g708(.A1(new_n1085), .A2(new_n1102), .A3(new_n1107), .A4(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1104), .A2(KEYINPUT54), .A3(new_n1106), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT125), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1072), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1085), .A2(KEYINPUT62), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1085), .A2(KEYINPUT62), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1138), .A2(new_n1101), .A3(new_n1139), .A4(new_n1133), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT63), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1129), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1077), .A2(G8), .A3(G168), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1128), .A2(new_n1073), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1142), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1147), .A2(new_n1124), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1141), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1116), .A2(G1976), .A3(G288), .ZN(new_n1150));
  NOR2_X1   g725(.A1(G305), .A2(G1981), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT118), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1108), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1144), .A2(KEYINPUT63), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n1130), .B2(new_n1146), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1153), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1149), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1137), .A2(new_n1140), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT112), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n1062), .B2(new_n1015), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1011), .A2(KEYINPUT112), .A3(new_n1028), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1163), .A2(KEYINPUT114), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1163), .A2(KEYINPUT114), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n742), .A2(new_n748), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n742), .A2(new_n748), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1166), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n766), .A2(G2067), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n764), .A2(new_n769), .A3(new_n765), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1170), .B(new_n1171), .C1(new_n1064), .C2(new_n807), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1166), .A2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1163), .A2(G1996), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(new_n807), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1169), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(KEYINPUT113), .B1(G290), .B2(G1986), .ZN(new_n1177));
  NAND2_X1  g752(.A1(G290), .A2(G1986), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1177), .B(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1179), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1159), .A2(new_n1176), .A3(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1173), .A2(new_n1168), .A3(new_n1175), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n1171), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(KEYINPUT126), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1182), .A2(new_n1185), .A3(new_n1171), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1184), .A2(new_n1166), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1170), .A2(new_n807), .A3(new_n1171), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1166), .A2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g764(.A1(KEYINPUT127), .A2(KEYINPUT46), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1174), .B(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(KEYINPUT127), .A2(KEYINPUT46), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1189), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT47), .ZN(new_n1194));
  NOR3_X1   g769(.A1(new_n1163), .A2(G1986), .A3(G290), .ZN(new_n1195));
  XOR2_X1   g770(.A(new_n1195), .B(KEYINPUT48), .Z(new_n1196));
  NAND2_X1  g771(.A1(new_n1176), .A2(new_n1196), .ZN(new_n1197));
  AND3_X1   g772(.A1(new_n1187), .A2(new_n1194), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1181), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g774(.A1(G229), .A2(G227), .ZN(new_n1201));
  NOR2_X1   g775(.A1(new_n999), .A2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g776(.A1(G401), .A2(new_n462), .ZN(new_n1203));
  NAND3_X1  g777(.A1(new_n1202), .A2(new_n906), .A3(new_n1203), .ZN(G225));
  INV_X1    g778(.A(G225), .ZN(G308));
endmodule


