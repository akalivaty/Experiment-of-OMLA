//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1172, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n204));
  AOI22_X1  g0004(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n205), .A2(KEYINPUT68), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(KEYINPUT68), .ZN(new_n207));
  OAI21_X1  g0007(.A(new_n204), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT69), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT67), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G77), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n203), .B1(new_n209), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT1), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n203), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n220), .B(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT65), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n222), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT66), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n218), .A2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G264), .ZN(new_n237));
  INV_X1    g0037(.A(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n248), .B1(G41), .B2(G45), .ZN(new_n249));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G97), .ZN(new_n252));
  INV_X1    g0052(.A(G232), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G1698), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(G226), .B2(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n252), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n251), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n262), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n249), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n263), .B1(new_n213), .B2(new_n265), .ZN(new_n266));
  OR2_X1    g0066(.A1(new_n266), .A2(KEYINPUT13), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(KEYINPUT13), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G169), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT14), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n267), .A2(G179), .A3(new_n268), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n224), .A2(G33), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT70), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n276), .A2(G77), .B1(G20), .B2(new_n212), .ZN(new_n277));
  INV_X1    g0077(.A(G50), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n223), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  XOR2_X1   g0084(.A(new_n284), .B(KEYINPUT11), .Z(new_n285));
  AND2_X1   g0085(.A1(new_n282), .A2(new_n223), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(G1), .B2(new_n224), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT12), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n248), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n288), .B1(new_n290), .B2(new_n212), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n289), .A2(KEYINPUT12), .A3(G68), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n287), .A2(new_n212), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n285), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n274), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g0096(.A(KEYINPUT8), .B(G58), .Z(new_n297));
  NAND2_X1  g0097(.A1(new_n276), .A2(new_n297), .ZN(new_n298));
  NOR3_X1   g0098(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n299));
  INV_X1    g0099(.A(G150), .ZN(new_n300));
  OAI221_X1 g0100(.A(new_n298), .B1(new_n224), .B2(new_n299), .C1(new_n300), .C2(new_n280), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n301), .A2(new_n283), .B1(new_n278), .B2(new_n290), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n283), .A2(KEYINPUT71), .B1(new_n248), .B2(G20), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(KEYINPUT71), .B2(new_n283), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n304), .A2(new_n278), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n265), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G226), .ZN(new_n308));
  INV_X1    g0108(.A(new_n251), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT3), .B(G33), .ZN(new_n310));
  INV_X1    g0110(.A(G1698), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G222), .ZN(new_n312));
  INV_X1    g0112(.A(G223), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n310), .B(new_n312), .C1(new_n313), .C2(new_n311), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n314), .B(new_n262), .C1(G77), .C2(new_n310), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n308), .A2(new_n309), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G169), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n316), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n306), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n306), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n323), .A2(KEYINPUT9), .B1(G190), .B2(new_n319), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT10), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT9), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n306), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n316), .A2(G200), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n324), .A2(new_n325), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G190), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n328), .B1(new_n330), .B2(new_n316), .C1(new_n306), .C2(new_n326), .ZN(new_n331));
  INV_X1    g0131(.A(new_n327), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT10), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n322), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n269), .A2(G200), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT74), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n335), .B(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n337), .B(new_n294), .C1(new_n330), .C2(new_n269), .ZN(new_n338));
  OR3_X1    g0138(.A1(new_n287), .A2(KEYINPUT73), .A3(new_n214), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT73), .B1(new_n287), .B2(new_n214), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n297), .A2(new_n279), .B1(G20), .B2(G77), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT15), .B(G87), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n341), .B1(new_n275), .B2(new_n342), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n339), .A2(new_n340), .B1(new_n343), .B2(new_n283), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n289), .A2(G77), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT72), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n260), .B1(G232), .B2(new_n311), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n213), .B2(new_n311), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n349), .B(new_n262), .C1(G107), .C2(new_n310), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n251), .B1(new_n307), .B2(G244), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n347), .B1(G190), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G200), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n353), .B1(new_n354), .B2(new_n352), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n296), .A2(new_n334), .A3(new_n338), .A4(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT75), .B1(new_n256), .B2(KEYINPUT3), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT75), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(new_n258), .A3(G33), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n257), .ZN(new_n361));
  XOR2_X1   g0161(.A(KEYINPUT76), .B(KEYINPUT7), .Z(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(new_n224), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n258), .A2(G33), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n357), .B2(new_n359), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(G20), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n363), .B(G68), .C1(new_n364), .C2(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(G58), .B(G68), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n369), .A2(G20), .B1(G159), .B2(new_n279), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(KEYINPUT16), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT16), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT7), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n310), .B2(G20), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n260), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n212), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n370), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n372), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n371), .A2(new_n378), .A3(new_n283), .ZN(new_n379));
  MUX2_X1   g0179(.A(new_n289), .B(new_n304), .S(new_n297), .Z(new_n380));
  AND2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G33), .A2(G87), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n382), .B(KEYINPUT77), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n366), .B1(G226), .B2(new_n311), .ZN(new_n384));
  NOR2_X1   g0184(.A1(G223), .A2(G1698), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n262), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n265), .A2(new_n253), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n309), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G200), .ZN(new_n391));
  AOI211_X1 g0191(.A(new_n251), .B(new_n388), .C1(new_n386), .C2(new_n262), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G190), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n381), .A2(KEYINPUT17), .A3(new_n391), .A4(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n393), .A2(new_n391), .A3(new_n379), .A4(new_n380), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT17), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n379), .A2(new_n380), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n387), .A2(G179), .A3(new_n309), .A4(new_n389), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n392), .B2(new_n317), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n398), .A2(KEYINPUT18), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT18), .B1(new_n398), .B2(new_n400), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n394), .B(new_n397), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n352), .A2(G169), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n352), .A2(new_n320), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n347), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n356), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT5), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT81), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(G41), .ZN(new_n411));
  INV_X1    g0211(.A(G45), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(G1), .ZN(new_n413));
  INV_X1    g0213(.A(G41), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n411), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n264), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(new_n238), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n366), .B1(G264), .B2(new_n311), .ZN(new_n419));
  NOR2_X1   g0219(.A1(G257), .A2(G1698), .ZN(new_n420));
  INV_X1    g0220(.A(G303), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n419), .A2(new_n420), .B1(new_n421), .B2(new_n310), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n418), .B1(new_n422), .B2(new_n262), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n416), .A2(new_n250), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G200), .ZN(new_n427));
  INV_X1    g0227(.A(G116), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(G20), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n283), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT85), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G283), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n432), .B(KEYINPUT80), .ZN(new_n433));
  AOI21_X1  g0233(.A(G20), .B1(new_n256), .B2(G97), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT20), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n430), .A2(KEYINPUT85), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT85), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(new_n283), .B2(new_n429), .ZN(new_n439));
  OAI211_X1 g0239(.A(KEYINPUT20), .B(new_n435), .C1(new_n437), .C2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n289), .A2(G116), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT86), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n286), .B(new_n289), .C1(G1), .C2(new_n256), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(KEYINPUT84), .A3(G116), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT84), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n446), .B2(new_n428), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n427), .A2(new_n444), .A3(new_n445), .A4(new_n451), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n423), .A2(new_n425), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G190), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n354), .B1(new_n423), .B2(new_n425), .ZN(new_n455));
  INV_X1    g0255(.A(new_n443), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n451), .B(new_n456), .C1(new_n436), .C2(new_n441), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT86), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n452), .A2(new_n454), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n310), .A2(new_n224), .A3(G87), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT22), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT23), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n224), .B2(G107), .ZN(new_n464));
  INV_X1    g0264(.A(G107), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(KEYINPUT23), .A3(G20), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n461), .A2(new_n462), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n366), .A2(KEYINPUT22), .A3(new_n224), .A4(G87), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n224), .A2(G33), .A3(G116), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT24), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT24), .A4(new_n469), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(new_n283), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n447), .A2(G107), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n289), .A2(G107), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n476), .B(KEYINPUT25), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G250), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n311), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n366), .B(new_n480), .C1(G257), .C2(new_n311), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G294), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n264), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n264), .A2(new_n416), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n484), .A2(G264), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n425), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n317), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(new_n320), .A3(new_n425), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n478), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n457), .A2(new_n426), .A3(G169), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT21), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n453), .A2(G179), .A3(new_n457), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n457), .A2(new_n426), .A3(KEYINPUT21), .A4(G169), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n490), .A2(new_n493), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT82), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n215), .A2(KEYINPUT4), .A3(G1698), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n257), .A2(new_n259), .A3(G244), .A4(new_n311), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n366), .A2(new_n499), .B1(new_n500), .B2(KEYINPUT4), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n310), .A2(G250), .A3(G1698), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n433), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n262), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n424), .B1(new_n484), .B2(G257), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(G179), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n317), .B1(new_n504), .B2(new_n505), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n289), .A2(G97), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(new_n447), .B2(G97), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT7), .B1(new_n260), .B2(new_n224), .ZN(new_n513));
  AOI211_X1 g0313(.A(new_n373), .B(G20), .C1(new_n257), .C2(new_n259), .ZN(new_n514));
  OAI21_X1  g0314(.A(G107), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT78), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n465), .A2(KEYINPUT6), .A3(G97), .ZN(new_n518));
  XOR2_X1   g0318(.A(G97), .B(G107), .Z(new_n519));
  OAI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(KEYINPUT6), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n520), .A2(G20), .B1(G77), .B2(new_n279), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n374), .A2(new_n375), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n522), .A2(KEYINPUT78), .A3(G107), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n517), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n512), .B1(new_n524), .B2(new_n283), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n498), .B1(new_n509), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n504), .A2(new_n505), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G169), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n506), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT78), .B1(new_n522), .B2(G107), .ZN(new_n530));
  AOI211_X1 g0330(.A(new_n516), .B(new_n465), .C1(new_n374), .C2(new_n375), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n286), .B1(new_n532), .B2(new_n521), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n529), .B(KEYINPUT82), .C1(new_n533), .C2(new_n512), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n526), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n342), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(new_n289), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n366), .A2(new_n224), .A3(G68), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT19), .ZN(new_n539));
  INV_X1    g0339(.A(G97), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n539), .B1(new_n275), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n224), .B1(new_n252), .B2(new_n539), .ZN(new_n542));
  XNOR2_X1  g0342(.A(new_n542), .B(KEYINPUT83), .ZN(new_n543));
  NOR3_X1   g0343(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n538), .B(new_n541), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n537), .B1(new_n545), .B2(new_n283), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n447), .A2(G87), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n413), .A2(new_n250), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n264), .B(new_n549), .C1(G250), .C2(new_n413), .ZN(new_n550));
  NOR2_X1   g0350(.A1(G238), .A2(G1698), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n215), .B2(G1698), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n366), .A2(new_n552), .B1(G33), .B2(G116), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n550), .B1(new_n553), .B2(new_n264), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(new_n330), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(G200), .B2(new_n554), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n447), .A2(new_n536), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n546), .A2(new_n557), .B1(new_n317), .B2(new_n554), .ZN(new_n558));
  OR2_X1    g0358(.A1(new_n554), .A2(G179), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n548), .A2(new_n556), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n527), .A2(new_n354), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(G190), .B2(new_n527), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n524), .A2(new_n283), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT79), .B1(new_n563), .B2(new_n511), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT79), .ZN(new_n565));
  AOI211_X1 g0365(.A(new_n565), .B(new_n512), .C1(new_n524), .C2(new_n283), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n562), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n474), .A2(new_n477), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n487), .A2(G200), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n486), .A2(G190), .A3(new_n425), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n568), .A2(new_n475), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n535), .A2(new_n560), .A3(new_n567), .A4(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  AND4_X1   g0373(.A1(new_n408), .A2(new_n460), .A3(new_n497), .A4(new_n573), .ZN(G372));
  INV_X1    g0374(.A(KEYINPUT26), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT88), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n564), .A2(new_n566), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(new_n529), .ZN(new_n578));
  NOR4_X1   g0378(.A1(new_n564), .A2(new_n566), .A3(new_n509), .A4(KEYINPUT88), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n575), .B(new_n560), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n558), .A2(new_n559), .ZN(new_n581));
  INV_X1    g0381(.A(new_n560), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT26), .B1(new_n582), .B2(new_n535), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n565), .B1(new_n533), .B2(new_n512), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n525), .A2(KEYINPUT79), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n587), .A2(new_n562), .B1(new_n526), .B2(new_n534), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT87), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n588), .A2(new_n589), .A3(new_n560), .A4(new_n571), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n572), .A2(KEYINPUT87), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(new_n591), .A3(new_n496), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n584), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n408), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT89), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n401), .B2(new_n402), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n398), .A2(new_n400), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT18), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n398), .A2(new_n400), .A3(KEYINPUT18), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(KEYINPUT89), .A3(new_n600), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n294), .B1(new_n272), .B2(new_n273), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n338), .B1(new_n603), .B2(new_n407), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n394), .A2(new_n397), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n602), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n329), .A2(new_n333), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n322), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n594), .A2(new_n609), .ZN(G369));
  NAND3_X1  g0410(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n459), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(G13), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n613), .A2(G20), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n248), .ZN(new_n615));
  XNOR2_X1  g0415(.A(KEYINPUT90), .B(KEYINPUT27), .ZN(new_n616));
  OR2_X1    g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(G213), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(G343), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n457), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g0422(.A(new_n622), .B(KEYINPUT91), .Z(new_n623));
  MUX2_X1   g0423(.A(new_n611), .B(new_n612), .S(new_n623), .Z(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(G330), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n478), .A2(new_n621), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n571), .A2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n628), .A2(new_n490), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n490), .A2(new_n621), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n621), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n611), .A2(new_n633), .ZN(new_n634));
  OAI22_X1  g0434(.A1(new_n629), .A2(new_n634), .B1(new_n490), .B2(new_n621), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n632), .A2(new_n636), .ZN(G399));
  INV_X1    g0437(.A(new_n219), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n638), .A2(G41), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n544), .A2(new_n428), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(G1), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n227), .B2(new_n640), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n643), .B(KEYINPUT28), .ZN(new_n644));
  INV_X1    g0444(.A(G330), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n453), .A2(G179), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n646), .A2(new_n487), .A3(new_n554), .A4(new_n527), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n483), .A2(new_n554), .A3(new_n485), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n453), .A2(new_n507), .A3(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n649), .A2(KEYINPUT30), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(KEYINPUT30), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT92), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT92), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n654), .B(new_n647), .C1(new_n650), .C2(new_n651), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n653), .A2(new_n621), .A3(new_n655), .ZN(new_n656));
  NOR4_X1   g0456(.A1(new_n572), .A2(new_n459), .A3(new_n496), .A4(new_n621), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT31), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n652), .A2(KEYINPUT31), .A3(new_n621), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n645), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n621), .B1(new_n584), .B2(new_n592), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT29), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n560), .A2(new_n526), .A3(new_n575), .A4(new_n534), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n664), .A2(new_n581), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n585), .A2(new_n529), .A3(new_n586), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT88), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n577), .A2(new_n576), .A3(new_n529), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n582), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n665), .B1(new_n669), .B2(new_n575), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n572), .A2(new_n497), .ZN(new_n671));
  OAI211_X1 g0471(.A(KEYINPUT29), .B(new_n633), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n661), .B1(new_n663), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n644), .B1(new_n673), .B2(G1), .ZN(G364));
  NAND2_X1  g0474(.A1(new_n614), .A2(G45), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n640), .A2(G1), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n626), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(G330), .B2(new_n624), .ZN(new_n679));
  NOR2_X1   g0479(.A1(G13), .A2(G33), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G20), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n677), .B1(new_n624), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n223), .B1(G20), .B2(new_n317), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n243), .A2(G45), .ZN(new_n687));
  XOR2_X1   g0487(.A(new_n687), .B(KEYINPUT93), .Z(new_n688));
  NOR2_X1   g0488(.A1(new_n366), .A2(new_n638), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(G45), .B2(new_n227), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT94), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n638), .A2(new_n260), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n688), .A2(new_n691), .B1(G355), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(G116), .B2(new_n219), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n684), .B1(new_n686), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n224), .A2(G190), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT95), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n697), .A2(G179), .A3(G200), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n699), .A2(KEYINPUT96), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(KEYINPUT96), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G159), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT32), .ZN(new_n705));
  NOR2_X1   g0505(.A1(G179), .A2(G200), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n224), .B1(new_n706), .B2(G190), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n707), .A2(KEYINPUT98), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(KEYINPUT98), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n330), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI22_X1  g0513(.A1(new_n710), .A2(new_n540), .B1(new_n278), .B2(new_n713), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n697), .A2(G179), .A3(new_n354), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G107), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n224), .A2(new_n330), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n354), .A2(G179), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G87), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n716), .A2(new_n310), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT97), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n711), .A2(G190), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n714), .B(new_n723), .C1(G68), .C2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(G58), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n320), .A2(G200), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n717), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n725), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n727), .A2(new_n696), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI211_X1 g0531(.A(new_n705), .B(new_n729), .C1(G77), .C2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G311), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G329), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n702), .A2(new_n735), .B1(new_n421), .B2(new_n719), .ZN(new_n736));
  INV_X1    g0536(.A(new_n710), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n734), .B(new_n736), .C1(G294), .C2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n728), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G322), .ZN(new_n740));
  INV_X1    g0540(.A(G317), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n741), .A2(KEYINPUT33), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(KEYINPUT33), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n724), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n310), .B1(new_n715), .B2(G283), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n738), .A2(new_n740), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(G326), .B2(new_n712), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n685), .B1(new_n732), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n695), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n679), .A2(new_n749), .ZN(G396));
  NAND2_X1  g0550(.A1(new_n347), .A2(new_n621), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n355), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n406), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n407), .A2(new_n633), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n662), .B(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n677), .B1(new_n759), .B2(new_n661), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n760), .A2(KEYINPUT100), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n759), .A2(new_n661), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(KEYINPUT100), .A3(new_n676), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n761), .B(new_n763), .C1(new_n661), .C2(new_n759), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n758), .A2(new_n680), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n739), .A2(G143), .B1(G150), .B2(new_n724), .ZN(new_n766));
  INV_X1    g0566(.A(G137), .ZN(new_n767));
  INV_X1    g0567(.A(G159), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n766), .B1(new_n767), .B2(new_n713), .C1(new_n768), .C2(new_n730), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT34), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n361), .B1(new_n703), .B2(G132), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n769), .A2(new_n770), .B1(G68), .B2(new_n715), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n772), .B(new_n773), .C1(new_n726), .C2(new_n710), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n771), .B(new_n774), .C1(G50), .C2(new_n720), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n310), .B1(new_n720), .B2(G107), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(KEYINPUT99), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n778), .B1(new_n540), .B2(new_n710), .C1(new_n702), .C2(new_n733), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n715), .A2(G87), .B1(G294), .B2(new_n739), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n780), .B1(KEYINPUT99), .B2(new_n777), .C1(new_n428), .C2(new_n730), .ZN(new_n781));
  INV_X1    g0581(.A(new_n724), .ZN(new_n782));
  INV_X1    g0582(.A(G283), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n713), .A2(new_n421), .ZN(new_n785));
  NOR4_X1   g0585(.A1(new_n779), .A2(new_n781), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n685), .B1(new_n775), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n685), .A2(new_n680), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n214), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n765), .A2(new_n787), .A3(new_n677), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n764), .A2(new_n790), .ZN(G384));
  INV_X1    g0591(.A(KEYINPUT40), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n605), .A2(new_n596), .A3(new_n601), .ZN(new_n793));
  INV_X1    g0593(.A(new_n619), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n398), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n597), .A2(new_n795), .A3(new_n395), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(KEYINPUT37), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT37), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n597), .A2(new_n795), .A3(new_n395), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(KEYINPUT38), .B1(new_n797), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n371), .A2(new_n283), .ZN(new_n805));
  AOI21_X1  g0605(.A(KEYINPUT16), .B1(new_n368), .B2(new_n370), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n380), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n403), .A2(new_n794), .A3(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n395), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n400), .A2(new_n794), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(new_n810), .B2(new_n807), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n801), .B1(new_n811), .B2(new_n800), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n808), .A2(new_n812), .A3(KEYINPUT38), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n792), .B1(new_n804), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n633), .B1(new_n652), .B2(KEYINPUT92), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n815), .A2(KEYINPUT31), .A3(new_n655), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n758), .B1(new_n659), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n295), .A2(new_n621), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n296), .A2(new_n338), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n603), .A2(new_n621), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n814), .A2(new_n817), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n808), .A2(new_n812), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT38), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n813), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n817), .A2(new_n826), .A3(new_n821), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n792), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n822), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n659), .A2(new_n816), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n408), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT101), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n829), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(G330), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n819), .A2(new_n820), .ZN(new_n835));
  AND3_X1   g0635(.A1(new_n590), .A2(new_n591), .A3(new_n496), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n633), .B(new_n757), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n835), .B1(new_n838), .B2(new_n755), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n826), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT39), .ZN(new_n841));
  INV_X1    g0641(.A(new_n813), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n841), .B1(new_n803), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n296), .A2(new_n621), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n825), .A2(KEYINPUT39), .A3(new_n813), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n602), .A2(new_n794), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n840), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n408), .B(new_n672), .C1(new_n662), .C2(KEYINPUT29), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n609), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n848), .B(new_n850), .Z(new_n851));
  XNOR2_X1  g0651(.A(new_n834), .B(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n248), .B2(new_n614), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n428), .B1(new_n520), .B2(KEYINPUT35), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n854), .B(new_n226), .C1(KEYINPUT35), .C2(new_n520), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT36), .ZN(new_n856));
  OAI21_X1  g0656(.A(G77), .B1(new_n726), .B2(new_n212), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n857), .A2(new_n227), .B1(G50), .B2(new_n212), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n858), .A2(G1), .A3(new_n613), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n853), .A2(new_n856), .A3(new_n859), .ZN(G367));
  OAI21_X1  g0660(.A(new_n560), .B1(new_n548), .B2(new_n633), .ZN(new_n861));
  OR3_X1    g0661(.A1(new_n581), .A2(new_n548), .A3(new_n633), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n863), .A2(KEYINPUT43), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n588), .B1(new_n587), .B2(new_n633), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n577), .A2(new_n529), .A3(new_n621), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n535), .B1(new_n868), .B2(new_n490), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n633), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n866), .A2(new_n867), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n871), .A2(new_n631), .A3(new_n611), .A4(new_n633), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT42), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT102), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT102), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n870), .A2(new_n876), .A3(new_n873), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n875), .B(new_n877), .C1(KEYINPUT42), .C2(new_n872), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n863), .A2(KEYINPUT43), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n865), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n632), .A2(new_n868), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n878), .A2(new_n865), .A3(new_n879), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n878), .A2(new_n865), .A3(new_n879), .ZN(new_n885));
  OAI22_X1  g0685(.A1(new_n885), .A2(new_n880), .B1(new_n632), .B2(new_n868), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n639), .B(KEYINPUT41), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  OR3_X1    g0688(.A1(new_n868), .A2(new_n635), .A3(KEYINPUT103), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT103), .B1(new_n868), .B2(new_n635), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT45), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n868), .A2(new_n635), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT44), .Z(new_n895));
  NAND3_X1  g0695(.A1(new_n889), .A2(KEYINPUT45), .A3(new_n890), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n893), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n632), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n893), .A2(new_n895), .A3(new_n632), .A4(new_n896), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n625), .A2(KEYINPUT104), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n631), .B(new_n634), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n625), .A2(KEYINPUT104), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n902), .B2(new_n901), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n899), .A2(new_n673), .A3(new_n900), .A4(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n888), .B1(new_n906), .B2(new_n673), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n675), .A2(G1), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n884), .B(new_n886), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT105), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n703), .A2(G137), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n737), .A2(G68), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n715), .A2(G77), .B1(G150), .B2(new_n739), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n310), .B1(new_n730), .B2(new_n278), .ZN(new_n914));
  INV_X1    g0714(.A(G143), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n713), .A2(new_n915), .B1(new_n719), .B2(new_n726), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n914), .B(new_n916), .C1(G159), .C2(new_n724), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n911), .A2(new_n912), .A3(new_n913), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n703), .A2(G317), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n731), .A2(G283), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n366), .B1(new_n739), .B2(G303), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n719), .A2(new_n428), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n922), .A2(KEYINPUT46), .B1(G311), .B2(new_n712), .ZN(new_n923));
  INV_X1    g0723(.A(G294), .ZN(new_n924));
  OAI221_X1 g0724(.A(new_n923), .B1(KEYINPUT46), .B2(new_n922), .C1(new_n924), .C2(new_n782), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(G97), .B2(new_n715), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n919), .A2(new_n920), .A3(new_n921), .A4(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n710), .A2(new_n465), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n918), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT47), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n685), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n861), .A2(new_n862), .A3(new_n682), .ZN(new_n932));
  INV_X1    g0732(.A(new_n689), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n686), .B1(new_n219), .B2(new_n342), .C1(new_n239), .C2(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n931), .A2(new_n677), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n909), .A2(new_n910), .A3(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n910), .B1(new_n909), .B2(new_n935), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n937), .A2(new_n938), .ZN(G387));
  NAND2_X1  g0739(.A1(new_n905), .A2(new_n908), .ZN(new_n940));
  INV_X1    g0740(.A(new_n715), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n361), .B1(new_n941), .B2(new_n428), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n737), .A2(G283), .B1(G294), .B2(new_n720), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n739), .A2(G317), .B1(G311), .B2(new_n724), .ZN(new_n944));
  INV_X1    g0744(.A(G322), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n944), .B1(new_n421), .B2(new_n730), .C1(new_n945), .C2(new_n713), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT48), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT107), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n946), .A2(new_n947), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT49), .Z(new_n952));
  AOI211_X1 g0752(.A(new_n942), .B(new_n952), .C1(G326), .C2(new_n703), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n703), .A2(G150), .B1(G97), .B2(new_n715), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n720), .A2(G77), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n955), .B1(new_n730), .B2(new_n212), .C1(new_n278), .C2(new_n728), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n297), .B2(new_n724), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n954), .B(new_n957), .C1(new_n768), .C2(new_n713), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n710), .A2(new_n342), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n958), .A2(new_n361), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n685), .B1(new_n953), .B2(new_n960), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n641), .B(new_n412), .C1(new_n212), .C2(new_n214), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT106), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n297), .A2(new_n278), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT50), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n689), .B1(new_n235), .B2(new_n412), .C1(new_n963), .C2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n692), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n966), .B1(G107), .B2(new_n219), .C1(new_n641), .C2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n676), .B1(new_n968), .B2(new_n686), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n961), .B(new_n969), .C1(new_n631), .C2(new_n683), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n905), .A2(new_n673), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n639), .B1(new_n905), .B2(new_n673), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n940), .B(new_n970), .C1(new_n972), .C2(new_n973), .ZN(G393));
  NAND2_X1  g0774(.A1(new_n899), .A2(new_n900), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n971), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(new_n639), .A3(new_n906), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n899), .A2(new_n908), .A3(new_n900), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n686), .B1(new_n540), .B2(new_n219), .C1(new_n246), .C2(new_n933), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n715), .A2(G87), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n980), .B(new_n366), .C1(new_n214), .C2(new_n710), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n713), .A2(new_n300), .B1(new_n728), .B2(new_n768), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT51), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n278), .B2(new_n782), .C1(new_n702), .C2(new_n915), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n981), .B(new_n984), .C1(G68), .C2(new_n720), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n731), .A2(new_n297), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n739), .A2(G311), .B1(G317), .B2(new_n712), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT52), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n260), .B(new_n716), .C1(new_n702), .C2(new_n945), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(G283), .C2(new_n720), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n737), .A2(G116), .B1(G294), .B2(new_n731), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n421), .B2(new_n782), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT108), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n985), .A2(new_n986), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n685), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n677), .B(new_n979), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n996), .A2(KEYINPUT109), .B1(new_n682), .B2(new_n868), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(KEYINPUT109), .B2(new_n996), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n977), .A2(new_n978), .A3(new_n998), .ZN(G390));
  NAND3_X1  g0799(.A1(new_n408), .A2(new_n830), .A3(G330), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n849), .A2(new_n609), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n573), .A2(new_n460), .A3(new_n497), .A4(new_n633), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n1003), .A2(KEYINPUT31), .B1(new_n655), .B2(new_n815), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n816), .ZN(new_n1005));
  OAI211_X1 g0805(.A(G330), .B(new_n757), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n835), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n661), .A2(new_n757), .A3(new_n821), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n633), .B1(new_n670), .B2(new_n671), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n755), .B1(new_n1009), .B2(new_n754), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n1007), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n756), .B1(new_n662), .B2(new_n757), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n660), .ZN(new_n1014));
  OAI21_X1  g0814(.A(G330), .B1(new_n1004), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n835), .B1(new_n1015), .B2(new_n758), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n817), .A2(G330), .A3(new_n821), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1013), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1002), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT111), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n843), .A2(new_n845), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n839), .B2(new_n844), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n844), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n803), .B2(new_n842), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n1011), .B2(new_n835), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1022), .A2(new_n1026), .A3(new_n1008), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1024), .B1(new_n821), .B2(new_n1010), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1023), .B1(new_n1013), .B2(new_n835), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1028), .B1(new_n1029), .B2(new_n1021), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1027), .B1(new_n1030), .B2(new_n1017), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT110), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n1031), .B2(new_n1019), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1013), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1006), .A2(new_n835), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n821), .B1(new_n661), .B2(new_n757), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1007), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1001), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n1035), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1039), .A2(new_n1041), .A3(KEYINPUT110), .A4(new_n1027), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1020), .A2(new_n1031), .B1(new_n1033), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n639), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT114), .ZN(new_n1045));
  AND3_X1   g0845(.A1(new_n1022), .A2(new_n1008), .A3(new_n1026), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1017), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT112), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1048), .A2(new_n1049), .A3(new_n908), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n908), .ZN(new_n1051));
  OAI21_X1  g0851(.A(KEYINPUT112), .B1(new_n1031), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n681), .B1(new_n843), .B2(new_n845), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n788), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1055), .A2(new_n297), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n260), .B1(new_n715), .B2(G50), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n720), .A2(new_n1058), .A3(G150), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1058), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n719), .B2(new_n300), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1057), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n703), .B2(G125), .ZN(new_n1063));
  INV_X1    g0863(.A(G132), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(KEYINPUT54), .B(G143), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n728), .A2(new_n1064), .B1(new_n730), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n737), .B2(G159), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1063), .B(new_n1067), .C1(new_n767), .C2(new_n782), .ZN(new_n1068));
  INV_X1    g0868(.A(G128), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n713), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n721), .B1(new_n713), .B2(new_n783), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n710), .A2(new_n214), .B1(new_n465), .B2(new_n782), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(G68), .C2(new_n715), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n310), .B1(new_n731), .B2(G97), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1073), .B(new_n1074), .C1(new_n924), .C2(new_n702), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n728), .A2(new_n428), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1068), .A2(new_n1070), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n685), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NOR4_X1   g0879(.A1(new_n1054), .A2(new_n676), .A3(new_n1056), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1045), .B1(new_n1053), .B2(new_n1081), .ZN(new_n1082));
  AOI211_X1 g0882(.A(KEYINPUT114), .B(new_n1080), .C1(new_n1050), .C2(new_n1052), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1044), .B1(new_n1082), .B2(new_n1083), .ZN(G378));
  XOR2_X1   g0884(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1085));
  XNOR2_X1  g0885(.A(new_n334), .B(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n323), .A2(new_n619), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1086), .B(new_n1087), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n817), .A2(new_n821), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1089), .A2(new_n814), .B1(new_n827), .B2(new_n792), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1088), .B1(new_n1090), .B2(G330), .ZN(new_n1091));
  AND4_X1   g0891(.A1(G330), .A2(new_n822), .A3(new_n828), .A4(new_n1088), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n848), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1088), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n829), .B2(new_n645), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1090), .A2(G330), .A3(new_n1088), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n848), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1093), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1033), .A2(new_n1042), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n1002), .ZN(new_n1101));
  OAI21_X1  g0901(.A(KEYINPUT118), .B1(new_n1101), .B2(KEYINPUT57), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n640), .B1(new_n1101), .B2(KEYINPUT57), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT118), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT57), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1001), .B1(new_n1033), .B2(new_n1042), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1104), .B(new_n1105), .C1(new_n1106), .C2(new_n1099), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1102), .A2(new_n1103), .A3(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1094), .A2(new_n681), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n715), .A2(G58), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT115), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n713), .A2(new_n428), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n912), .A2(new_n361), .A3(new_n955), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n414), .B1(new_n730), .B2(new_n342), .C1(new_n782), .C2(new_n540), .ZN(new_n1115));
  NOR4_X1   g0915(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1116), .B1(new_n465), .B2(new_n728), .C1(new_n783), .C2(new_n702), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT58), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n360), .A2(G33), .ZN(new_n1119));
  AOI21_X1  g0919(.A(G50), .B1(new_n1119), .B2(new_n414), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n719), .A2(new_n1065), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n737), .A2(G150), .B1(KEYINPUT117), .B2(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n731), .A2(G137), .B1(G132), .B2(new_n724), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT116), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n712), .A2(G125), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n1121), .A2(KEYINPUT117), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(G128), .B2(new_n739), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT59), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(G41), .B1(new_n703), .B2(G124), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n256), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G159), .B2(new_n715), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1120), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n995), .B1(new_n1118), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1055), .A2(G50), .ZN(new_n1138));
  NOR4_X1   g0938(.A1(new_n1109), .A2(new_n676), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1099), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1139), .B1(new_n1140), .B2(new_n908), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1108), .A2(new_n1141), .ZN(G375));
  NAND3_X1  g0942(.A1(new_n1037), .A2(new_n1001), .A3(new_n1038), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1020), .A2(new_n887), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n959), .B1(new_n703), .B2(G303), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1145), .B1(new_n214), .B2(new_n941), .C1(new_n540), .C2(new_n719), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n713), .A2(new_n924), .B1(new_n730), .B2(new_n465), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G116), .B2(new_n724), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT119), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n783), .B2(new_n728), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1146), .A2(new_n310), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1111), .B1(new_n702), .B2(new_n1069), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n713), .A2(new_n1064), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n782), .A2(new_n1065), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n361), .B1(G150), .B2(new_n731), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G137), .A2(new_n739), .B1(new_n720), .B2(G159), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(new_n710), .C2(new_n278), .ZN(new_n1157));
  NOR4_X1   g0957(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .A4(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n685), .B1(new_n1151), .B2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n677), .B(new_n1159), .C1(new_n821), .C2(new_n681), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n212), .B2(new_n788), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1161), .B1(new_n1162), .B2(new_n908), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1144), .A2(new_n1163), .ZN(G381));
  XOR2_X1   g0964(.A(G375), .B(KEYINPUT120), .Z(new_n1165));
  INV_X1    g0965(.A(new_n1082), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1083), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1166), .A2(new_n1167), .B1(new_n639), .B2(new_n1043), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(G387), .A2(G384), .A3(G381), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(G390), .A2(G396), .A3(G393), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1165), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(G407));
  NAND3_X1  g0971(.A1(new_n1165), .A2(new_n620), .A3(new_n1168), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(G407), .A2(G213), .A3(new_n1172), .ZN(G409));
  NAND3_X1  g0973(.A1(new_n1108), .A2(G378), .A3(new_n1141), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT122), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT110), .B1(new_n1048), .B2(new_n1039), .ZN(new_n1176));
  AND4_X1   g0976(.A1(KEYINPUT110), .A2(new_n1039), .A3(new_n1041), .A4(new_n1027), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1002), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1178), .A2(new_n887), .A3(new_n1140), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1139), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT121), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1099), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1093), .A2(new_n1098), .A3(KEYINPUT121), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1182), .A2(new_n908), .A3(new_n1183), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1179), .A2(new_n1180), .A3(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1175), .B1(new_n1185), .B2(G378), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1179), .A2(new_n1180), .A3(new_n1184), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1168), .A2(KEYINPUT122), .A3(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1174), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n620), .A2(G213), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT60), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n640), .B1(new_n1143), .B2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1192), .B(new_n1019), .C1(new_n1191), .C2(new_n1143), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n1163), .ZN(new_n1194));
  INV_X1    g0994(.A(G384), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(G384), .A2(new_n1193), .A3(new_n1163), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT123), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1196), .A2(KEYINPUT123), .A3(new_n1197), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1189), .A2(new_n1190), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(KEYINPUT62), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n620), .A2(G213), .A3(G2897), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1200), .A2(new_n1206), .A3(new_n1201), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1198), .A2(new_n1206), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1205), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT61), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT62), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1189), .A2(new_n1212), .A3(new_n1190), .A4(new_n1202), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1204), .A2(new_n1210), .A3(new_n1211), .A4(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT126), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(G390), .A2(new_n1215), .ZN(new_n1216));
  OR2_X1    g1016(.A1(G390), .A2(new_n1215), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(new_n937), .C2(new_n938), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(G393), .B(G396), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n909), .A2(new_n935), .A3(G390), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1219), .ZN(new_n1222));
  AOI21_X1  g1022(.A(G390), .B1(new_n909), .B2(new_n935), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT125), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(new_n1224), .B2(new_n1220), .ZN(new_n1225));
  AOI211_X1 g1025(.A(KEYINPUT125), .B(G390), .C1(new_n909), .C2(new_n935), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1222), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1221), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1214), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT127), .B1(new_n1228), .B2(new_n1211), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT127), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1232), .B(KEYINPUT61), .C1(new_n1221), .C2(new_n1227), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1189), .A2(new_n1190), .A3(new_n1202), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT63), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT63), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT124), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1207), .A2(new_n1238), .A3(new_n1208), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1238), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1237), .B1(new_n1241), .B2(new_n1205), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1234), .B(new_n1236), .C1(new_n1242), .C2(new_n1235), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1230), .A2(new_n1243), .ZN(G405));
  NAND2_X1  g1044(.A1(G375), .A2(new_n1168), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1174), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1202), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1198), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1247), .B1(new_n1248), .B2(new_n1246), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(new_n1229), .ZN(G402));
endmodule


