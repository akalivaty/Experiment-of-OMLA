//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1104, new_n1105, new_n1106;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT68), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT69), .Z(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(KEYINPUT70), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n470), .A2(new_n472), .A3(KEYINPUT3), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n476), .A2(G137), .A3(new_n477), .A4(new_n463), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  AND3_X1   g055(.A1(new_n476), .A2(new_n477), .A3(new_n463), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n477), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n476), .A2(G2105), .A3(new_n463), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT71), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n485), .B1(G124), .B2(new_n487), .ZN(new_n488));
  XOR2_X1   g063(.A(new_n488), .B(KEYINPUT72), .Z(G162));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n490), .A2(new_n477), .A3(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n466), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n477), .A2(G138), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n476), .A2(new_n463), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n492), .B1(new_n494), .B2(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n476), .A2(G126), .A3(G2105), .A4(new_n463), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n498), .A2(KEYINPUT73), .A3(G2105), .ZN(new_n499));
  AOI21_X1  g074(.A(KEYINPUT73), .B1(new_n498), .B2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(G2104), .B(new_n497), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  OR2_X1    g077(.A1(new_n495), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(KEYINPUT74), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .A3(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G62), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT76), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n511), .A2(new_n512), .B1(G75), .B2(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n513), .B1(new_n512), .B2(new_n511), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT75), .B(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n521), .B2(G50), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n515), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  AND2_X1   g099(.A1(new_n518), .A2(G89), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n526), .B(new_n528), .C1(new_n520), .C2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n525), .A2(new_n530), .ZN(G168));
  AOI22_X1  g106(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n533));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  OR3_X1    g109(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n532), .B2(new_n534), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n518), .A2(G90), .B1(new_n521), .B2(G52), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  AOI22_X1  g114(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n534), .ZN(new_n541));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  INV_X1    g117(.A(G43), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n517), .A2(new_n542), .B1(new_n520), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT78), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n541), .A2(new_n545), .A3(KEYINPUT78), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  AOI22_X1  g131(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n534), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT79), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n521), .A2(G53), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n560), .B1(new_n521), .B2(G53), .ZN(new_n562));
  AND3_X1   g137(.A1(new_n518), .A2(KEYINPUT80), .A3(G91), .ZN(new_n563));
  AOI21_X1  g138(.A(KEYINPUT80), .B1(new_n518), .B2(G91), .ZN(new_n564));
  OAI221_X1 g139(.A(new_n558), .B1(new_n561), .B2(new_n562), .C1(new_n563), .C2(new_n564), .ZN(G299));
  INV_X1    g140(.A(G168), .ZN(G286));
  NAND2_X1  g141(.A1(new_n518), .A2(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n521), .A2(G49), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(G288));
  AOI22_X1  g145(.A1(new_n518), .A2(G86), .B1(new_n521), .B2(G48), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n572), .A2(new_n534), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(G305));
  AOI22_X1  g149(.A1(new_n518), .A2(G85), .B1(new_n521), .B2(G47), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT81), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n534), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT82), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n576), .A2(KEYINPUT82), .A3(new_n578), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n518), .A2(G92), .ZN(new_n585));
  XOR2_X1   g160(.A(KEYINPUT83), .B(KEYINPUT10), .Z(new_n586));
  XNOR2_X1  g161(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(new_n510), .ZN(new_n589));
  INV_X1    g164(.A(G66), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(G54), .B2(new_n521), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n584), .B1(new_n594), .B2(G868), .ZN(G284));
  OAI21_X1  g170(.A(new_n584), .B1(new_n594), .B2(G868), .ZN(G321));
  INV_X1    g171(.A(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(G299), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(new_n597), .B2(G168), .ZN(G297));
  OAI21_X1  g174(.A(new_n598), .B1(new_n597), .B2(G168), .ZN(G280));
  NOR2_X1   g175(.A1(new_n593), .A2(G559), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(G860), .B2(new_n594), .ZN(new_n602));
  XOR2_X1   g177(.A(new_n602), .B(KEYINPUT84), .Z(G148));
  NAND2_X1  g178(.A1(new_n550), .A2(new_n597), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n601), .B(KEYINPUT85), .Z(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n597), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT86), .Z(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g183(.A1(new_n487), .A2(G123), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n477), .A2(G111), .ZN(new_n610));
  OAI21_X1  g185(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n481), .A2(G135), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(G2096), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(G2096), .ZN(new_n616));
  INV_X1    g191(.A(new_n466), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(new_n473), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT87), .B(KEYINPUT13), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n619), .B(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n615), .A2(new_n616), .A3(new_n622), .ZN(G156));
  INV_X1    g198(.A(KEYINPUT14), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2430), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n627), .B2(new_n626), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n629), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  AND3_X1   g212(.A1(new_n636), .A2(G14), .A3(new_n637), .ZN(G401));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT17), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT88), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  INV_X1    g219(.A(new_n642), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n644), .B1(new_n645), .B2(new_n639), .ZN(new_n646));
  AOI22_X1  g221(.A1(new_n641), .A2(new_n642), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n643), .B2(new_n646), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT89), .Z(new_n649));
  INV_X1    g224(.A(new_n639), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n650), .A2(new_n644), .A3(new_n642), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT18), .Z(new_n652));
  NAND3_X1  g227(.A1(new_n640), .A2(new_n644), .A3(new_n645), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n649), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2096), .B(G2100), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(G227));
  XOR2_X1   g231(.A(G1971), .B(G1976), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1961), .B(G1966), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n658), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n658), .A2(new_n661), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  AOI211_X1 g241(.A(new_n663), .B(new_n666), .C1(new_n658), .C2(new_n662), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G229));
  MUX2_X1   g248(.A(G6), .B(G305), .S(G16), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT32), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G1981), .ZN(new_n676));
  NAND2_X1  g251(.A1(G166), .A2(G16), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(G16), .B2(G22), .ZN(new_n678));
  INV_X1    g253(.A(G1971), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  MUX2_X1   g256(.A(G23), .B(G288), .S(G16), .Z(new_n682));
  XOR2_X1   g257(.A(KEYINPUT33), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NOR4_X1   g259(.A1(new_n676), .A2(new_n680), .A3(new_n681), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT34), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n581), .A2(new_n582), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G16), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G16), .B2(G24), .ZN(new_n689));
  INV_X1    g264(.A(G1986), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n691), .A2(KEYINPUT93), .A3(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT35), .B(G1991), .Z(new_n694));
  OR2_X1    g269(.A1(G25), .A2(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n481), .A2(G131), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n477), .A2(G107), .ZN(new_n697));
  OAI21_X1  g272(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G119), .B2(new_n487), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT91), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT92), .Z(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n695), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n693), .B1(new_n694), .B2(new_n704), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n704), .A2(new_n694), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n686), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT36), .ZN(new_n708));
  NOR2_X1   g283(.A1(G4), .A2(G16), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n594), .B2(G16), .ZN(new_n710));
  INV_X1    g285(.A(G1348), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n487), .A2(G129), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n481), .A2(G141), .ZN(new_n714));
  NAND3_X1  g289(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT26), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n473), .A2(G105), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n713), .A2(new_n714), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  MUX2_X1   g293(.A(G32), .B(new_n718), .S(G29), .Z(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT27), .B(G1996), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT97), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n712), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n703), .A2(G27), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G164), .B2(new_n703), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT98), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n609), .A2(G29), .A3(new_n613), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n724), .A2(G2078), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n725), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n727), .B(new_n728), .C1(G2078), .C2(new_n724), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT24), .B(G34), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(new_n703), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT96), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n479), .B2(new_n703), .ZN(new_n733));
  INV_X1    g308(.A(G2084), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G16), .ZN(new_n736));
  NOR2_X1   g311(.A1(G168), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n736), .B2(G21), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n735), .B1(new_n739), .B2(G1966), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n733), .A2(new_n734), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n481), .A2(G139), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT25), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n617), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n742), .B(new_n745), .C1(new_n477), .C2(new_n746), .ZN(new_n747));
  MUX2_X1   g322(.A(G33), .B(new_n747), .S(G29), .Z(new_n748));
  XOR2_X1   g323(.A(KEYINPUT95), .B(G2072), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT30), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n751), .A2(G28), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n703), .B1(new_n751), .B2(G28), .ZN(new_n753));
  AND2_X1   g328(.A1(KEYINPUT31), .A2(G11), .ZN(new_n754));
  NOR2_X1   g329(.A1(KEYINPUT31), .A2(G11), .ZN(new_n755));
  OAI22_X1  g330(.A1(new_n752), .A2(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G1966), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n756), .B1(new_n738), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n740), .A2(new_n741), .A3(new_n750), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n703), .A2(G26), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT28), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n487), .A2(G128), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n477), .A2(G116), .ZN(new_n763));
  OAI21_X1  g338(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n481), .A2(G140), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n761), .B1(new_n767), .B2(G29), .ZN(new_n768));
  INV_X1    g343(.A(G2067), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NOR4_X1   g345(.A1(new_n722), .A2(new_n729), .A3(new_n759), .A4(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G29), .A2(G35), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G162), .B2(G29), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT29), .B(G2090), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(G1961), .ZN(new_n776));
  NOR2_X1   g351(.A1(G5), .A2(G16), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT99), .Z(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G301), .B2(new_n736), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n719), .A2(new_n721), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n736), .A2(G20), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT23), .Z(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G299), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1956), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n780), .B(new_n784), .C1(new_n776), .C2(new_n779), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n773), .A2(new_n774), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n736), .A2(G19), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n551), .B2(new_n736), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT94), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1341), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n771), .A2(new_n775), .A3(new_n787), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT100), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n708), .A2(new_n793), .ZN(G150));
  INV_X1    g369(.A(G150), .ZN(G311));
  NAND2_X1  g370(.A1(new_n594), .A2(G559), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT38), .ZN(new_n797));
  NAND2_X1  g372(.A1(G80), .A2(G543), .ZN(new_n798));
  INV_X1    g373(.A(G67), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n589), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n534), .B1(new_n800), .B2(KEYINPUT101), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(KEYINPUT101), .B2(new_n800), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n518), .A2(G93), .B1(new_n521), .B2(G55), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n802), .A2(new_n546), .A3(new_n803), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n550), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(KEYINPUT102), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT102), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n808), .B(new_n804), .C1(new_n805), .C2(new_n550), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n797), .B(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(KEYINPUT39), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT103), .ZN(new_n813));
  AOI21_X1  g388(.A(G860), .B1(new_n811), .B2(KEYINPUT39), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n805), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G860), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n815), .A2(new_n819), .ZN(G145));
  NAND2_X1  g395(.A1(new_n481), .A2(G142), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n477), .A2(G118), .ZN(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G130), .B2(new_n487), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(new_n619), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n718), .B(new_n747), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n767), .B(new_n503), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n701), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n828), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n614), .B(G160), .ZN(new_n832));
  XNOR2_X1  g407(.A(G162), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n831), .B(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT105), .B(G37), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g412(.A(new_n810), .B(KEYINPUT106), .Z(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(new_n605), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n605), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n593), .B(G299), .Z(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n842), .B(KEYINPUT41), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n839), .A2(new_n840), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n687), .A2(G303), .ZN(new_n847));
  NAND2_X1  g422(.A1(G290), .A2(G166), .ZN(new_n848));
  XOR2_X1   g423(.A(G288), .B(KEYINPUT107), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G305), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n850), .B1(new_n847), .B2(new_n848), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT42), .Z(new_n854));
  AND3_X1   g429(.A1(new_n844), .A2(new_n846), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n854), .B1(new_n844), .B2(new_n846), .ZN(new_n856));
  OAI21_X1  g431(.A(G868), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(G868), .B2(new_n805), .ZN(G295));
  OAI21_X1  g433(.A(new_n857), .B1(G868), .B2(new_n805), .ZN(G331));
  INV_X1    g434(.A(new_n853), .ZN(new_n860));
  XNOR2_X1  g435(.A(G301), .B(G168), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n810), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n842), .ZN(new_n863));
  INV_X1    g438(.A(new_n861), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n807), .A2(new_n809), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT109), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n807), .A2(KEYINPUT109), .A3(new_n809), .A4(new_n864), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n845), .B1(new_n862), .B2(new_n865), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n860), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n862), .A2(new_n842), .A3(new_n865), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n867), .A2(new_n868), .B1(new_n810), .B2(new_n861), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n853), .B(new_n872), .C1(new_n845), .C2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n871), .A2(new_n874), .A3(new_n835), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT43), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n872), .B1(new_n873), .B2(new_n845), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n860), .ZN(new_n878));
  INV_X1    g453(.A(G37), .ZN(new_n879));
  XNOR2_X1  g454(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .A4(new_n874), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n876), .A2(KEYINPUT44), .A3(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT111), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n878), .A2(new_n879), .A3(new_n874), .ZN(new_n886));
  INV_X1    g461(.A(new_n880), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT110), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n871), .A2(new_n874), .A3(new_n835), .A4(new_n880), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n888), .B1(new_n891), .B2(KEYINPUT110), .ZN(new_n892));
  OAI22_X1  g467(.A1(new_n884), .A2(new_n885), .B1(new_n892), .B2(KEYINPUT44), .ZN(G397));
  XOR2_X1   g468(.A(new_n701), .B(new_n694), .Z(new_n894));
  NAND2_X1  g469(.A1(new_n767), .A2(G2067), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n762), .A2(new_n769), .A3(new_n766), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(G1996), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n718), .B(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n894), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(KEYINPUT112), .B(G1384), .Z(new_n901));
  NAND2_X1  g476(.A1(new_n503), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT45), .B1(new_n902), .B2(KEYINPUT113), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(KEYINPUT113), .B2(new_n902), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n469), .A2(G40), .A3(new_n478), .A4(new_n474), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT114), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n900), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n687), .A3(new_n690), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n911), .B1(KEYINPUT48), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(KEYINPUT48), .B2(new_n913), .ZN(new_n915));
  INV_X1    g490(.A(new_n897), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n909), .B1(new_n916), .B2(new_n718), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n909), .A2(new_n898), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n918), .A2(KEYINPUT46), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(KEYINPUT46), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT47), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n899), .A2(new_n694), .A3(new_n897), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n896), .B1(new_n702), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n909), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n915), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT63), .ZN(new_n927));
  NAND2_X1  g502(.A1(G303), .A2(G8), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT55), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  OAI211_X1 g505(.A(KEYINPUT45), .B(new_n901), .C1(new_n495), .C2(new_n502), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT115), .ZN(new_n932));
  INV_X1    g507(.A(G1384), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(new_n495), .B2(new_n502), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n932), .A2(new_n907), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT116), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT116), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n932), .A2(new_n939), .A3(new_n907), .A4(new_n936), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n679), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n934), .A2(KEYINPUT117), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT117), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n943), .B(new_n933), .C1(new_n495), .C2(new_n502), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT50), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n946), .B(new_n907), .C1(KEYINPUT50), .C2(new_n934), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n941), .B1(G2090), .B2(new_n947), .ZN(new_n948));
  XOR2_X1   g523(.A(KEYINPUT119), .B(G8), .Z(new_n949));
  AOI21_X1  g524(.A(new_n930), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G1981), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n952), .B1(new_n571), .B2(new_n573), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n571), .A2(new_n573), .A3(new_n952), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT49), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n955), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT49), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n957), .A2(new_n958), .A3(new_n953), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n945), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n907), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n962), .A3(new_n949), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT120), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n962), .A2(new_n949), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n966), .A2(KEYINPUT120), .A3(new_n960), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1976), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n966), .B1(new_n969), .B2(G288), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT52), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT52), .B1(G288), .B2(new_n969), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n966), .B(new_n972), .C1(new_n969), .C2(G288), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n968), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G8), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n942), .A2(new_n976), .A3(new_n944), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n934), .A2(KEYINPUT50), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n907), .A3(new_n978), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n979), .A2(G2090), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n975), .B1(new_n941), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT118), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n981), .A2(new_n982), .A3(new_n930), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n982), .B1(new_n981), .B2(new_n930), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n951), .B(new_n974), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n475), .A2(new_n906), .A3(G40), .A4(new_n478), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n905), .A2(KEYINPUT114), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n987), .B(new_n988), .C1(new_n935), .C2(new_n934), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT45), .B1(new_n942), .B2(new_n944), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n757), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n991), .B1(new_n979), .B2(G2084), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n949), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n993), .A2(G286), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n927), .B1(new_n986), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(KEYINPUT63), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n941), .A2(new_n980), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(G8), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n997), .B1(new_n929), .B2(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n1000), .B(new_n974), .C1(new_n985), .C2(new_n984), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n996), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT118), .B1(new_n999), .B2(new_n929), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1003), .A2(new_n983), .A3(new_n974), .ZN(new_n1004));
  AOI211_X1 g579(.A(G1976), .B(G288), .C1(new_n965), .C2(new_n967), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n966), .B1(new_n1005), .B2(new_n957), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n992), .A2(G286), .A3(new_n949), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n992), .A2(G8), .ZN(new_n1009));
  NAND2_X1  g584(.A1(G286), .A2(new_n949), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n1010), .B(KEYINPUT126), .Z(new_n1011));
  OAI211_X1 g586(.A(KEYINPUT51), .B(new_n1008), .C1(new_n1009), .C2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n993), .A2(new_n1013), .A3(new_n1010), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1012), .A2(KEYINPUT62), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT62), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n1017));
  OR4_X1    g592(.A1(new_n1017), .A2(new_n989), .A3(new_n990), .A4(G2078), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT121), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n942), .A2(new_n976), .A3(new_n944), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n987), .A2(new_n978), .A3(new_n988), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n977), .A2(new_n907), .A3(KEYINPUT121), .A4(new_n978), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n776), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(G2078), .B1(new_n938), .B2(new_n940), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1018), .B(new_n1024), .C1(new_n1025), .C2(KEYINPUT53), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G171), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1015), .A2(new_n1016), .A3(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n968), .A2(new_n971), .A3(new_n973), .ZN(new_n1029));
  AOI211_X1 g604(.A(new_n1029), .B(new_n950), .C1(new_n1003), .C2(new_n983), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1007), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1002), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n905), .A2(new_n1017), .A3(G2078), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n904), .A2(new_n932), .A3(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1024), .B(new_n1035), .C1(new_n1025), .C2(KEYINPUT53), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1027), .B1(G171), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1033), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OR2_X1    g614(.A1(new_n1026), .A2(G171), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT127), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1036), .A2(new_n1041), .A3(G171), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1041), .B1(new_n1036), .B2(G171), .ZN(new_n1043));
  OAI211_X1 g618(.A(KEYINPUT54), .B(new_n1040), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1030), .A2(new_n1039), .A3(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1022), .A2(new_n711), .A3(new_n1023), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n961), .A2(new_n769), .A3(new_n907), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT122), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT122), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1046), .A2(new_n1050), .A3(new_n1047), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n594), .B1(new_n1052), .B2(KEYINPUT60), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT124), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n1052), .B2(KEYINPUT60), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1046), .A2(new_n1050), .A3(new_n1047), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1050), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1054), .B(KEYINPUT60), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1053), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT60), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n593), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT60), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT124), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1063), .A2(new_n1065), .A3(new_n1058), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT61), .ZN(new_n1067));
  INV_X1    g642(.A(G1956), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n947), .A2(new_n1068), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n932), .A2(new_n907), .A3(new_n936), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT56), .B(G2072), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  XOR2_X1   g647(.A(G299), .B(KEYINPUT57), .Z(new_n1073));
  AND3_X1   g648(.A1(new_n1069), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1073), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1067), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1073), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1069), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(KEYINPUT61), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1076), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n551), .B1(KEYINPUT123), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1070), .A2(new_n898), .ZN(new_n1085));
  XOR2_X1   g660(.A(KEYINPUT58), .B(G1341), .Z(new_n1086));
  NAND2_X1  g661(.A1(new_n962), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1084), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1083), .A2(KEYINPUT123), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1088), .B(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1082), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1060), .A2(new_n1066), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1079), .B1(new_n1052), .B2(new_n593), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1080), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT125), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1045), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1092), .A2(KEYINPUT125), .A3(new_n1094), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1032), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(G290), .B(new_n690), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n910), .B1(new_n900), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n926), .B1(new_n1099), .B2(new_n1101), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g677(.A(G319), .ZN(new_n1104));
  NOR4_X1   g678(.A1(G229), .A2(new_n1104), .A3(G401), .A4(G227), .ZN(new_n1105));
  NAND2_X1  g679(.A1(new_n1105), .A2(new_n836), .ZN(new_n1106));
  NOR2_X1   g680(.A1(new_n892), .A2(new_n1106), .ZN(G308));
  INV_X1    g681(.A(G308), .ZN(G225));
endmodule


