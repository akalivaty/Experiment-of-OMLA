//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1028, new_n1029, new_n1030, new_n1031;
  INV_X1    g000(.A(KEYINPUT103), .ZN(new_n202));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT7), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G92gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT98), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G85gat), .ZN(new_n210));
  INV_X1    g009(.A(G85gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(KEYINPUT98), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n208), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G99gat), .ZN(new_n214));
  INV_X1    g013(.A(G106gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT8), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT99), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n211), .A2(KEYINPUT98), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n209), .A2(G85gat), .ZN(new_n219));
  AOI21_X1  g018(.A(G92gat), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT99), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT8), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n222), .B1(G99gat), .B2(G106gat), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n220), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n207), .B1(new_n217), .B2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(G99gat), .B(G106gat), .Z(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G64gat), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n228), .A2(G57gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(G57gat), .ZN(new_n230));
  AND2_X1   g029(.A1(G71gat), .A2(G78gat), .ZN(new_n231));
  OAI22_X1  g030(.A1(new_n229), .A2(new_n230), .B1(KEYINPUT9), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G71gat), .B(G78gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n221), .B1(new_n220), .B2(new_n223), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT98), .B(G85gat), .ZN(new_n236));
  OAI211_X1 g035(.A(KEYINPUT99), .B(new_n216), .C1(new_n236), .C2(G92gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n226), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n239), .A3(new_n207), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n227), .A2(new_n234), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n234), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n239), .B1(new_n238), .B2(new_n207), .ZN(new_n243));
  AOI211_X1 g042(.A(new_n226), .B(new_n206), .C1(new_n235), .C2(new_n237), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT101), .B(KEYINPUT10), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n241), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n227), .A2(KEYINPUT10), .A3(new_n234), .A4(new_n240), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n204), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n203), .B1(new_n241), .B2(new_n245), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n202), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT102), .B(G176gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(G204gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(G120gat), .B(G148gat), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n253), .B(new_n254), .Z(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n202), .B(new_n255), .C1(new_n249), .C2(new_n250), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G113gat), .B(G120gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n260), .A2(KEYINPUT1), .ZN(new_n261));
  XNOR2_X1  g060(.A(G127gat), .B(G134gat), .ZN(new_n262));
  OR2_X1    g061(.A1(KEYINPUT73), .A2(KEYINPUT1), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n263), .B(new_n262), .C1(new_n260), .C2(KEYINPUT1), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G183gat), .A2(G190gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT24), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n269), .B1(new_n270), .B2(KEYINPUT64), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT64), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n272), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n273));
  INV_X1    g072(.A(G183gat), .ZN(new_n274));
  INV_X1    g073(.A(G190gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n270), .A2(KEYINPUT64), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n271), .A2(new_n273), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT23), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n279), .A2(G176gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n281), .A2(G169gat), .ZN(new_n282));
  INV_X1    g081(.A(G169gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(KEYINPUT65), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n280), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  OR2_X1    g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n279), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n278), .A2(new_n285), .A3(new_n286), .A4(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT25), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT66), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n289), .A2(KEYINPUT66), .A3(new_n290), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n269), .A2(KEYINPUT68), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT24), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n269), .A2(KEYINPUT68), .A3(new_n270), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n296), .A2(new_n276), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n290), .B1(new_n280), .B2(new_n283), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n286), .B(KEYINPUT67), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n298), .A2(new_n288), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n293), .A2(new_n294), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT69), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n293), .A2(new_n304), .A3(new_n294), .A4(new_n301), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n275), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(KEYINPUT70), .A2(KEYINPUT28), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI221_X1 g110(.A(new_n275), .B1(KEYINPUT70), .B2(KEYINPUT28), .C1(new_n307), .C2(new_n308), .ZN(new_n312));
  NAND2_X1  g111(.A1(KEYINPUT70), .A2(KEYINPUT28), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(new_n286), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT71), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n315), .A2(new_n318), .A3(new_n286), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n317), .B(new_n319), .C1(KEYINPUT26), .C2(new_n287), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n314), .A2(new_n320), .A3(new_n269), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT72), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n314), .A2(new_n320), .A3(new_n323), .A4(new_n269), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n268), .B1(new_n306), .B2(new_n326), .ZN(new_n327));
  AOI211_X1 g126(.A(new_n267), .B(new_n325), .C1(new_n303), .C2(new_n305), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G227gat), .ZN(new_n330));
  INV_X1    g129(.A(G233gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT34), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT34), .ZN(new_n334));
  INV_X1    g133(.A(new_n332), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n334), .B(new_n335), .C1(new_n327), .C2(new_n328), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT33), .B1(new_n329), .B2(new_n332), .ZN(new_n337));
  XNOR2_X1  g136(.A(G15gat), .B(G43gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(G71gat), .B(G99gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n333), .B(new_n336), .C1(new_n337), .C2(new_n340), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n289), .A2(KEYINPUT66), .A3(new_n290), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT66), .B1(new_n289), .B2(new_n290), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n304), .B1(new_n344), .B2(new_n301), .ZN(new_n345));
  INV_X1    g144(.A(new_n305), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n326), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n267), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n325), .B1(new_n303), .B2(new_n305), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n268), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n332), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT33), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n340), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n350), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n334), .B1(new_n354), .B2(new_n335), .ZN(new_n355));
  INV_X1    g154(.A(new_n336), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n351), .A2(KEYINPUT32), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G141gat), .B(G148gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362));
  NOR2_X1   g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT2), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n361), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n362), .B1(new_n361), .B2(KEYINPUT2), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n363), .A2(KEYINPUT79), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(G155gat), .B2(G162gat), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT80), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n362), .ZN(new_n373));
  INV_X1    g172(.A(G148gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G141gat), .ZN(new_n375));
  INV_X1    g174(.A(G141gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G148gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n373), .B1(new_n378), .B2(new_n364), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n368), .A2(new_n370), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n366), .B1(new_n372), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT29), .ZN(new_n384));
  XOR2_X1   g183(.A(G211gat), .B(G218gat), .Z(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G211gat), .A2(G218gat), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT74), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n387), .B1(new_n388), .B2(KEYINPUT22), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT22), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n390), .A2(KEYINPUT74), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT75), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n390), .A2(KEYINPUT74), .B1(G211gat), .B2(G218gat), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT75), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n388), .A2(KEYINPUT22), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  XOR2_X1   g196(.A(G197gat), .B(G204gat), .Z(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n386), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  AOI211_X1 g199(.A(new_n385), .B(new_n398), .C1(new_n392), .C2(new_n396), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n384), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n383), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n383), .A2(new_n403), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT77), .B(KEYINPUT29), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n400), .A2(new_n401), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n406), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n404), .B2(new_n405), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n366), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n367), .A2(new_n371), .A3(KEYINPUT80), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n380), .B1(new_n379), .B2(new_n381), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n390), .A2(KEYINPUT74), .ZN(new_n422));
  AND4_X1   g221(.A1(new_n394), .A2(new_n395), .A3(new_n422), .A4(new_n387), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n394), .B1(new_n393), .B2(new_n395), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n399), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n385), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n397), .A2(new_n386), .A3(new_n399), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n408), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n403), .B1(new_n428), .B2(KEYINPUT84), .ZN(new_n429));
  OAI211_X1 g228(.A(KEYINPUT84), .B(new_n409), .C1(new_n400), .C2(new_n401), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n421), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT85), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n409), .B1(new_n400), .B2(new_n401), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT84), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n437), .A2(new_n403), .A3(new_n430), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(KEYINPUT85), .A3(new_n421), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n434), .A2(new_n412), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n417), .B1(new_n440), .B2(new_n414), .ZN(new_n441));
  INV_X1    g240(.A(G22gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(KEYINPUT88), .A3(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(G78gat), .B(G106gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT31), .B(G50gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT88), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n447), .B1(new_n441), .B2(new_n442), .ZN(new_n448));
  AOI211_X1 g247(.A(G22gat), .B(new_n417), .C1(new_n440), .C2(new_n414), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n443), .B(new_n446), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT3), .B1(new_n435), .B2(new_n436), .ZN(new_n452));
  AOI211_X1 g251(.A(new_n433), .B(new_n383), .C1(new_n452), .C2(new_n430), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT85), .B1(new_n438), .B2(new_n421), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n415), .B1(new_n455), .B2(new_n412), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n451), .B(G22gat), .C1(new_n456), .C2(new_n417), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT87), .B1(new_n441), .B2(new_n442), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n442), .ZN(new_n459));
  INV_X1    g258(.A(new_n446), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n359), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n341), .A2(new_n357), .A3(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n360), .A2(new_n450), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n267), .B(new_n418), .C1(new_n419), .C2(new_n420), .ZN(new_n465));
  NAND2_X1  g264(.A1(G225gat), .A2(G233gat), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(KEYINPUT4), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT4), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n383), .A2(new_n468), .A3(new_n267), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n421), .A2(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(new_n407), .A3(new_n268), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n466), .ZN(new_n474));
  INV_X1    g273(.A(new_n465), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n383), .A2(new_n267), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n473), .A2(KEYINPUT5), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n469), .A2(KEYINPUT81), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT81), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n383), .A2(new_n480), .A3(new_n468), .A4(new_n267), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n465), .A2(KEYINPUT4), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n474), .A2(KEYINPUT5), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n472), .ZN(new_n485));
  XNOR2_X1  g284(.A(G1gat), .B(G29gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(new_n211), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT0), .B(G57gat), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n487), .B(new_n488), .Z(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n478), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT82), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n485), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n489), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n491), .A2(KEYINPUT82), .A3(new_n492), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT83), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n496), .A2(KEYINPUT6), .A3(new_n489), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n495), .A2(KEYINPUT83), .A3(new_n497), .A4(new_n498), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G8gat), .B(G36gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(G64gat), .B(G92gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n411), .ZN(new_n508));
  NAND2_X1  g307(.A1(G226gat), .A2(G233gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT76), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(new_n349), .B2(new_n408), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n302), .A2(new_n321), .ZN(new_n512));
  INV_X1    g311(.A(new_n509), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n508), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n510), .B1(new_n306), .B2(new_n326), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n513), .B1(new_n512), .B2(new_n384), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n516), .A2(new_n411), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n507), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT78), .ZN(new_n520));
  INV_X1    g319(.A(new_n517), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n521), .B(new_n508), .C1(new_n349), .C2(new_n510), .ZN(new_n522));
  INV_X1    g321(.A(new_n507), .ZN(new_n523));
  INV_X1    g322(.A(new_n514), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n347), .A2(new_n409), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n524), .B1(new_n525), .B2(new_n510), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n522), .B(new_n523), .C1(new_n526), .C2(new_n508), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT78), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n530), .B(new_n507), .C1(new_n515), .C2(new_n518), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n511), .A2(new_n514), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n411), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n533), .A2(KEYINPUT30), .A3(new_n522), .A4(new_n523), .ZN(new_n534));
  AND4_X1   g333(.A1(new_n520), .A2(new_n529), .A3(new_n531), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n504), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT35), .B1(new_n464), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n450), .A2(new_n461), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n341), .A2(new_n357), .A3(new_n462), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n462), .B1(new_n341), .B2(new_n357), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n491), .A2(new_n492), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT89), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n543), .B1(new_n496), .B2(new_n489), .ZN(new_n544));
  AOI211_X1 g343(.A(KEYINPUT89), .B(new_n490), .C1(new_n478), .C2(new_n485), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT90), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n542), .B(KEYINPUT90), .C1(new_n544), .C2(new_n545), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(new_n502), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT35), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n535), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n541), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n536), .A2(new_n538), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT36), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n556), .B1(new_n539), .B2(new_n540), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n360), .A2(KEYINPUT36), .A3(new_n463), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT37), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n533), .A2(new_n560), .A3(new_n522), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT37), .B1(new_n515), .B2(new_n518), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(new_n562), .A3(new_n507), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT38), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n527), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n515), .A2(new_n518), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n523), .B1(new_n566), .B2(new_n560), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT38), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n521), .B(new_n411), .C1(new_n349), .C2(new_n510), .ZN(new_n569));
  OAI211_X1 g368(.A(KEYINPUT37), .B(new_n569), .C1(new_n526), .C2(new_n411), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NOR3_X1   g371(.A1(new_n565), .A2(new_n572), .A3(new_n550), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n450), .A2(new_n461), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n529), .A2(new_n520), .A3(new_n531), .A4(new_n534), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n544), .A2(new_n545), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n466), .B1(new_n483), .B2(new_n472), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT39), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n489), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR3_X1   g378(.A1(new_n475), .A2(new_n476), .A3(new_n474), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n581), .B2(new_n578), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT40), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n575), .A2(new_n576), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n574), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n555), .B(new_n559), .C1(new_n573), .C2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n259), .B1(new_n554), .B2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G113gat), .B(G141gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(G197gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT11), .B(G169gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(KEYINPUT91), .B(KEYINPUT12), .Z(new_n592));
  XOR2_X1   g391(.A(new_n591), .B(new_n592), .Z(new_n593));
  INV_X1    g392(.A(G15gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n442), .ZN(new_n595));
  INV_X1    g394(.A(G1gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(G15gat), .A2(G22gat), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n595), .A2(new_n597), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT93), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT16), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n600), .B1(new_n601), .B2(G1gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n596), .A2(KEYINPUT93), .A3(KEYINPUT16), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n598), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(G8gat), .B1(new_n598), .B2(KEYINPUT94), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI221_X1 g406(.A(new_n598), .B1(KEYINPUT94), .B2(G8gat), .C1(new_n599), .C2(new_n604), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G29gat), .A2(G36gat), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NOR3_X1   g411(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(G43gat), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(G50gat), .ZN(new_n616));
  INV_X1    g415(.A(G50gat), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(G43gat), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n614), .A2(KEYINPUT15), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT14), .ZN(new_n621));
  INV_X1    g420(.A(G29gat), .ZN(new_n622));
  INV_X1    g421(.A(G36gat), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AOI22_X1  g423(.A1(new_n624), .A2(new_n611), .B1(G29gat), .B2(G36gat), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT15), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n616), .B2(new_n618), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n617), .A2(G43gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n615), .A2(G50gat), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(new_n629), .A3(KEYINPUT15), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n625), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n620), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n609), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n620), .A2(new_n631), .A3(KEYINPUT17), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT95), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT95), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n620), .A2(new_n631), .A3(new_n636), .A4(KEYINPUT17), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n631), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT17), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n639), .A2(new_n640), .B1(new_n607), .B2(new_n608), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n633), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G229gat), .A2(G233gat), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n642), .A2(KEYINPUT18), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT18), .B1(new_n642), .B2(new_n643), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n643), .B(KEYINPUT13), .ZN(new_n646));
  INV_X1    g445(.A(new_n633), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n609), .A2(new_n632), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n644), .A2(new_n645), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT92), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n593), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n645), .ZN(new_n653));
  INV_X1    g452(.A(new_n649), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n642), .A2(KEYINPUT18), .A3(new_n643), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n593), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(KEYINPUT92), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G127gat), .B(G155gat), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n660), .B(KEYINPUT20), .Z(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n234), .A2(KEYINPUT21), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(new_n274), .A3(new_n609), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n274), .B1(new_n663), .B2(new_n609), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n667));
  OAI22_X1  g466(.A1(new_n665), .A2(new_n666), .B1(new_n234), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n666), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n234), .A2(new_n667), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n664), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n662), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G211gat), .ZN(new_n675));
  NAND2_X1  g474(.A1(G231gat), .A2(G233gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(new_n677));
  NAND3_X1  g476(.A1(new_n668), .A2(new_n671), .A3(new_n662), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n673), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n677), .ZN(new_n680));
  INV_X1    g479(.A(new_n678), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n680), .B1(new_n681), .B2(new_n672), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n227), .A2(new_n240), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n639), .A2(new_n640), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n638), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT100), .ZN(new_n688));
  NAND3_X1  g487(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n227), .A2(new_n639), .A3(new_n240), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n685), .A2(new_n638), .A3(new_n691), .A4(new_n686), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n688), .A2(new_n689), .A3(new_n690), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(G134gat), .B(G162gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(G190gat), .B(G218gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n693), .A2(new_n699), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n684), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n587), .A2(new_n659), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n504), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n504), .A2(new_n707), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(new_n596), .ZN(G1324gat));
  INV_X1    g511(.A(new_n706), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT42), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(KEYINPUT105), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT16), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n713), .A2(new_n575), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(G8gat), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n713), .A2(new_n575), .ZN(new_n720));
  AOI21_X1  g519(.A(G8gat), .B1(new_n720), .B2(new_n714), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n719), .B1(new_n721), .B2(new_n717), .ZN(G1325gat));
  NOR3_X1   g521(.A1(new_n706), .A2(new_n594), .A3(new_n559), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n539), .A2(new_n540), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n713), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n723), .B1(new_n725), .B2(new_n594), .ZN(G1326gat));
  OR3_X1    g525(.A1(new_n706), .A2(KEYINPUT106), .A3(new_n574), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT106), .B1(new_n706), .B2(new_n574), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(KEYINPUT43), .B(G22gat), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(G1327gat));
  AOI21_X1  g533(.A(new_n703), .B1(new_n554), .B2(new_n586), .ZN(new_n735));
  INV_X1    g534(.A(new_n659), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n736), .A2(new_n259), .A3(new_n683), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n708), .A2(new_n709), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(new_n622), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT45), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n554), .A2(new_n586), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n743), .B2(new_n704), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n701), .B2(new_n702), .ZN(new_n746));
  INV_X1    g545(.A(new_n702), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(KEYINPUT107), .A3(new_n700), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  AOI211_X1 g548(.A(KEYINPUT44), .B(new_n749), .C1(new_n554), .C2(new_n586), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n739), .B(new_n737), .C1(new_n744), .C2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n504), .A2(new_n535), .B1(new_n450), .B2(new_n461), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n574), .A2(new_n584), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n548), .A2(new_n549), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n563), .A2(KEYINPUT38), .B1(new_n566), .B2(new_n523), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n756), .A2(new_n502), .A3(new_n757), .A4(new_n571), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n754), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n759), .A2(new_n559), .B1(new_n537), .B2(new_n553), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT44), .B1(new_n760), .B2(new_n703), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n746), .A2(new_n748), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n743), .A2(new_n742), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n764), .A2(KEYINPUT108), .A3(new_n739), .A4(new_n737), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n753), .A2(new_n765), .A3(G29gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n741), .A2(new_n766), .ZN(G1328gat));
  NAND3_X1  g566(.A1(new_n764), .A2(new_n575), .A3(new_n737), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G36gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n738), .A2(new_n623), .A3(new_n575), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT46), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(KEYINPUT109), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n771), .A2(KEYINPUT109), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n769), .B(new_n774), .C1(new_n772), .C2(new_n770), .ZN(G1329gat));
  NOR2_X1   g574(.A1(new_n559), .A2(new_n615), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n764), .A2(new_n737), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n738), .A2(new_n724), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n615), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT47), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT47), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n777), .A2(new_n779), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(G1330gat));
  INV_X1    g583(.A(KEYINPUT48), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n785), .A2(KEYINPUT110), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n735), .A2(new_n617), .A3(new_n538), .A4(new_n737), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(KEYINPUT110), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n538), .B(new_n737), .C1(new_n744), .C2(new_n750), .ZN(new_n790));
  AOI211_X1 g589(.A(new_n786), .B(new_n789), .C1(new_n790), .C2(G50gat), .ZN(new_n791));
  INV_X1    g590(.A(new_n786), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(G50gat), .ZN(new_n793));
  INV_X1    g592(.A(new_n789), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n791), .A2(new_n795), .ZN(G1331gat));
  INV_X1    g595(.A(new_n259), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n683), .A2(new_n703), .A3(new_n658), .A4(new_n652), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n760), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n739), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g602(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n799), .A2(new_n575), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT112), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n799), .A2(new_n807), .A3(new_n575), .A4(new_n804), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT49), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n228), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n806), .A2(new_n810), .A3(new_n228), .A4(new_n808), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(G1333gat));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n724), .ZN(new_n815));
  INV_X1    g614(.A(G71gat), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n559), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n799), .A2(G71gat), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT50), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n817), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(G1334gat));
  NAND2_X1  g623(.A1(new_n799), .A2(new_n538), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g625(.A1(new_n659), .A2(new_n683), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n797), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(new_n761), .B2(new_n763), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n236), .B1(new_n832), .B2(new_n710), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n735), .A2(KEYINPUT51), .A3(new_n827), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT51), .B1(new_n735), .B2(new_n827), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n259), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n739), .B1(new_n210), .B2(new_n212), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n833), .B1(new_n837), .B2(new_n838), .ZN(G1336gat));
  OAI211_X1 g638(.A(new_n575), .B(new_n829), .C1(new_n744), .C2(new_n750), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G92gat), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n535), .A2(G92gat), .A3(new_n797), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n842), .B1(new_n835), .B2(new_n836), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT51), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n743), .A2(new_n704), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n828), .ZN(new_n848));
  AOI22_X1  g647(.A1(new_n848), .A2(new_n834), .B1(KEYINPUT113), .B2(new_n842), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n842), .A2(KEYINPUT113), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n849), .A2(new_n850), .B1(G92gat), .B2(new_n840), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n845), .B1(new_n851), .B2(new_n844), .ZN(G1337gat));
  XNOR2_X1  g651(.A(KEYINPUT114), .B(G99gat), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n853), .B1(new_n832), .B2(new_n559), .ZN(new_n854));
  OR3_X1    g653(.A1(new_n539), .A2(new_n540), .A3(new_n853), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n854), .B1(new_n837), .B2(new_n855), .ZN(G1338gat));
  AOI21_X1  g655(.A(new_n215), .B1(new_n831), .B2(new_n538), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n538), .A2(new_n215), .A3(new_n259), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT115), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n860), .B1(new_n848), .B2(new_n834), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT53), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n861), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n538), .B(new_n829), .C1(new_n744), .C2(new_n750), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(G106gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n862), .A2(new_n867), .ZN(G1339gat));
  INV_X1    g667(.A(G113gat), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n705), .A2(KEYINPUT116), .A3(new_n736), .A4(new_n797), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n871), .B1(new_n798), .B2(new_n259), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  OR3_X1    g672(.A1(new_n249), .A2(new_n250), .A3(new_n255), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n247), .A2(new_n248), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n203), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n247), .A2(new_n204), .A3(new_n248), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(KEYINPUT54), .A3(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n256), .B1(new_n249), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(KEYINPUT55), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n878), .A2(new_n880), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT55), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n659), .A2(new_n874), .A3(new_n881), .A4(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n647), .A2(new_n648), .A3(new_n646), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n886), .B1(new_n642), .B2(new_n643), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n650), .A2(new_n593), .B1(new_n591), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n259), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n762), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n884), .A2(new_n874), .A3(new_n881), .A4(new_n888), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n749), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n684), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n464), .B1(new_n873), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n739), .A3(new_n535), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n896), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n869), .B1(new_n899), .B2(new_n659), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n801), .A2(new_n535), .A3(new_n894), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n901), .A2(G113gat), .A3(new_n736), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n900), .A2(new_n902), .ZN(G1340gat));
  OR3_X1    g702(.A1(new_n901), .A2(G120gat), .A3(new_n797), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n897), .A2(new_n259), .A3(new_n898), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G120gat), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT118), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n904), .A2(new_n909), .A3(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1341gat));
  NAND3_X1  g710(.A1(new_n899), .A2(G127gat), .A3(new_n683), .ZN(new_n912));
  INV_X1    g711(.A(G127gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n913), .B1(new_n901), .B2(new_n684), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n912), .A2(new_n914), .ZN(G1342gat));
  NOR3_X1   g714(.A1(new_n901), .A2(G134gat), .A3(new_n703), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT56), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n899), .A2(new_n704), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n918), .A2(KEYINPUT119), .A3(G134gat), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT119), .B1(new_n918), .B2(G134gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(G1343gat));
  AOI21_X1  g720(.A(new_n574), .B1(new_n873), .B2(new_n893), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n575), .B1(new_n557), .B2(new_n558), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n801), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n924), .A2(G141gat), .A3(new_n736), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n925), .A2(KEYINPUT58), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT57), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n889), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n259), .A2(new_n888), .A3(KEYINPUT120), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n885), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n892), .B1(new_n931), .B2(new_n703), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT121), .B1(new_n932), .B2(new_n683), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n259), .A2(KEYINPUT120), .A3(new_n888), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT120), .B1(new_n259), .B2(new_n888), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n704), .B1(new_n937), .B2(new_n885), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n934), .B(new_n684), .C1(new_n938), .C2(new_n892), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n933), .A2(new_n939), .A3(new_n873), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n927), .B1(new_n940), .B2(new_n538), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n885), .A2(new_n889), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n749), .ZN(new_n943));
  INV_X1    g742(.A(new_n892), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n683), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n870), .A2(new_n872), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n927), .B(new_n538), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n923), .A3(new_n739), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n941), .A2(new_n736), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n926), .B1(new_n376), .B2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT58), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT122), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n940), .A2(new_n538), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT57), .ZN(new_n954));
  INV_X1    g753(.A(new_n948), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n941), .A2(KEYINPUT122), .A3(new_n948), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n659), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n925), .B1(new_n958), .B2(G141gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n950), .B1(new_n951), .B2(new_n959), .ZN(G1344gat));
  INV_X1    g759(.A(new_n924), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(new_n374), .A3(new_n259), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT59), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n922), .A2(KEYINPUT57), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n964), .A2(KEYINPUT123), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(KEYINPUT123), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n891), .A2(new_n703), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n684), .B1(new_n938), .B2(new_n967), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n798), .A2(new_n259), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n574), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n965), .B(new_n966), .C1(KEYINPUT57), .C2(new_n970), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n971), .A2(new_n739), .A3(new_n259), .A4(new_n923), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n963), .B1(new_n972), .B2(G148gat), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n954), .A2(new_n952), .A3(new_n955), .ZN(new_n974));
  OAI21_X1  g773(.A(KEYINPUT122), .B1(new_n941), .B2(new_n948), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n797), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n976), .A2(KEYINPUT59), .A3(new_n374), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n962), .B1(new_n973), .B2(new_n977), .ZN(G1345gat));
  AOI21_X1  g777(.A(G155gat), .B1(new_n961), .B2(new_n683), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n684), .B1(new_n974), .B2(new_n975), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n979), .B1(G155gat), .B2(new_n980), .ZN(G1346gat));
  OAI21_X1  g780(.A(new_n762), .B1(new_n956), .B2(new_n957), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(KEYINPUT124), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n984), .B(new_n762), .C1(new_n956), .C2(new_n957), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n983), .A2(G162gat), .A3(new_n985), .ZN(new_n986));
  OR3_X1    g785(.A1(new_n924), .A2(G162gat), .A3(new_n703), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(G1347gat));
  XNOR2_X1  g787(.A(new_n739), .B(KEYINPUT111), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n989), .A2(new_n575), .A3(new_n894), .ZN(new_n990));
  OAI21_X1  g789(.A(G169gat), .B1(new_n990), .B2(new_n736), .ZN(new_n991));
  OAI211_X1 g790(.A(new_n709), .B(new_n708), .C1(new_n945), .C2(new_n946), .ZN(new_n992));
  NOR3_X1   g791(.A1(new_n992), .A2(new_n464), .A3(new_n535), .ZN(new_n993));
  OAI211_X1 g792(.A(new_n993), .B(new_n659), .C1(new_n282), .C2(new_n284), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n991), .A2(new_n994), .ZN(G1348gat));
  AOI21_X1  g794(.A(G176gat), .B1(new_n993), .B2(new_n259), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n990), .A2(new_n797), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n996), .B1(new_n997), .B2(G176gat), .ZN(G1349gat));
  OAI21_X1  g797(.A(G183gat), .B1(new_n990), .B2(new_n684), .ZN(new_n999));
  OAI211_X1 g798(.A(new_n993), .B(new_n683), .C1(new_n308), .C2(new_n307), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g800(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n1002));
  XNOR2_X1  g801(.A(new_n1001), .B(new_n1002), .ZN(G1350gat));
  OAI21_X1  g802(.A(G190gat), .B1(new_n990), .B2(new_n703), .ZN(new_n1004));
  XNOR2_X1  g803(.A(new_n1004), .B(KEYINPUT61), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n993), .A2(new_n275), .A3(new_n762), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1005), .A2(new_n1006), .ZN(G1351gat));
  NOR3_X1   g806(.A1(new_n801), .A2(new_n535), .A3(new_n818), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n971), .A2(new_n659), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g810(.A1(new_n971), .A2(KEYINPUT126), .A3(new_n659), .A4(new_n1008), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n1011), .A2(G197gat), .A3(new_n1012), .ZN(new_n1013));
  OR4_X1    g812(.A1(new_n574), .A2(new_n992), .A3(new_n535), .A4(new_n818), .ZN(new_n1014));
  OR3_X1    g813(.A1(new_n1014), .A2(G197gat), .A3(new_n736), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1013), .A2(new_n1015), .ZN(G1352gat));
  XNOR2_X1  g815(.A(KEYINPUT127), .B(G204gat), .ZN(new_n1017));
  NOR3_X1   g816(.A1(new_n1014), .A2(new_n797), .A3(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1018), .B(KEYINPUT62), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n971), .A2(new_n259), .A3(new_n1008), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1020), .A2(new_n1017), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1019), .A2(new_n1021), .ZN(G1353gat));
  OR3_X1    g821(.A1(new_n1014), .A2(G211gat), .A3(new_n684), .ZN(new_n1023));
  NAND3_X1  g822(.A1(new_n971), .A2(new_n683), .A3(new_n1008), .ZN(new_n1024));
  AND3_X1   g823(.A1(new_n1024), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1025));
  AOI21_X1  g824(.A(KEYINPUT63), .B1(new_n1024), .B2(G211gat), .ZN(new_n1026));
  OAI21_X1  g825(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(G1354gat));
  AND2_X1   g826(.A1(new_n971), .A2(new_n1008), .ZN(new_n1028));
  INV_X1    g827(.A(G218gat), .ZN(new_n1029));
  NOR2_X1   g828(.A1(new_n703), .A2(new_n1029), .ZN(new_n1030));
  OR2_X1    g829(.A1(new_n1014), .A2(new_n749), .ZN(new_n1031));
  AOI22_X1  g830(.A1(new_n1028), .A2(new_n1030), .B1(new_n1031), .B2(new_n1029), .ZN(G1355gat));
endmodule


