//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n634, new_n635, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1208, new_n1209,
    new_n1210, new_n1211;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  AND2_X1   g017(.A1(G2072), .A2(G2078), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G101), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n462), .ZN(new_n473));
  NAND3_X1  g048(.A1(KEYINPUT68), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n471), .B1(new_n475), .B2(G137), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n467), .A2(new_n476), .ZN(G160));
  AND3_X1   g052(.A1(KEYINPUT68), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(KEYINPUT3), .B1(KEYINPUT68), .B2(G2104), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n468), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G136), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n468), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  OAI22_X1  g058(.A1(new_n480), .A2(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n485));
  OAI21_X1  g060(.A(G2105), .B1(new_n478), .B2(new_n479), .ZN(new_n486));
  INV_X1    g061(.A(G124), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n489), .A2(KEYINPUT69), .A3(G124), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n484), .B1(new_n488), .B2(new_n490), .ZN(G162));
  OAI211_X1 g066(.A(G138), .B(new_n468), .C1(new_n478), .C2(new_n479), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT3), .B(G2104), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n494), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n492), .A2(KEYINPUT4), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n468), .A2(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  OAI22_X1  g074(.A1(new_n486), .A2(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n496), .A2(new_n500), .ZN(G164));
  OR2_X1    g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(new_n506), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n504), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n513), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n507), .A2(new_n517), .ZN(G166));
  NAND2_X1  g093(.A1(new_n515), .A2(G89), .ZN(new_n519));
  NAND2_X1  g094(.A1(G63), .A2(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(new_n504), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT70), .B(G51), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n512), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n525), .B(new_n526), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n522), .A2(new_n524), .A3(new_n527), .ZN(G168));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n502), .A2(new_n503), .ZN(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n532), .A2(KEYINPUT72), .A3(G651), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n535), .B2(new_n506), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n512), .A2(G52), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n504), .A2(new_n515), .A3(G90), .ZN(new_n539));
  AOI21_X1  g114(.A(KEYINPUT73), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n539), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n537), .B1(new_n540), .B2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n546), .B1(new_n502), .B2(new_n503), .ZN(new_n547));
  AND2_X1   g122(.A1(G68), .A2(G543), .ZN(new_n548));
  OAI21_X1  g123(.A(G651), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n512), .A2(G43), .ZN(new_n550));
  XOR2_X1   g125(.A(KEYINPUT74), .B(G81), .Z(new_n551));
  NAND3_X1  g126(.A1(new_n551), .A2(new_n504), .A3(new_n515), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(KEYINPUT75), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n549), .A2(new_n555), .A3(new_n552), .A4(new_n550), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(G188));
  AOI22_X1  g139(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n565), .A2(new_n506), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n567));
  INV_X1    g142(.A(new_n511), .ZN(new_n568));
  NOR2_X1   g143(.A1(KEYINPUT6), .A2(G651), .ZN(new_n569));
  OAI211_X1 g144(.A(G53), .B(G543), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n567), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR3_X1   g148(.A1(new_n570), .A2(KEYINPUT77), .A3(KEYINPUT9), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT76), .B1(new_n571), .B2(new_n572), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n570), .A2(new_n577), .A3(KEYINPUT9), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n566), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n516), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n504), .A2(new_n515), .A3(KEYINPUT78), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n582), .A2(G91), .A3(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n582), .A2(KEYINPUT79), .A3(G91), .A4(new_n583), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n580), .A2(new_n588), .ZN(G299));
  NAND3_X1  g164(.A1(new_n522), .A2(new_n524), .A3(new_n527), .ZN(G286));
  INV_X1    g165(.A(G166), .ZN(G303));
  NAND2_X1  g166(.A1(new_n512), .A2(G49), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n582), .A2(G87), .A3(new_n583), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G288));
  NAND3_X1  g172(.A1(new_n515), .A2(G48), .A3(G543), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G73), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G61), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n530), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n599), .B1(new_n604), .B2(G651), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n582), .A2(G86), .A3(new_n583), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(G305));
  INV_X1    g182(.A(new_n516), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G85), .B1(G47), .B2(new_n512), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n506), .B2(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  XNOR2_X1  g187(.A(KEYINPUT82), .B(G66), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n504), .A2(new_n613), .B1(G79), .B2(G543), .ZN(new_n614));
  INV_X1    g189(.A(new_n512), .ZN(new_n615));
  INV_X1    g190(.A(G54), .ZN(new_n616));
  OAI22_X1  g191(.A1(new_n614), .A2(new_n506), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI221_X1 g194(.A(KEYINPUT83), .B1(new_n615), .B2(new_n616), .C1(new_n614), .C2(new_n506), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n582), .A2(G92), .A3(new_n583), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT10), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g199(.A1(new_n582), .A2(KEYINPUT10), .A3(G92), .A4(new_n583), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(KEYINPUT84), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT84), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n621), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  AND2_X1   g205(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n612), .B1(new_n631), .B2(G868), .ZN(G284));
  XNOR2_X1  g207(.A(G284), .B(KEYINPUT85), .ZN(G321));
  INV_X1    g208(.A(G868), .ZN(new_n634));
  NAND2_X1  g209(.A1(G299), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(new_n634), .B2(G168), .ZN(G297));
  OAI21_X1  g211(.A(new_n635), .B1(new_n634), .B2(G168), .ZN(G280));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n631), .B1(new_n638), .B2(G860), .ZN(G148));
  NAND3_X1  g214(.A1(new_n628), .A2(new_n630), .A3(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(KEYINPUT86), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n640), .A2(KEYINPUT86), .ZN(new_n643));
  OAI21_X1  g218(.A(G868), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g220(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g221(.A1(new_n489), .A2(G123), .ZN(new_n647));
  OR2_X1    g222(.A1(G99), .A2(G2105), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n648), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(G135), .B2(new_n475), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2096), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n468), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT12), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT13), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2100), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n656), .ZN(G156));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT87), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2427), .B(G2430), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(KEYINPUT14), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2451), .B(G2454), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT16), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n666), .B(new_n667), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n664), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2443), .B(G2446), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(G14), .B1(new_n669), .B2(new_n671), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(G401));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  XNOR2_X1  g250(.A(G2072), .B(G2078), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT18), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n676), .B(KEYINPUT17), .Z(new_n680));
  INV_X1    g255(.A(new_n675), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n681), .A2(new_n677), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n679), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n677), .B1(new_n676), .B2(KEYINPUT88), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(KEYINPUT88), .B2(new_n676), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n685), .A2(KEYINPUT89), .A3(new_n681), .ZN(new_n686));
  INV_X1    g261(.A(new_n677), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(new_n680), .ZN(new_n688));
  AOI21_X1  g263(.A(KEYINPUT89), .B1(new_n685), .B2(new_n681), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n683), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G2096), .B(G2100), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(G227));
  XNOR2_X1  g267(.A(G1971), .B(G1976), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT19), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT90), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1961), .B(G1966), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n695), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT20), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n695), .B1(new_n697), .B2(new_n699), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n697), .A2(new_n699), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n701), .B(new_n704), .C1(new_n694), .C2(new_n703), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT91), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n705), .B(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(G1991), .B(G1996), .Z(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(new_n710), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(G1981), .B(G1986), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n711), .A2(new_n714), .A3(new_n712), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(G229));
  INV_X1    g293(.A(KEYINPUT93), .ZN(new_n719));
  NAND2_X1  g294(.A1(G305), .A2(G16), .ZN(new_n720));
  INV_X1    g295(.A(G6), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(G16), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n719), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  AOI211_X1 g299(.A(KEYINPUT93), .B(new_n722), .C1(G305), .C2(G16), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT32), .B(G1981), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n727), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n724), .B2(new_n725), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n732), .A2(G23), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G288), .B2(G16), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT33), .B(G1976), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G16), .A2(G22), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G166), .B2(G16), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT94), .B(G1971), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n734), .A2(new_n735), .ZN(new_n741));
  NOR3_X1   g316(.A1(new_n736), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n731), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT34), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n731), .A2(new_n742), .A3(KEYINPUT34), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n489), .A2(G119), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n475), .A2(G131), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n468), .A2(G107), .ZN(new_n750));
  OAI21_X1  g325(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n748), .B(new_n749), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT92), .ZN(new_n753));
  MUX2_X1   g328(.A(G25), .B(new_n753), .S(G29), .Z(new_n754));
  XOR2_X1   g329(.A(KEYINPUT35), .B(G1991), .Z(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n754), .B(new_n756), .ZN(new_n757));
  MUX2_X1   g332(.A(G24), .B(G290), .S(G16), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1986), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n747), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(KEYINPUT95), .A2(KEYINPUT36), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT96), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n763), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n747), .A2(new_n760), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n732), .A2(G4), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n631), .B2(new_n732), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT97), .B(G1348), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(G29), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n772), .A2(G33), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT25), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G139), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(new_n480), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT100), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n493), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n782));
  OAI22_X1  g357(.A1(new_n780), .A2(new_n781), .B1(new_n468), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n773), .B1(new_n783), .B2(G29), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n784), .A2(G2072), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(G2072), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n772), .A2(G32), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT103), .B(KEYINPUT26), .Z(new_n789));
  NAND3_X1  g364(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n489), .A2(G129), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n793));
  AND3_X1   g368(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n475), .A2(G141), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT102), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n788), .B1(new_n798), .B2(new_n772), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT27), .B(G1996), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(G301), .A2(G16), .ZN(new_n803));
  INV_X1    g378(.A(G1961), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n732), .A2(G5), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT99), .B(KEYINPUT28), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n772), .A2(G26), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n489), .A2(G128), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n475), .A2(G140), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n468), .A2(G116), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n809), .B1(new_n814), .B2(G29), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G2067), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n802), .A2(new_n806), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(G27), .A2(G29), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G164), .B2(G29), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(G2078), .Z(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT101), .B(KEYINPUT24), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G34), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(G29), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G160), .B2(G29), .ZN(new_n824));
  INV_X1    g399(.A(G2084), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n820), .B(new_n826), .C1(new_n799), .C2(new_n801), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n772), .A2(G35), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G162), .B2(new_n772), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT29), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n829), .A2(KEYINPUT29), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n832), .A2(G2090), .A3(new_n833), .ZN(new_n834));
  NOR4_X1   g409(.A1(new_n787), .A2(new_n817), .A3(new_n827), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n732), .A2(G21), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G168), .B2(new_n732), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G1966), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n651), .A2(G29), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT30), .B(G28), .ZN(new_n840));
  OR2_X1    g415(.A1(KEYINPUT31), .A2(G11), .ZN(new_n841));
  NAND2_X1  g416(.A1(KEYINPUT31), .A2(G11), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n840), .A2(new_n772), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(G1966), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n845), .B(new_n836), .C1(G168), .C2(new_n732), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n838), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n804), .B1(new_n803), .B2(new_n805), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT104), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OR3_X1    g424(.A1(new_n847), .A2(new_n848), .A3(KEYINPUT104), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n557), .A2(G16), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n732), .A2(G19), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n852), .B1(new_n851), .B2(new_n853), .ZN(new_n855));
  INV_X1    g430(.A(G1341), .ZN(new_n856));
  OR3_X1    g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n856), .B1(new_n854), .B2(new_n855), .ZN(new_n858));
  AND4_X1   g433(.A1(new_n849), .A2(new_n850), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n771), .A2(new_n835), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n732), .A2(G20), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT23), .Z(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(G299), .B2(G16), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(G1956), .ZN(new_n864));
  OAI21_X1  g439(.A(G2090), .B1(new_n832), .B2(new_n833), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n864), .A2(KEYINPUT105), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(KEYINPUT105), .B1(new_n864), .B2(new_n865), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n860), .A2(new_n868), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n767), .A2(new_n869), .ZN(G311));
  INV_X1    g445(.A(KEYINPUT106), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n765), .B1(new_n747), .B2(new_n760), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n747), .A2(new_n760), .A3(new_n765), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n869), .B(new_n871), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n871), .B1(new_n767), .B2(new_n869), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(G150));
  INV_X1    g452(.A(KEYINPUT109), .ZN(new_n878));
  INV_X1    g453(.A(G860), .ZN(new_n879));
  NAND2_X1  g454(.A1(G80), .A2(G543), .ZN(new_n880));
  INV_X1    g455(.A(G67), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(new_n530), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n883), .A3(G651), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT107), .B1(new_n885), .B2(new_n506), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AOI22_X1  g462(.A1(new_n608), .A2(G93), .B1(G55), .B2(new_n512), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n557), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n552), .A2(new_n550), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n887), .A2(new_n549), .A3(new_n891), .A4(new_n888), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n631), .A2(G559), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n879), .B1(new_n898), .B2(KEYINPUT39), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(KEYINPUT39), .A3(new_n897), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(KEYINPUT108), .A3(KEYINPUT39), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n889), .A2(G860), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT37), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n878), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n906), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n903), .A2(new_n902), .ZN(new_n909));
  OAI211_X1 g484(.A(KEYINPUT109), .B(new_n908), .C1(new_n909), .C2(new_n899), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(G145));
  XNOR2_X1  g486(.A(new_n783), .B(new_n797), .ZN(new_n912));
  OAI21_X1  g487(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n913));
  INV_X1    g488(.A(G118), .ZN(new_n914));
  AOI22_X1  g489(.A1(new_n913), .A2(KEYINPUT111), .B1(new_n914), .B2(G2105), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(KEYINPUT111), .B2(new_n913), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n489), .A2(G130), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n475), .A2(G142), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  XOR2_X1   g494(.A(new_n919), .B(new_n654), .Z(new_n920));
  XNOR2_X1  g495(.A(new_n912), .B(new_n920), .ZN(new_n921));
  XOR2_X1   g496(.A(G164), .B(new_n814), .Z(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(new_n753), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n921), .B(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(G160), .B(KEYINPUT110), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n925), .B(new_n651), .Z(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(G162), .ZN(new_n927));
  AOI21_X1  g502(.A(G37), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n927), .B2(new_n924), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g505(.A1(G299), .A2(new_n627), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n580), .A2(new_n588), .A3(new_n621), .A4(new_n626), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n642), .A2(new_n643), .A3(new_n893), .ZN(new_n935));
  INV_X1    g510(.A(new_n893), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n640), .A2(KEYINPUT86), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n936), .B1(new_n937), .B2(new_n641), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n934), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n893), .B1(new_n642), .B2(new_n643), .ZN(new_n940));
  INV_X1    g515(.A(new_n932), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n580), .A2(new_n588), .B1(new_n621), .B2(new_n626), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT41), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT41), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n931), .A2(new_n944), .A3(new_n932), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n937), .A2(new_n641), .A3(new_n936), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n940), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(G288), .B(G305), .ZN(new_n949));
  XNOR2_X1  g524(.A(G303), .B(G290), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n950), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT42), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n939), .A2(new_n948), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n939), .B2(new_n948), .ZN(new_n956));
  OAI21_X1  g531(.A(G868), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n889), .A2(new_n634), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(G295));
  INV_X1    g534(.A(new_n954), .ZN(new_n960));
  INV_X1    g535(.A(new_n948), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n933), .B1(new_n940), .B2(new_n947), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n939), .A2(new_n948), .A3(new_n954), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n634), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n958), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT112), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n957), .A2(new_n968), .A3(new_n958), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(G331));
  NAND2_X1  g545(.A1(G301), .A2(G168), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n537), .B(G286), .C1(new_n540), .C2(new_n543), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n893), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n971), .A2(new_n890), .A3(new_n972), .A4(new_n892), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n946), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n933), .B1(new_n975), .B2(new_n974), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(new_n953), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G37), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n931), .A2(KEYINPUT115), .A3(new_n944), .A4(new_n932), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n982), .A2(new_n975), .A3(new_n974), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n943), .A2(new_n984), .A3(new_n945), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n978), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n980), .B(new_n981), .C1(new_n986), .C2(new_n953), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n988));
  INV_X1    g563(.A(new_n953), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n974), .A2(new_n975), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(new_n945), .B2(new_n943), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n991), .B2(new_n978), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n992), .A2(new_n981), .A3(new_n980), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n988), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n993), .A2(KEYINPUT114), .A3(KEYINPUT43), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(new_n987), .B2(KEYINPUT43), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n986), .A2(new_n953), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n978), .B1(new_n946), .B2(new_n976), .ZN(new_n1002));
  AOI21_X1  g577(.A(G37), .B1(new_n1002), .B2(new_n953), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1001), .A2(new_n1003), .A3(KEYINPUT116), .A4(new_n1004), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n997), .A2(new_n998), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(KEYINPUT113), .B(KEYINPUT44), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n994), .B1(new_n1006), .B2(new_n1007), .ZN(G397));
  NAND2_X1  g583(.A1(G286), .A2(G8), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1384), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(new_n496), .B2(new_n500), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(KEYINPUT45), .B(new_n1012), .C1(new_n496), .C2(new_n500), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n467), .A2(new_n476), .A3(G40), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n845), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1017), .B1(new_n1013), .B2(KEYINPUT50), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1022), .B(new_n1012), .C1(new_n496), .C2(new_n500), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n825), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1011), .B1(new_n1025), .B2(G8), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT124), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1013), .A2(KEYINPUT50), .ZN(new_n1028));
  AND4_X1   g603(.A1(new_n825), .A2(new_n1028), .A3(new_n1018), .A4(new_n1023), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1017), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1966), .B1(new_n1030), .B2(new_n1016), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1027), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1020), .A2(KEYINPUT124), .A3(new_n1024), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(G168), .ZN(new_n1035));
  INV_X1    g610(.A(G8), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1010), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1026), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1009), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1032), .A2(new_n1033), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT125), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT125), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1032), .A2(new_n1033), .A3(new_n1042), .A4(new_n1039), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT62), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1026), .ZN(new_n1046));
  AOI21_X1  g621(.A(G286), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1037), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1046), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT62), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1049), .A2(new_n1050), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1051));
  NAND3_X1  g626(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(G1971), .B1(new_n1030), .B2(new_n1016), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1028), .A2(new_n1018), .A3(new_n1023), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1057), .A2(G2090), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1055), .B(G8), .C1(new_n1056), .C2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(G8), .B1(new_n1058), .B2(new_n1056), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT120), .B1(new_n1064), .B2(new_n1036), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1066), .B(G8), .C1(new_n1013), .C2(new_n1017), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1976), .ZN(new_n1069));
  OR2_X1    g644(.A1(G288), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT52), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT52), .B1(G288), .B2(new_n1069), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1068), .A2(new_n1070), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1981), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n605), .A2(new_n1075), .A3(new_n606), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n600), .B(KEYINPUT81), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n603), .B1(new_n502), .B2(new_n503), .ZN(new_n1078));
  OAI21_X1  g653(.A(G651), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n504), .A2(new_n515), .A3(G86), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(new_n598), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G1981), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1076), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(KEYINPUT121), .A2(KEYINPUT49), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT49), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1083), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(new_n1068), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1072), .A2(new_n1074), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n1093));
  OR3_X1    g668(.A1(new_n1019), .A2(new_n1093), .A3(G2078), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1093), .B1(new_n1019), .B2(G2078), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1057), .A2(new_n804), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(G171), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1063), .A2(new_n1092), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1045), .A2(new_n1051), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT126), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1045), .A2(new_n1051), .A3(KEYINPUT126), .A4(new_n1099), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(G299), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G1956), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1057), .A2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT56), .B(G2072), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1030), .A2(new_n1016), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n580), .A2(new_n588), .A3(new_n1104), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1106), .A2(new_n1108), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(G2067), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1057), .A2(new_n770), .B1(new_n1113), .B2(new_n1064), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1114), .A2(new_n627), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1111), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1104), .B1(new_n580), .B2(new_n588), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1110), .ZN(new_n1119));
  AOI21_X1  g694(.A(G1956), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n1117), .A2(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1116), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1112), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1114), .A2(new_n627), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT60), .B1(new_n1126), .B2(new_n1115), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1121), .A2(new_n1112), .A3(KEYINPUT61), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n627), .A2(KEYINPUT60), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1114), .A2(new_n1130), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT58), .B(G1341), .Z(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT123), .ZN(new_n1135));
  INV_X1    g710(.A(G1996), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1030), .A2(new_n1136), .A3(new_n1016), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1132), .A2(new_n1138), .A3(new_n1133), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1135), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1140), .A2(new_n1141), .A3(new_n558), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1141), .B1(new_n1140), .B2(new_n558), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1131), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1122), .B1(new_n1129), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1049), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1094), .A2(G301), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1098), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT54), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT54), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1098), .A2(new_n1150), .A3(new_n1147), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1063), .A2(new_n1092), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1145), .A2(new_n1146), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1072), .A2(new_n1074), .A3(new_n1091), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1059), .ZN(new_n1156));
  NOR2_X1   g731(.A1(G288), .A2(G1976), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1091), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1076), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1155), .A2(new_n1156), .B1(new_n1159), .B2(new_n1068), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1060), .B(new_n1055), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT63), .ZN(new_n1162));
  AOI211_X1 g737(.A(new_n1036), .B(G286), .C1(new_n1020), .C2(new_n1024), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1161), .A2(new_n1155), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1162), .B1(new_n1153), .B2(new_n1163), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1102), .A2(new_n1103), .A3(new_n1154), .A4(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1136), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1170), .A2(new_n797), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT117), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1169), .A2(G1996), .A3(new_n797), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1173), .B(KEYINPUT118), .Z(new_n1174));
  INV_X1    g749(.A(new_n1169), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n814), .B(new_n1113), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1172), .A2(new_n1174), .A3(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n753), .B(new_n755), .ZN(new_n1179));
  OR2_X1    g754(.A1(new_n1179), .A2(KEYINPUT119), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(KEYINPUT119), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1180), .A2(new_n1169), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(G290), .B(G1986), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1183), .B1(new_n1169), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1168), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1175), .B1(new_n798), .B2(new_n1176), .ZN(new_n1187));
  OR2_X1    g762(.A1(new_n1170), .A2(KEYINPUT46), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1170), .A2(KEYINPUT46), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  XOR2_X1   g765(.A(new_n1190), .B(KEYINPUT47), .Z(new_n1191));
  NOR3_X1   g766(.A1(new_n1175), .A2(G1986), .A3(G290), .ZN(new_n1192));
  XOR2_X1   g767(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1193));
  XNOR2_X1  g768(.A(new_n1192), .B(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1191), .B1(new_n1183), .B2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n753), .A2(new_n756), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1178), .A2(new_n1196), .ZN(new_n1197));
  OR2_X1    g772(.A1(new_n814), .A2(G2067), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1175), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1186), .A2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g776(.A(G319), .B1(new_n672), .B2(new_n673), .ZN(new_n1203));
  OR2_X1    g777(.A1(new_n1203), .A2(G227), .ZN(new_n1204));
  AOI21_X1  g778(.A(new_n1204), .B1(new_n716), .B2(new_n717), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n929), .A2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g780(.A1(new_n1006), .A2(new_n1206), .ZN(G308));
  INV_X1    g781(.A(new_n998), .ZN(new_n1208));
  AOI21_X1  g782(.A(KEYINPUT114), .B1(new_n993), .B2(KEYINPUT43), .ZN(new_n1209));
  NOR2_X1   g783(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  AND2_X1   g784(.A1(new_n1000), .A2(new_n1005), .ZN(new_n1211));
  OAI211_X1 g785(.A(new_n929), .B(new_n1205), .C1(new_n1210), .C2(new_n1211), .ZN(G225));
endmodule


