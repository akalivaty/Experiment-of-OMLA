//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  INV_X1    g003(.A(G176gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT26), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n204), .A2(new_n205), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT26), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(KEYINPUT27), .B(G183gat), .Z(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT68), .ZN(new_n214));
  INV_X1    g013(.A(G183gat), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n215), .A2(KEYINPUT27), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n217));
  AOI21_X1  g016(.A(G190gat), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT28), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT28), .ZN(new_n220));
  NOR3_X1   g019(.A1(new_n213), .A2(new_n220), .A3(G190gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n203), .B(new_n212), .C1(new_n219), .C2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n210), .A2(KEYINPUT66), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(new_n208), .B2(KEYINPUT23), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n206), .B1(KEYINPUT23), .B2(new_n208), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n232), .A2(KEYINPUT65), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(KEYINPUT65), .ZN(new_n234));
  NAND3_X1  g033(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(G183gat), .B2(G190gat), .ZN(new_n236));
  OR3_X1    g035(.A1(new_n233), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n223), .B1(new_n231), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239));
  OR2_X1    g038(.A1(new_n203), .A2(KEYINPUT67), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT24), .B1(new_n203), .B2(KEYINPUT67), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n236), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NOR3_X1   g041(.A1(new_n230), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n222), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(KEYINPUT69), .B2(KEYINPUT1), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G120gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n247), .A2(KEYINPUT1), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n246), .B(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n249), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n251), .B(new_n222), .C1(new_n238), .C2(new_n243), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G227gat), .ZN(new_n254));
  INV_X1    g053(.A(G233gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n202), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT34), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT32), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n261), .B1(new_n253), .B2(new_n257), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n250), .A2(KEYINPUT70), .A3(new_n256), .A4(new_n252), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT33), .B1(new_n262), .B2(new_n263), .ZN(new_n265));
  XOR2_X1   g064(.A(G15gat), .B(G43gat), .Z(new_n266));
  XNOR2_X1  g065(.A(G71gat), .B(G99gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NOR3_X1   g068(.A1(new_n264), .A2(new_n265), .A3(new_n269), .ZN(new_n270));
  AOI221_X4 g069(.A(new_n260), .B1(KEYINPUT33), .B2(new_n268), .C1(new_n262), .C2(new_n263), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n259), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n264), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n262), .A2(new_n263), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT33), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n273), .A2(new_n276), .A3(new_n268), .ZN(new_n277));
  INV_X1    g076(.A(new_n271), .ZN(new_n278));
  INV_X1    g077(.A(new_n259), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n272), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  OAI211_X1 g081(.A(KEYINPUT72), .B(new_n259), .C1(new_n270), .C2(new_n271), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AND2_X1   g083(.A1(G226gat), .A2(G233gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT29), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n285), .B1(new_n244), .B2(new_n286), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n287), .A2(KEYINPUT74), .ZN(new_n288));
  XNOR2_X1  g087(.A(G197gat), .B(G204gat), .ZN(new_n289));
  INV_X1    g088(.A(G211gat), .ZN(new_n290));
  INV_X1    g089(.A(G218gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n289), .B1(KEYINPUT22), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G211gat), .B(G218gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n244), .A2(new_n285), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n287), .A2(KEYINPUT74), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n288), .A2(new_n296), .A3(new_n297), .A4(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G8gat), .B(G36gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(G64gat), .B(G92gat), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n300), .B(new_n301), .Z(new_n302));
  XOR2_X1   g101(.A(KEYINPUT73), .B(KEYINPUT29), .Z(new_n303));
  AND2_X1   g102(.A1(new_n244), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n297), .B1(new_n304), .B2(new_n285), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(new_n295), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n299), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT30), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n302), .B1(new_n299), .B2(new_n306), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n299), .A2(KEYINPUT30), .A3(new_n302), .A4(new_n306), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G225gat), .A2(G233gat), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n314), .B(KEYINPUT78), .Z(new_n315));
  NOR2_X1   g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT75), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT2), .ZN(new_n318));
  INV_X1    g117(.A(G141gat), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n319), .A2(G148gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(G148gat), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n318), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n317), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT76), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT76), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n317), .A2(new_n322), .A3(new_n326), .A4(new_n323), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT77), .B(G148gat), .ZN(new_n329));
  MUX2_X1   g128(.A(G148gat), .B(new_n329), .S(G141gat), .Z(new_n330));
  INV_X1    g129(.A(new_n316), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n323), .B1(new_n331), .B2(KEYINPUT2), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n334), .A2(new_n251), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n325), .A2(new_n327), .B1(new_n330), .B2(new_n332), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(new_n249), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n315), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n334), .A2(KEYINPUT3), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n251), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n315), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n336), .A2(new_n344), .A3(new_n345), .A4(new_n249), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n342), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT4), .B1(new_n334), .B2(new_n251), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n336), .A2(new_n345), .A3(new_n249), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n348), .A2(KEYINPUT79), .A3(new_n349), .ZN(new_n350));
  OAI211_X1 g149(.A(KEYINPUT5), .B(new_n338), .C1(new_n347), .C2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT5), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n342), .A2(new_n352), .A3(new_n343), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n335), .A2(new_n355), .A3(new_n345), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n349), .A2(KEYINPUT80), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT81), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n336), .A2(new_n249), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(KEYINPUT4), .ZN(new_n360));
  AOI211_X1 g159(.A(KEYINPUT81), .B(new_n345), .C1(new_n336), .C2(new_n249), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n356), .B(new_n357), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n354), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n351), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G1gat), .B(G29gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(KEYINPUT0), .ZN(new_n366));
  XNOR2_X1  g165(.A(G57gat), .B(G85gat), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n366), .B(new_n367), .Z(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n364), .A2(KEYINPUT6), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n364), .A2(new_n369), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT6), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n351), .A2(new_n363), .A3(new_n368), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n313), .B1(new_n370), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G78gat), .B(G106gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT31), .B(G50gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(G22gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n303), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT82), .B1(new_n295), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n340), .ZN(new_n382));
  NOR3_X1   g181(.A1(new_n295), .A2(KEYINPUT82), .A3(new_n380), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n334), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT83), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n386), .B(new_n334), .C1(new_n382), .C2(new_n383), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n296), .B1(new_n341), .B2(new_n303), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n385), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G228gat), .A2(G233gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT84), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n340), .B1(new_n295), .B2(KEYINPUT29), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n391), .B1(new_n334), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n393), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n395), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n397), .A2(new_n388), .A3(KEYINPUT84), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n379), .B1(new_n392), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n378), .B1(new_n400), .B2(KEYINPUT85), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n392), .A2(new_n399), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(G22gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n392), .A2(new_n399), .A3(new_n379), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n403), .A2(KEYINPUT85), .A3(new_n404), .A4(new_n378), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n284), .A2(new_n375), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT35), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n272), .A2(new_n280), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT35), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n408), .A2(new_n375), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n411), .A2(KEYINPUT36), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n415), .B1(KEYINPUT36), .B2(new_n284), .ZN(new_n416));
  INV_X1    g215(.A(new_n408), .ZN(new_n417));
  INV_X1    g216(.A(new_n375), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n313), .A2(new_n371), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT86), .ZN(new_n421));
  AOI211_X1 g220(.A(KEYINPUT39), .B(new_n343), .C1(new_n362), .C2(new_n342), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(new_n369), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n343), .B1(new_n362), .B2(new_n342), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT39), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n426), .A2(KEYINPUT86), .A3(new_n368), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n335), .A2(new_n337), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT39), .B1(new_n429), .B2(new_n315), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT40), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT87), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n435), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n428), .A2(new_n437), .A3(new_n432), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n420), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  XOR2_X1   g238(.A(KEYINPUT88), .B(KEYINPUT38), .Z(new_n440));
  INV_X1    g239(.A(KEYINPUT37), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n302), .A2(new_n441), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n310), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n299), .A2(new_n306), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT37), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n440), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n288), .A2(new_n295), .A3(new_n297), .A4(new_n298), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n441), .B1(new_n305), .B2(new_n296), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n440), .B(new_n449), .C1(new_n310), .C2(new_n442), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n374), .A2(new_n450), .A3(new_n370), .A4(new_n307), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n408), .B1(new_n446), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n419), .B1(new_n439), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n414), .B1(new_n416), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(G50gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(G43gat), .ZN(new_n456));
  INV_X1    g255(.A(G43gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(G50gat), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT15), .ZN(new_n459));
  OR3_X1    g258(.A1(new_n456), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  XOR2_X1   g259(.A(KEYINPUT91), .B(G36gat), .Z(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(G29gat), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT92), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(new_n455), .A3(G43gat), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT92), .B1(new_n457), .B2(G50gat), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n459), .B(new_n464), .C1(new_n465), .C2(new_n456), .ZN(new_n466));
  OR3_X1    g265(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AND4_X1   g268(.A1(new_n460), .A2(new_n462), .A3(new_n466), .A4(new_n469), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n468), .A2(KEYINPUT90), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n468), .A2(KEYINPUT90), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n460), .B1(new_n473), .B2(new_n462), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G15gat), .B(G22gat), .ZN(new_n476));
  INV_X1    g275(.A(G1gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT16), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n476), .A2(G1gat), .ZN(new_n481));
  OAI21_X1  g280(.A(G8gat), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(G8gat), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n479), .B(new_n483), .C1(G1gat), .C2(new_n476), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT93), .B1(new_n475), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n473), .A2(new_n462), .ZN(new_n487));
  INV_X1    g286(.A(new_n460), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n460), .A2(new_n462), .A3(new_n466), .A4(new_n469), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT93), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n482), .A2(new_n484), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n486), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n475), .A2(new_n485), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n498));
  NAND2_X1  g297(.A1(G229gat), .A2(G233gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n491), .A2(KEYINPUT17), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT17), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n504), .B1(new_n489), .B2(new_n490), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n485), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n506), .A2(new_n495), .A3(KEYINPUT18), .A4(new_n499), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT18), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n495), .ZN(new_n510));
  INV_X1    g309(.A(new_n499), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT94), .ZN(new_n513));
  XNOR2_X1  g312(.A(G113gat), .B(G141gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(G169gat), .B(G197gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n518), .B(KEYINPUT12), .Z(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n508), .B(new_n512), .C1(new_n513), .C2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n512), .A2(new_n502), .A3(new_n507), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n502), .A2(new_n513), .A3(new_n507), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n523), .A3(new_n519), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G57gat), .B(G64gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G71gat), .ZN(new_n528));
  INV_X1    g327(.A(G78gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G71gat), .A2(G78gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT9), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n527), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n531), .B(new_n530), .C1(new_n526), .C2(new_n533), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n538), .A2(KEYINPUT21), .ZN(new_n539));
  NAND2_X1  g338(.A1(G231gat), .A2(G233gat), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n539), .B(new_n540), .Z(new_n541));
  INV_X1    g340(.A(G127gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n493), .B1(KEYINPUT21), .B2(new_n538), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n546));
  INV_X1    g345(.A(G155gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G183gat), .B(G211gat), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n548), .B(new_n549), .Z(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n545), .A2(new_n551), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n543), .A2(new_n544), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n543), .A2(new_n544), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n554), .A3(new_n550), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n557), .A2(KEYINPUT41), .ZN(new_n558));
  XNOR2_X1  g357(.A(G134gat), .B(G162gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT99), .ZN(new_n562));
  AND2_X1   g361(.A1(G99gat), .A2(G106gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(G99gat), .A2(G106gat), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n566));
  NAND2_X1  g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n562), .A2(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n571));
  INV_X1    g370(.A(G85gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT97), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT97), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(G85gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n571), .A2(new_n573), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n566), .A2(new_n567), .B1(new_n578), .B2(KEYINPUT8), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT99), .B1(new_n563), .B2(new_n564), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n570), .A2(new_n577), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  OR2_X1    g380(.A1(G99gat), .A2(G106gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(new_n562), .A3(new_n578), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT7), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AND2_X1   g385(.A1(G85gat), .A2(G92gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n587), .A3(new_n569), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n577), .A2(new_n579), .A3(new_n583), .A4(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n580), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n581), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT100), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n581), .A2(new_n591), .A3(KEYINPUT100), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n594), .B(new_n595), .C1(new_n503), .C2(new_n505), .ZN(new_n596));
  XOR2_X1   g395(.A(G190gat), .B(G218gat), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n491), .A2(new_n592), .B1(KEYINPUT41), .B2(new_n557), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n598), .B1(new_n596), .B2(new_n599), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n561), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n602), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n604), .A2(new_n560), .A3(new_n600), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n581), .A2(new_n591), .A3(new_n537), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n537), .B1(new_n581), .B2(new_n591), .ZN(new_n608));
  NOR3_X1   g407(.A1(new_n607), .A2(new_n608), .A3(KEYINPUT10), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(KEYINPUT10), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(KEYINPUT101), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n589), .A2(new_n590), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n589), .A2(new_n590), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n538), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n581), .A2(new_n591), .A3(new_n537), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n620), .A3(new_n610), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n612), .A2(new_n613), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n613), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n623), .B1(new_n607), .B2(new_n608), .ZN(new_n624));
  XNOR2_X1  g423(.A(G120gat), .B(G148gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT102), .ZN(new_n626));
  XNOR2_X1  g425(.A(G176gat), .B(G204gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n622), .A2(new_n624), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n613), .B1(new_n609), .B2(new_n611), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n624), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n628), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n556), .A2(new_n606), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n454), .A2(new_n525), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n374), .A2(new_n370), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(new_n477), .ZN(G1324gat));
  INV_X1    g439(.A(new_n313), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT103), .ZN(new_n643));
  AOI21_X1  g442(.A(KEYINPUT42), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT16), .B(G8gat), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n646), .ZN(new_n648));
  OAI21_X1  g447(.A(G8gat), .B1(new_n637), .B2(new_n641), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n647), .B(new_n648), .C1(new_n651), .C2(new_n652), .ZN(G1325gat));
  NAND2_X1  g452(.A1(new_n284), .A2(KEYINPUT36), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(KEYINPUT36), .B2(new_n411), .ZN(new_n655));
  OAI21_X1  g454(.A(G15gat), .B1(new_n637), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n411), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n657), .A2(G15gat), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n637), .B2(new_n658), .ZN(G1326gat));
  NOR2_X1   g458(.A1(new_n637), .A2(new_n408), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT43), .B(G22gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(G1327gat));
  NOR2_X1   g461(.A1(new_n408), .A2(new_n375), .ZN(new_n663));
  AND4_X1   g462(.A1(new_n370), .A2(new_n374), .A3(new_n450), .A4(new_n307), .ZN(new_n664));
  INV_X1    g463(.A(new_n446), .ZN(new_n665));
  AOI22_X1  g464(.A1(new_n664), .A2(new_n665), .B1(new_n407), .B2(new_n406), .ZN(new_n666));
  INV_X1    g465(.A(new_n420), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n437), .B1(new_n428), .B2(new_n432), .ZN(new_n668));
  AOI211_X1 g467(.A(new_n435), .B(new_n431), .C1(new_n423), .C2(new_n427), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n663), .B1(new_n666), .B2(new_n670), .ZN(new_n671));
  AOI22_X1  g470(.A1(new_n671), .A2(new_n655), .B1(new_n410), .B2(new_n413), .ZN(new_n672));
  INV_X1    g471(.A(new_n606), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n556), .ZN(new_n675));
  INV_X1    g474(.A(new_n525), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n675), .A2(new_n676), .A3(new_n635), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(G29gat), .ZN(new_n679));
  INV_X1    g478(.A(new_n638), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT45), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n683), .B1(new_n672), .B2(new_n673), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n453), .A2(new_n416), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n408), .A2(new_n411), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n418), .A2(KEYINPUT35), .ZN(new_n688));
  AOI22_X1  g487(.A1(new_n687), .A2(new_n688), .B1(new_n409), .B2(KEYINPUT35), .ZN(new_n689));
  OAI211_X1 g488(.A(KEYINPUT44), .B(new_n606), .C1(new_n685), .C2(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n684), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n677), .B(KEYINPUT105), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(G29gat), .B1(new_n693), .B2(new_n638), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n682), .A2(new_n694), .ZN(G1328gat));
  NOR2_X1   g494(.A1(new_n641), .A2(new_n461), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n678), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n461), .B1(new_n693), .B2(new_n641), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(G1329gat));
  NAND4_X1  g500(.A1(new_n684), .A2(new_n690), .A3(new_n416), .A4(new_n692), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(G43gat), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n657), .A2(G43gat), .ZN(new_n704));
  AND4_X1   g503(.A1(new_n454), .A2(new_n606), .A3(new_n704), .A4(new_n677), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT47), .B1(new_n707), .B2(KEYINPUT106), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n705), .B1(new_n702), .B2(G43gat), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT47), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n708), .A2(new_n712), .ZN(G1330gat));
  NAND3_X1  g512(.A1(new_n678), .A2(new_n455), .A3(new_n417), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n684), .A2(new_n690), .A3(new_n417), .A4(new_n692), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(G50gat), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT48), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1331gat));
  NAND2_X1  g518(.A1(new_n676), .A2(new_n635), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n556), .A2(new_n720), .A3(new_n606), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n454), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n638), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT107), .B(G57gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1332gat));
  INV_X1    g524(.A(new_n722), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n313), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT49), .B(G64gat), .Z(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT108), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n728), .B(new_n732), .C1(new_n727), .C2(new_n729), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(G1333gat));
  NOR3_X1   g533(.A1(new_n722), .A2(G71gat), .A3(new_n657), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n726), .A2(new_n416), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(G71gat), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n408), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(new_n529), .ZN(G1335gat));
  NOR2_X1   g539(.A1(new_n675), .A2(new_n525), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT51), .B1(new_n674), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n674), .A2(KEYINPUT51), .A3(new_n741), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n674), .A2(KEYINPUT51), .A3(new_n741), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT109), .B1(new_n747), .B2(new_n742), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n573), .A2(new_n575), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n638), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n746), .A2(new_n748), .A3(new_n635), .A4(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n675), .A2(new_n720), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n691), .A2(new_n680), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n749), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n754), .ZN(G1336gat));
  NOR3_X1   g554(.A1(new_n641), .A2(G92gat), .A3(new_n634), .ZN(new_n756));
  XOR2_X1   g555(.A(new_n756), .B(KEYINPUT110), .Z(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n747), .B2(new_n742), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n684), .A2(new_n690), .A3(new_n313), .A4(new_n752), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n571), .A2(new_n576), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT52), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n758), .A2(new_n764), .A3(new_n761), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(G1337gat));
  NOR2_X1   g565(.A1(new_n657), .A2(G99gat), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n746), .A2(new_n748), .A3(new_n635), .A4(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n691), .A2(new_n416), .A3(new_n752), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G99gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(G1338gat));
  NOR3_X1   g570(.A1(new_n408), .A2(G106gat), .A3(new_n634), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n772), .B(KEYINPUT111), .Z(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n747), .B2(new_n742), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n684), .A2(new_n690), .A3(new_n417), .A4(new_n752), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G106gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT53), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n774), .A2(new_n779), .A3(new_n776), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(G1339gat));
  NAND4_X1  g580(.A1(new_n675), .A2(new_n676), .A3(new_n673), .A4(new_n634), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n619), .A2(new_n623), .A3(new_n610), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n783), .A2(KEYINPUT54), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n622), .A2(new_n784), .ZN(new_n785));
  AOI211_X1 g584(.A(KEYINPUT54), .B(new_n623), .C1(new_n619), .C2(new_n610), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n786), .A2(new_n787), .A3(new_n629), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n789), .B(new_n613), .C1(new_n609), .C2(new_n611), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT112), .B1(new_n790), .B2(new_n628), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n785), .B(KEYINPUT55), .C1(new_n788), .C2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(new_n793), .A3(new_n630), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n793), .B1(new_n792), .B2(new_n630), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n495), .A2(new_n496), .A3(new_n500), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n510), .A2(new_n511), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n495), .A2(KEYINPUT114), .A3(new_n496), .A4(new_n500), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n518), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n512), .A2(new_n502), .A3(new_n507), .A4(new_n520), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n803), .A2(new_n605), .A3(new_n603), .A4(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n787), .B1(new_n786), .B2(new_n629), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n790), .A2(KEYINPUT112), .A3(new_n628), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n806), .A2(new_n807), .B1(new_n622), .B2(new_n784), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n808), .A2(KEYINPUT55), .ZN(new_n809));
  NOR4_X1   g608(.A1(new_n795), .A2(new_n796), .A3(new_n805), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n792), .A2(new_n630), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT113), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n785), .B1(new_n788), .B2(new_n791), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n812), .A2(new_n525), .A3(new_n794), .A4(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n635), .A2(new_n803), .A3(new_n804), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n810), .B1(new_n818), .B2(new_n673), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n782), .B1(new_n819), .B2(new_n675), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(new_n687), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n638), .A2(new_n313), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(G113gat), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n823), .A2(new_n824), .A3(new_n676), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n820), .A2(new_n680), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n408), .A3(new_n284), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n829), .A2(new_n641), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n525), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n825), .B1(new_n832), .B2(new_n824), .ZN(G1340gat));
  INV_X1    g632(.A(G120gat), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n823), .A2(new_n834), .A3(new_n634), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n831), .A2(new_n635), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(new_n834), .ZN(G1341gat));
  OAI21_X1  g636(.A(G127gat), .B1(new_n823), .B2(new_n556), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n829), .A2(new_n641), .A3(new_n830), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n675), .A2(new_n542), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(G1342gat));
  INV_X1    g640(.A(KEYINPUT56), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n673), .A2(G134gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n831), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n823), .B2(new_n673), .ZN(new_n845));
  XOR2_X1   g644(.A(new_n845), .B(KEYINPUT116), .Z(new_n846));
  INV_X1    g645(.A(new_n843), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT56), .B1(new_n839), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n844), .A2(new_n846), .A3(new_n848), .ZN(G1343gat));
  AND2_X1   g648(.A1(new_n655), .A2(new_n822), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n820), .A2(new_n417), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n417), .A2(KEYINPUT57), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT117), .B1(new_n808), .B2(KEYINPUT55), .ZN(new_n855));
  INV_X1    g654(.A(new_n630), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n808), .B2(KEYINPUT55), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n813), .A2(new_n858), .A3(new_n814), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n855), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n855), .A2(new_n857), .A3(KEYINPUT118), .A4(new_n859), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n525), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n606), .B1(new_n864), .B2(new_n817), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n556), .B1(new_n865), .B2(new_n810), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n854), .B1(new_n866), .B2(new_n782), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n853), .B1(new_n867), .B2(KEYINPUT119), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n869));
  AOI211_X1 g668(.A(new_n869), .B(new_n854), .C1(new_n866), .C2(new_n782), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n525), .B(new_n850), .C1(new_n868), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(G141gat), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n416), .A2(new_n408), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n826), .A2(new_n641), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n676), .A2(G141gat), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT120), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT58), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n872), .A2(new_n879), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(G1344gat));
  NAND3_X1  g680(.A1(new_n874), .A2(new_n329), .A3(new_n635), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT121), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n782), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n408), .A2(KEYINPUT57), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n884), .A2(new_n885), .B1(new_n851), .B2(KEYINPUT57), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n635), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n850), .B(KEYINPUT122), .ZN(new_n888));
  OAI211_X1 g687(.A(KEYINPUT59), .B(G148gat), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n850), .B1(new_n868), .B2(new_n870), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n634), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n329), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n883), .B(new_n889), .C1(new_n892), .C2(KEYINPUT59), .ZN(G1345gat));
  OAI21_X1  g692(.A(G155gat), .B1(new_n890), .B2(new_n556), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n874), .A2(new_n547), .A3(new_n675), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1346gat));
  INV_X1    g695(.A(G162gat), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n890), .A2(new_n897), .A3(new_n673), .ZN(new_n898));
  AOI21_X1  g697(.A(G162gat), .B1(new_n874), .B2(new_n606), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(G1347gat));
  AND2_X1   g699(.A1(new_n820), .A2(new_n638), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n284), .A2(new_n313), .A3(new_n408), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n204), .A3(new_n525), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n638), .A2(new_n313), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT123), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n821), .A2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n525), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n909), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT124), .B1(new_n909), .B2(G169gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n904), .B1(new_n910), .B2(new_n911), .ZN(G1348gat));
  NAND3_X1  g711(.A1(new_n903), .A2(new_n205), .A3(new_n635), .ZN(new_n913));
  OAI21_X1  g712(.A(G176gat), .B1(new_n907), .B2(new_n634), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1349gat));
  NOR2_X1   g714(.A1(new_n556), .A2(new_n213), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n903), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(G183gat), .B1(new_n907), .B2(new_n556), .ZN(new_n918));
  NAND2_X1  g717(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT126), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n920), .B(new_n923), .ZN(G1350gat));
  INV_X1    g723(.A(G190gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n903), .A2(new_n925), .A3(new_n606), .ZN(new_n926));
  OAI21_X1  g725(.A(G190gat), .B1(new_n907), .B2(new_n673), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n927), .A2(KEYINPUT61), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(KEYINPUT61), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(G1351gat));
  AND3_X1   g729(.A1(new_n901), .A2(new_n313), .A3(new_n873), .ZN(new_n931));
  INV_X1    g730(.A(G197gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n931), .A2(new_n932), .A3(new_n525), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n655), .A2(new_n906), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n886), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT127), .B1(new_n936), .B2(new_n676), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G197gat), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n936), .A2(KEYINPUT127), .A3(new_n676), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n933), .B1(new_n938), .B2(new_n939), .ZN(G1352gat));
  INV_X1    g739(.A(G204gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n931), .A2(new_n941), .A3(new_n635), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n942), .A2(KEYINPUT62), .ZN(new_n943));
  OAI21_X1  g742(.A(G204gat), .B1(new_n887), .B2(new_n934), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(KEYINPUT62), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(G1353gat));
  NAND3_X1  g745(.A1(new_n931), .A2(new_n290), .A3(new_n675), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n886), .A2(new_n675), .A3(new_n935), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n948), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT63), .B1(new_n948), .B2(G211gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(G1354gat));
  OAI21_X1  g750(.A(G218gat), .B1(new_n936), .B2(new_n673), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n931), .A2(new_n291), .A3(new_n606), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1355gat));
endmodule


