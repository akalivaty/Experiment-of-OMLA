//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT66), .Z(new_n211));
  NAND2_X1  g0011(.A1(G107), .A2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G68), .B2(G238), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G87), .A2(G250), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G58), .A2(G232), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n211), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  AND2_X1   g0019(.A1(G97), .A2(G257), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n209), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT65), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n203), .A2(G50), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n209), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT0), .Z(new_n231));
  NOR3_X1   g0031(.A1(new_n222), .A2(new_n228), .A3(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT76), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT76), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G294), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT67), .B(G1698), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n255), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n251), .A2(KEYINPUT3), .A3(new_n252), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n254), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT86), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G1), .A3(G13), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI211_X1 g0066(.A(KEYINPUT86), .B(new_n254), .C1(new_n256), .C2(new_n260), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n263), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT5), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT5), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G1), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n270), .A2(new_n272), .A3(new_n273), .A4(G45), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  OR2_X1    g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n274), .A2(new_n265), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G264), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n268), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G190), .ZN(new_n280));
  OR2_X1    g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n259), .A2(new_n283), .A3(new_n224), .A4(G87), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT22), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n206), .A2(G20), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT23), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n287), .B(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n253), .A2(G116), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n286), .B(new_n289), .C1(G20), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n224), .A2(G87), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n260), .A2(new_n285), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n282), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n295));
  AND2_X1   g0095(.A1(KEYINPUT76), .A2(G33), .ZN(new_n296));
  NOR2_X1   g0096(.A1(KEYINPUT76), .A2(G33), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n295), .B1(new_n298), .B2(KEYINPUT3), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n299), .A2(KEYINPUT22), .A3(new_n224), .A4(G87), .ZN(new_n300));
  INV_X1    g0100(.A(G116), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n302), .A2(new_n224), .B1(new_n285), .B2(new_n284), .ZN(new_n303));
  INV_X1    g0103(.A(new_n282), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n300), .A2(new_n303), .A3(new_n289), .A4(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n223), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n294), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n307), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n273), .A2(G33), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n273), .A2(G13), .A3(G20), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G107), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n311), .A2(G107), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT25), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n308), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n279), .A2(G200), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n281), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n279), .A2(G169), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT87), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n268), .A2(G179), .A3(new_n276), .A4(new_n278), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n322), .B1(new_n321), .B2(new_n323), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n308), .A2(new_n314), .A3(new_n316), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n320), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT14), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n273), .B1(G41), .B2(G45), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n265), .A2(G238), .A3(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n273), .B(G274), .C1(G41), .C2(G45), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n331), .A2(KEYINPUT72), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(KEYINPUT72), .B1(new_n331), .B2(new_n332), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n258), .A2(G33), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n295), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G226), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT67), .ZN(new_n339));
  INV_X1    g0139(.A(G1698), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n338), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n234), .A2(new_n340), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n337), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G33), .A2(G97), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT71), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(KEYINPUT71), .A2(G33), .A3(G97), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n265), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT13), .B1(new_n335), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n259), .A2(new_n283), .ZN(new_n354));
  AND2_X1   g0154(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n355));
  NOR2_X1   g0155(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n356));
  OAI21_X1  g0156(.A(G226), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n344), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n354), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n266), .B1(new_n359), .B2(new_n350), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT13), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n360), .B(new_n361), .C1(new_n334), .C2(new_n333), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n353), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n329), .B1(new_n363), .B2(G169), .ZN(new_n364));
  INV_X1    g0164(.A(G169), .ZN(new_n365));
  AOI211_X1 g0165(.A(KEYINPUT14), .B(new_n365), .C1(new_n353), .C2(new_n362), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n353), .A2(KEYINPUT73), .A3(new_n362), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT73), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n370), .B(KEYINPUT13), .C1(new_n335), .C2(new_n352), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n368), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n250), .A2(G20), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G77), .ZN(new_n376));
  INV_X1    g0176(.A(G50), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n224), .A2(new_n250), .ZN(new_n378));
  OAI221_X1 g0178(.A(new_n376), .B1(new_n224), .B2(G68), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n307), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT11), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT74), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n307), .B1(new_n273), .B2(G20), .ZN(new_n383));
  OR3_X1    g0183(.A1(new_n311), .A2(KEYINPUT12), .A3(G68), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT12), .B1(new_n311), .B2(G68), .ZN(new_n385));
  AOI22_X1  g0185(.A1(G68), .A2(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n381), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n382), .B1(new_n381), .B2(new_n386), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n374), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n381), .A2(new_n386), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n369), .A2(new_n371), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(G190), .ZN(new_n395));
  INV_X1    g0195(.A(G200), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n353), .B2(new_n362), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n392), .A2(new_n399), .ZN(new_n400));
  XOR2_X1   g0200(.A(new_n400), .B(KEYINPUT75), .Z(new_n401));
  NOR2_X1   g0201(.A1(new_n311), .A2(G77), .ZN(new_n402));
  INV_X1    g0202(.A(new_n383), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(new_n213), .ZN(new_n404));
  XOR2_X1   g0204(.A(KEYINPUT15), .B(G87), .Z(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n375), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT70), .ZN(new_n407));
  XOR2_X1   g0207(.A(KEYINPUT8), .B(G58), .Z(new_n408));
  INV_X1    g0208(.A(new_n378), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n408), .A2(new_n409), .B1(G20), .B2(G77), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  AOI211_X1 g0211(.A(new_n402), .B(new_n404), .C1(new_n411), .C2(new_n307), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G238), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n355), .A2(new_n356), .ZN(new_n415));
  OAI221_X1 g0215(.A(new_n337), .B1(new_n414), .B2(new_n340), .C1(new_n234), .C2(new_n415), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n416), .B(new_n266), .C1(G107), .C2(new_n337), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n265), .A2(new_n330), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n417), .B(new_n332), .C1(new_n214), .C2(new_n419), .ZN(new_n420));
  XNOR2_X1  g0220(.A(KEYINPUT68), .B(G179), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n365), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n413), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n401), .A2(new_n425), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n408), .A2(new_n375), .B1(G150), .B2(new_n409), .ZN(new_n427));
  OAI21_X1  g0227(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n311), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n429), .A2(new_n307), .B1(new_n377), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n383), .A2(G50), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT9), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n255), .A2(G222), .B1(G223), .B2(G1698), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n265), .B1(new_n435), .B2(new_n337), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(G77), .B2(new_n337), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n437), .B(new_n332), .C1(new_n338), .C2(new_n419), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G200), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n434), .B(new_n439), .C1(new_n280), .C2(new_n438), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT10), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n438), .A2(new_n422), .ZN(new_n442));
  XNOR2_X1  g0242(.A(new_n442), .B(KEYINPUT69), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n438), .A2(new_n365), .B1(new_n432), .B2(new_n431), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n420), .A2(G200), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n412), .B(new_n447), .C1(new_n280), .C2(new_n420), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT16), .ZN(new_n450));
  INV_X1    g0250(.A(G68), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT3), .B1(new_n251), .B2(new_n252), .ZN(new_n452));
  OAI211_X1 g0252(.A(KEYINPUT7), .B(new_n224), .C1(new_n452), .C2(new_n336), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT7), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n337), .B2(G20), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n451), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G58), .A2(G68), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT77), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT77), .B1(G58), .B2(G68), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n459), .A2(new_n202), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G159), .ZN(new_n462));
  OAI22_X1  g0262(.A1(new_n461), .A2(new_n224), .B1(new_n462), .B2(new_n378), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n450), .B1(new_n456), .B2(new_n463), .ZN(new_n464));
  OR3_X1    g0264(.A1(new_n459), .A2(new_n202), .A3(new_n460), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n465), .A2(G20), .B1(G159), .B2(new_n409), .ZN(new_n466));
  AOI21_X1  g0266(.A(G20), .B1(new_n257), .B2(new_n259), .ZN(new_n467));
  OAI21_X1  g0267(.A(G68), .B1(new_n467), .B2(new_n454), .ZN(new_n468));
  AOI211_X1 g0268(.A(KEYINPUT7), .B(G20), .C1(new_n257), .C2(new_n259), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n466), .B(KEYINPUT16), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n464), .A2(new_n307), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n403), .A2(new_n408), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n430), .B2(new_n408), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n418), .A2(G232), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G87), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(G223), .B1(new_n355), .B2(new_n356), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G226), .A2(G1698), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n477), .B1(new_n299), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n332), .B(new_n475), .C1(new_n481), .C2(new_n265), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G169), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n255), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n476), .B1(new_n484), .B2(new_n260), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n266), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n486), .A2(new_n422), .A3(new_n332), .A4(new_n475), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n474), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT18), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(KEYINPUT78), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT78), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n471), .A2(new_n473), .B1(new_n483), .B2(new_n487), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n492), .B1(new_n493), .B2(KEYINPUT18), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(KEYINPUT18), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n491), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n482), .A2(new_n396), .ZN(new_n497));
  XNOR2_X1  g0297(.A(KEYINPUT79), .B(G190), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n486), .A2(new_n499), .A3(new_n332), .A4(new_n475), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(new_n471), .A3(new_n473), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT17), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n501), .A2(new_n471), .A3(KEYINPUT17), .A4(new_n473), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n504), .A2(KEYINPUT80), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT80), .B1(new_n504), .B2(new_n505), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n496), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OR3_X1    g0308(.A1(new_n446), .A2(new_n449), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n426), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n430), .A2(new_n301), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n309), .A2(G116), .A3(new_n310), .A4(new_n311), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n306), .A2(new_n223), .B1(G20), .B2(new_n301), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G283), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n514), .B(new_n224), .C1(G33), .C2(new_n205), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n513), .A2(KEYINPUT20), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT20), .B1(new_n513), .B2(new_n515), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n511), .B(new_n512), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n274), .A2(G270), .A3(new_n265), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(G257), .B1(new_n355), .B2(new_n356), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G264), .A2(G1698), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n299), .A2(new_n524), .B1(G303), .B2(new_n354), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n276), .B(new_n521), .C1(new_n525), .C2(new_n265), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n519), .B1(new_n526), .B2(new_n499), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n354), .A2(G303), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n255), .A2(G257), .B1(G264), .B2(G1698), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n529), .B2(new_n260), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n520), .B1(new_n530), .B2(new_n266), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n396), .B1(new_n531), .B2(new_n276), .ZN(new_n532));
  OAI21_X1  g0332(.A(KEYINPUT83), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n526), .A2(G200), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n531), .A2(new_n276), .A3(new_n498), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT83), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n519), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n526), .A2(G169), .A3(new_n518), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT21), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n526), .A2(new_n368), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n518), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n526), .A2(KEYINPUT21), .A3(G169), .A4(new_n518), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT84), .B1(new_n538), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n533), .A2(new_n537), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT84), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n214), .B1(new_n341), .B2(new_n342), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT4), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n552), .A2(new_n257), .A3(new_n553), .A4(new_n259), .ZN(new_n554));
  OAI21_X1  g0354(.A(G244), .B1(new_n355), .B2(new_n356), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT4), .B1(new_n555), .B2(new_n354), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n337), .A2(G250), .A3(G1698), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n514), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT82), .ZN(new_n560));
  INV_X1    g0360(.A(new_n514), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n561), .B1(new_n554), .B2(new_n556), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT82), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n563), .A3(new_n558), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n560), .A2(new_n266), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n277), .A2(G257), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n276), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n365), .ZN(new_n570));
  XNOR2_X1  g0370(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G97), .A2(G107), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n207), .A3(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n205), .A2(G107), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n573), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  OAI22_X1  g0375(.A1(new_n575), .A2(new_n224), .B1(new_n213), .B2(new_n378), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n206), .B1(new_n453), .B2(new_n455), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n307), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n313), .A2(G97), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n430), .A2(new_n205), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n565), .A2(new_n421), .A3(new_n568), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n570), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n581), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n565), .A2(G190), .A3(new_n568), .ZN(new_n585));
  AND4_X1   g0385(.A1(new_n563), .A2(new_n557), .A3(new_n514), .A4(new_n558), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n563), .B1(new_n562), .B2(new_n558), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n567), .B1(new_n588), .B2(new_n266), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n584), .B(new_n585), .C1(new_n589), .C2(new_n396), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n405), .A2(new_n311), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT19), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n346), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n257), .A2(new_n224), .A3(G68), .A4(new_n259), .ZN(new_n594));
  AOI21_X1  g0394(.A(G20), .B1(new_n350), .B2(KEYINPUT19), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n207), .A2(G87), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n593), .B(new_n594), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n591), .B1(new_n597), .B2(new_n307), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n313), .A2(new_n405), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(G45), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n601), .A2(new_n275), .A3(G1), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n265), .B(G250), .C1(G1), .C2(new_n601), .ZN(new_n604));
  OAI22_X1  g0404(.A1(new_n415), .A2(new_n414), .B1(new_n214), .B2(new_n340), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n302), .B1(new_n605), .B2(new_n299), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n603), .B(new_n604), .C1(new_n606), .C2(new_n265), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n365), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n255), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n290), .B1(new_n609), .B2(new_n260), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n266), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n611), .A2(new_n421), .A3(new_n603), .A4(new_n604), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n600), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n607), .A2(G200), .ZN(new_n614));
  INV_X1    g0414(.A(G87), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n312), .A2(new_n615), .ZN(new_n616));
  AOI211_X1 g0416(.A(new_n591), .B(new_n616), .C1(new_n597), .C2(new_n307), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n611), .A2(G190), .A3(new_n603), .A4(new_n604), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n614), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n583), .A2(new_n590), .A3(new_n621), .ZN(new_n622));
  AND4_X1   g0422(.A1(new_n328), .A2(new_n510), .A3(new_n551), .A4(new_n622), .ZN(G372));
  NOR2_X1   g0423(.A1(new_n489), .A2(new_n490), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n493), .A2(KEYINPUT18), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n504), .A2(new_n505), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT80), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n504), .A2(KEYINPUT80), .A3(new_n505), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n425), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n399), .A2(new_n634), .B1(new_n374), .B2(new_n391), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n627), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n636), .A2(new_n441), .B1(new_n444), .B2(new_n443), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n426), .A2(new_n509), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT88), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n317), .B1(new_n321), .B2(new_n323), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n639), .B1(new_n640), .B2(new_n545), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n321), .A2(new_n323), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n327), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(KEYINPUT88), .A3(new_n547), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n583), .A2(new_n590), .A3(new_n319), .A4(new_n621), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n582), .A2(new_n581), .ZN(new_n648));
  AOI21_X1  g0448(.A(G169), .B1(new_n565), .B2(new_n568), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT26), .B1(new_n650), .B2(new_n621), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  NOR4_X1   g0452(.A1(new_n648), .A2(new_n620), .A3(new_n649), .A4(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n613), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n637), .B1(new_n638), .B2(new_n655), .ZN(G369));
  INV_X1    g0456(.A(G330), .ZN(new_n657));
  INV_X1    g0457(.A(G13), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(G20), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n273), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G213), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(new_n519), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n549), .B1(new_n547), .B2(new_n548), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n547), .A2(new_n668), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n657), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n642), .A2(KEYINPUT87), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(new_n327), .A3(new_n676), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n317), .A2(KEYINPUT89), .A3(new_n666), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT89), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n327), .B2(new_n665), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n677), .A2(new_n681), .A3(new_n319), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n326), .A2(new_n327), .A3(new_n665), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n674), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n640), .A2(new_n666), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n547), .A2(new_n665), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n677), .A2(new_n681), .A3(new_n319), .A4(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n685), .A2(new_n686), .A3(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n229), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n596), .A2(new_n301), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n691), .A2(new_n692), .A3(new_n273), .ZN(new_n693));
  INV_X1    g0493(.A(new_n227), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(new_n691), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT28), .Z(new_n696));
  NAND4_X1  g0496(.A1(new_n328), .A2(new_n551), .A3(new_n622), .A4(new_n666), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n268), .A2(new_n278), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n531), .A2(G179), .A3(new_n276), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n698), .A2(new_n699), .A3(new_n607), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(new_n589), .A3(KEYINPUT30), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  INV_X1    g0502(.A(new_n607), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n542), .A2(new_n703), .A3(new_n278), .A4(new_n268), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n702), .B1(new_n704), .B2(new_n569), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n422), .B1(new_n531), .B2(new_n276), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n569), .A2(new_n706), .A3(new_n279), .A4(new_n607), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n701), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT31), .B1(new_n708), .B2(new_n665), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT91), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI211_X1 g0511(.A(KEYINPUT91), .B(KEYINPUT31), .C1(new_n708), .C2(new_n665), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n697), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n708), .A2(KEYINPUT31), .A3(new_n665), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT90), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n714), .B(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(G330), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n646), .B1(new_n677), .B2(new_n547), .ZN(new_n718));
  OAI211_X1 g0518(.A(KEYINPUT29), .B(new_n666), .C1(new_n718), .C2(new_n654), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n622), .A2(new_n319), .A3(new_n641), .A4(new_n644), .ZN(new_n720));
  INV_X1    g0520(.A(new_n613), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n652), .B1(new_n583), .B2(new_n620), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n650), .A2(KEYINPUT26), .A3(new_n621), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n665), .B1(new_n720), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n719), .B1(KEYINPUT29), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n717), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n696), .B1(new_n728), .B2(G1), .ZN(G364));
  NOR2_X1   g0529(.A1(new_n224), .A2(G179), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(new_n280), .A3(G200), .ZN(new_n731));
  INV_X1    g0531(.A(G283), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n280), .A2(G179), .A3(G200), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(new_n224), .ZN(new_n734));
  INV_X1    g0534(.A(G294), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n354), .B1(new_n731), .B2(new_n732), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G311), .ZN(new_n737));
  OR3_X1    g0537(.A1(new_n421), .A2(KEYINPUT93), .A3(new_n224), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT93), .B1(new_n421), .B2(new_n224), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n396), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G190), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n741), .A2(new_n499), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G322), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n737), .A2(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n730), .A2(new_n280), .A3(new_n396), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n736), .B(new_n747), .C1(G329), .C2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n730), .A2(G190), .A3(G200), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(KEYINPUT96), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(KEYINPUT96), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G303), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n396), .B1(new_n738), .B2(new_n739), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(KEYINPUT94), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(KEYINPUT94), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n758), .A2(new_n498), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT95), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n758), .A2(KEYINPUT95), .A3(new_n498), .A4(new_n759), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G326), .ZN(new_n765));
  AND3_X1   g0565(.A1(new_n758), .A2(new_n280), .A3(new_n759), .ZN(new_n766));
  XNOR2_X1  g0566(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(G317), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n750), .A2(new_n756), .A3(new_n765), .A4(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n764), .A2(G50), .B1(G87), .B2(new_n755), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n734), .A2(new_n205), .B1(new_n731), .B2(new_n206), .ZN(new_n772));
  OR3_X1    g0572(.A1(new_n748), .A2(KEYINPUT32), .A3(new_n462), .ZN(new_n773));
  OAI21_X1  g0573(.A(KEYINPUT32), .B1(new_n748), .B2(new_n462), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n773), .A2(new_n337), .A3(new_n774), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n772), .B(new_n775), .C1(new_n742), .C2(G77), .ZN(new_n776));
  INV_X1    g0576(.A(new_n766), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n771), .B(new_n776), .C1(new_n451), .C2(new_n777), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n744), .A2(G58), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n770), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n223), .B1(G20), .B2(new_n365), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G20), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n781), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n694), .A2(new_n601), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n299), .A2(new_n690), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n786), .B(new_n787), .C1(new_n247), .C2(new_n601), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n337), .A2(G355), .A3(new_n229), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n788), .B(new_n789), .C1(G116), .C2(new_n229), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n780), .A2(new_n781), .B1(new_n785), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n659), .A2(G45), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n792), .A2(KEYINPUT92), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(KEYINPUT92), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n793), .A2(G1), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n691), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n671), .A2(new_n673), .A3(new_n784), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n791), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n667), .B1(new_n546), .B2(new_n550), .ZN(new_n799));
  OAI21_X1  g0599(.A(G330), .B1(new_n799), .B2(new_n672), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n671), .A2(new_n657), .A3(new_n673), .ZN(new_n801));
  INV_X1    g0601(.A(new_n796), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n798), .A2(new_n803), .ZN(G396));
  NOR2_X1   g0604(.A1(new_n412), .A2(new_n666), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n425), .B1(new_n449), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n634), .A2(new_n666), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(KEYINPUT98), .B1(new_n725), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n725), .A2(new_n808), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n809), .B(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(new_n717), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n796), .ZN(new_n813));
  INV_X1    g0613(.A(new_n781), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n764), .A2(G137), .B1(G150), .B2(new_n766), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n462), .B2(new_n743), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G143), .B2(new_n744), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT34), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G50), .B2(new_n755), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n749), .A2(G132), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n731), .A2(new_n451), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n260), .ZN(new_n822));
  INV_X1    g0622(.A(new_n734), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G58), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n819), .A2(new_n820), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n764), .A2(G303), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n354), .B1(new_n745), .B2(new_n735), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G283), .B2(new_n766), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n742), .A2(G116), .ZN(new_n829));
  INV_X1    g0629(.A(new_n731), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(G87), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n754), .B2(new_n206), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n734), .A2(new_n205), .B1(new_n748), .B2(new_n737), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n826), .A2(new_n828), .A3(new_n829), .A4(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n814), .B1(new_n825), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n781), .A2(new_n782), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n808), .A2(new_n783), .B1(G77), .B2(new_n838), .ZN(new_n839));
  NOR3_X1   g0639(.A1(new_n836), .A2(new_n802), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n813), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G384));
  INV_X1    g0642(.A(KEYINPUT38), .ZN(new_n843));
  INV_X1    g0643(.A(new_n663), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n470), .A2(new_n307), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT7), .B1(new_n299), .B2(G20), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n467), .A2(new_n454), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n846), .A2(G68), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT16), .B1(new_n848), .B2(new_n466), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n473), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n844), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n632), .B2(new_n496), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n464), .A2(new_n307), .A3(new_n470), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n854), .A2(new_n851), .B1(new_n488), .B2(new_n844), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT37), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n855), .A2(new_n856), .A3(new_n502), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n850), .A2(new_n851), .B1(new_n488), .B2(new_n844), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n856), .B1(new_n858), .B2(new_n502), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n843), .B1(new_n853), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n852), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n508), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n860), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(KEYINPUT38), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n397), .B(new_n393), .C1(new_n394), .C2(G190), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n391), .B(new_n665), .C1(new_n374), .C2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n665), .B1(new_n388), .B2(new_n389), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n372), .A2(new_n364), .A3(new_n366), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n399), .B(new_n869), .C1(new_n870), .C2(new_n390), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n808), .ZN(new_n873));
  INV_X1    g0673(.A(new_n714), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n874), .A2(new_n709), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n873), .B1(new_n875), .B2(new_n697), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n866), .A2(new_n876), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n877), .A2(KEYINPUT40), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n474), .B(new_n844), .C1(new_n626), .C2(new_n628), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n856), .B1(new_n855), .B2(new_n502), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n857), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g0682(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n865), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(new_n876), .A3(KEYINPUT40), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT102), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n885), .A2(new_n876), .A3(KEYINPUT102), .A4(KEYINPUT40), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n875), .A2(new_n697), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n878), .A2(new_n890), .A3(new_n510), .A4(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n878), .A2(new_n890), .A3(G330), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n510), .A2(G330), .A3(new_n891), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n892), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n861), .B2(new_n865), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n843), .B(new_n860), .C1(new_n508), .C2(new_n862), .ZN(new_n899));
  INV_X1    g0699(.A(new_n883), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n879), .B2(new_n881), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n899), .A2(KEYINPUT39), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT101), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n392), .A2(new_n665), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n863), .B2(new_n864), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT39), .B1(new_n905), .B2(new_n899), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT101), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n884), .A2(new_n865), .A3(new_n897), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n903), .A2(new_n904), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n807), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n725), .B2(new_n806), .ZN(new_n912));
  INV_X1    g0712(.A(new_n872), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n914), .A2(new_n866), .B1(new_n626), .B2(new_n663), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n896), .B(new_n916), .Z(new_n917));
  OR2_X1    g0717(.A1(new_n638), .A2(new_n726), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n637), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n917), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n273), .B2(new_n659), .ZN(new_n921));
  NOR4_X1   g0721(.A1(new_n227), .A2(new_n459), .A3(new_n213), .A4(new_n460), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n201), .A2(new_n451), .ZN(new_n923));
  OAI211_X1 g0723(.A(G1), .B(new_n658), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT35), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n226), .B1(new_n575), .B2(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n926), .B(G116), .C1(new_n925), .C2(new_n575), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT99), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT36), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n921), .A2(new_n924), .A3(new_n929), .ZN(G367));
  INV_X1    g0730(.A(new_n785), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n240), .B2(new_n787), .ZN(new_n932));
  INV_X1    g0732(.A(new_n405), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n932), .B1(new_n229), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT103), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n617), .A2(new_n666), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n935), .B1(new_n621), .B2(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n936), .A2(new_n613), .ZN(new_n938));
  MUX2_X1   g0738(.A(new_n935), .B(new_n937), .S(new_n938), .Z(new_n939));
  AOI21_X1  g0739(.A(new_n802), .B1(new_n939), .B2(new_n784), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n830), .A2(G77), .B1(new_n749), .B2(G137), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n777), .B2(new_n462), .ZN(new_n942));
  AOI211_X1 g0742(.A(new_n354), .B(new_n942), .C1(G58), .C2(new_n755), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n744), .A2(G150), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n764), .A2(G143), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n742), .A2(new_n201), .B1(G68), .B2(new_n823), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n943), .A2(new_n944), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n731), .A2(new_n205), .ZN(new_n948));
  INV_X1    g0748(.A(new_n764), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n949), .A2(new_n737), .B1(new_n206), .B2(new_n734), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n948), .B(new_n950), .C1(G317), .C2(new_n749), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n744), .A2(G303), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT46), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n754), .B2(new_n301), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n755), .A2(KEYINPUT46), .A3(G116), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n954), .B(new_n955), .C1(new_n777), .C2(new_n735), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT108), .Z(new_n957));
  NAND4_X1  g0757(.A1(new_n951), .A2(new_n260), .A3(new_n952), .A4(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n743), .A2(new_n732), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n947), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT47), .Z(new_n961));
  OAI211_X1 g0761(.A(new_n934), .B(new_n940), .C1(new_n961), .C2(new_n814), .ZN(new_n962));
  INV_X1    g0762(.A(new_n687), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n682), .A2(new_n683), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n688), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT106), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n965), .A2(new_n966), .A3(new_n800), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n688), .B(new_n964), .C1(new_n674), .C2(KEYINPUT106), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(KEYINPUT107), .B1(new_n727), .B2(new_n969), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n967), .A2(new_n968), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT107), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n971), .A2(new_n972), .A3(new_n717), .A4(new_n726), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT45), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n688), .A2(new_n686), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n583), .A2(new_n590), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n581), .A2(new_n665), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n570), .A2(new_n581), .A3(new_n582), .A4(new_n665), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(KEYINPUT104), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n582), .A2(new_n581), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT104), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n980), .A2(new_n981), .A3(new_n570), .A4(new_n665), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n976), .A2(new_n977), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n974), .B1(new_n975), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NOR3_X1   g0785(.A1(new_n975), .A2(new_n983), .A3(new_n974), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n975), .A2(new_n983), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT44), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT44), .B1(new_n975), .B2(new_n983), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n985), .A2(new_n986), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n685), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n685), .B1(new_n989), .B2(new_n990), .C1(new_n986), .C2(new_n985), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n970), .A2(new_n973), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n728), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n691), .B(KEYINPUT41), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n795), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(KEYINPUT42), .B1(new_n983), .B2(new_n688), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n979), .A2(new_n982), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n583), .A2(new_n590), .A3(new_n977), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n677), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n650), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n999), .B1(new_n1004), .B2(new_n665), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT105), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OR3_X1    g0807(.A1(new_n983), .A2(KEYINPUT42), .A3(new_n688), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n999), .B(KEYINPUT105), .C1(new_n1004), .C2(new_n665), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT43), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n939), .A2(new_n1011), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n939), .A2(new_n1011), .ZN(new_n1013));
  AND3_X1   g0813(.A1(new_n1010), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1012), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1014), .A2(new_n1015), .B1(new_n685), .B2(new_n983), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1017), .A2(new_n1011), .A3(new_n939), .A4(new_n1008), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1010), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1018), .A2(new_n992), .A3(new_n1002), .A4(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n962), .B1(new_n998), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(KEYINPUT109), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT109), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1024), .B(new_n962), .C1(new_n998), .C2(new_n1021), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1025), .ZN(G387));
  AOI22_X1  g0826(.A1(new_n764), .A2(G322), .B1(G311), .B2(new_n766), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n744), .A2(G317), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n742), .A2(G303), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT48), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n823), .A2(G283), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n755), .A2(G294), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n731), .A2(new_n301), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n299), .B(new_n1038), .C1(G326), .C2(new_n749), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n408), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n777), .A2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n948), .B(new_n1043), .C1(G159), .C2(new_n764), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n823), .A2(new_n405), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n755), .A2(G77), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n745), .B2(new_n377), .C1(new_n451), .C2(new_n743), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(G150), .B2(new_n749), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1044), .A2(new_n299), .A3(new_n1045), .A4(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n814), .B1(new_n1041), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n787), .B1(new_n237), .B2(new_n601), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n692), .A2(new_n229), .A3(new_n337), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AOI211_X1 g0853(.A(G45), .B(new_n692), .C1(G68), .C2(G77), .ZN(new_n1054));
  OAI21_X1  g0854(.A(KEYINPUT50), .B1(new_n1042), .B2(G50), .ZN(new_n1055));
  OR3_X1    g0855(.A1(new_n1042), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1053), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n690), .A2(new_n206), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n931), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n1050), .A2(new_n802), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n682), .A2(new_n683), .A3(new_n784), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1061), .A2(new_n1062), .B1(new_n795), .B2(new_n971), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n970), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n973), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n691), .B1(new_n728), .B2(new_n971), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1063), .A2(new_n1066), .ZN(G393));
  NAND2_X1  g0867(.A1(new_n993), .A2(new_n994), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1069), .A2(new_n691), .A3(new_n995), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n802), .B1(new_n983), .B2(new_n784), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n787), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1072), .A2(new_n244), .B1(new_n205), .B2(new_n229), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1071), .B1(new_n931), .B2(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n354), .B1(new_n746), .B2(new_n748), .C1(new_n754), .C2(new_n732), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n764), .A2(G317), .B1(G311), .B2(new_n744), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  XOR2_X1   g0877(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n1078));
  AOI21_X1  g0878(.A(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n766), .A2(G303), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n742), .A2(G294), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n734), .A2(new_n301), .B1(new_n731), .B2(new_n206), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1078), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1082), .B1(new_n1076), .B2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .A4(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n764), .A2(G150), .B1(G159), .B2(new_n744), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT51), .Z(new_n1087));
  NAND2_X1  g0887(.A1(new_n749), .A2(G143), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n742), .A2(new_n408), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n831), .B1(new_n754), .B2(new_n451), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n734), .A2(new_n213), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1090), .A2(new_n260), .A3(new_n1091), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .A4(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n201), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n777), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1085), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1074), .B1(new_n1096), .B2(new_n781), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1068), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1097), .B1(new_n1098), .B2(new_n795), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1070), .A2(new_n1099), .ZN(G390));
  NAND2_X1  g0900(.A1(new_n806), .A2(new_n807), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n871), .B2(new_n868), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n891), .A2(G330), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(KEYINPUT112), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT112), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n876), .A2(new_n1105), .A3(G330), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n666), .B1(new_n647), .B2(new_n654), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n807), .B1(new_n1109), .B2(new_n1101), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n904), .B1(new_n1110), .B2(new_n872), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n903), .B2(new_n909), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n904), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n885), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n718), .A2(new_n654), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1115), .A2(new_n665), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n911), .B1(new_n1116), .B2(new_n806), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1114), .B1(new_n1118), .B2(new_n872), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1108), .B1(new_n1112), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1113), .B1(new_n912), .B2(new_n913), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n907), .B1(new_n906), .B2(new_n908), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1113), .B(new_n885), .C1(new_n1117), .C2(new_n913), .ZN(new_n1125));
  OAI211_X1 g0925(.A(G330), .B(new_n808), .C1(new_n713), .C2(new_n716), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1126), .A2(new_n913), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1120), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1127), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n891), .A2(G330), .A3(new_n808), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n913), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1130), .A2(new_n1117), .A3(new_n1132), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1126), .A2(new_n913), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1110), .B1(new_n1134), .B2(new_n1107), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(KEYINPUT113), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1126), .A2(new_n913), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1137), .A2(new_n1106), .A3(new_n1104), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT113), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(new_n1139), .A3(new_n1110), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1133), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n918), .A2(new_n637), .A3(new_n894), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1129), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1130), .A2(new_n1117), .A3(new_n1132), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1140), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1139), .B1(new_n1138), .B2(new_n1110), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1144), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1120), .A2(new_n1128), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1142), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1143), .A2(new_n691), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n783), .B1(new_n903), .B2(new_n909), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n1042), .B2(new_n837), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n745), .A2(new_n301), .B1(new_n615), .B2(new_n754), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1091), .B(new_n1154), .C1(G294), .C2(new_n749), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n337), .B(new_n821), .C1(new_n742), .C2(G97), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(new_n206), .C2(new_n777), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G283), .B2(new_n764), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n766), .A2(G137), .ZN(new_n1159));
  INV_X1    g0959(.A(G128), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1159), .B1(new_n949), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n354), .B1(new_n749), .B2(G125), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n1094), .B2(new_n731), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT114), .Z(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT54), .B(G143), .Z(new_n1165));
  AOI22_X1  g0965(.A1(new_n742), .A2(new_n1165), .B1(G159), .B2(new_n823), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n744), .A2(G132), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1164), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n755), .A2(G150), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1169), .B(new_n1170), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1161), .A2(new_n1168), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n781), .B1(new_n1158), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1153), .A2(new_n796), .A3(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT116), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1148), .A2(new_n795), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1151), .A2(new_n1175), .A3(new_n1176), .ZN(G378));
  INV_X1    g0977(.A(KEYINPUT57), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n878), .A2(new_n890), .A3(G330), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n433), .A2(new_n844), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n446), .B(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1181), .B(new_n1182), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n910), .A2(new_n915), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1183), .B1(new_n910), .B2(new_n915), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1179), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1183), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n916), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n910), .A2(new_n915), .A3(new_n1183), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(new_n893), .A3(new_n1189), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1186), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1142), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1178), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1149), .B1(new_n1129), .B2(new_n1141), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1186), .A2(new_n1190), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(KEYINPUT57), .A3(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1193), .A2(new_n691), .A3(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n764), .A2(G125), .B1(G150), .B2(new_n823), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT119), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n744), .A2(G128), .B1(new_n755), .B2(new_n1165), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT118), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n766), .A2(G132), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n742), .A2(G137), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1199), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  XOR2_X1   g1004(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1205));
  XNOR2_X1  g1005(.A(new_n1204), .B(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(G41), .B1(new_n830), .B2(G159), .ZN(new_n1207));
  AOI21_X1  g1007(.A(G33), .B1(new_n749), .B2(G124), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n299), .B1(new_n766), .B2(G97), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n745), .A2(new_n206), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(KEYINPUT117), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(new_n269), .A3(new_n1212), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n743), .A2(new_n933), .B1(new_n451), .B2(new_n734), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n830), .A2(G58), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1046), .B(new_n1215), .C1(new_n732), .C2(new_n748), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1216), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(KEYINPUT117), .B2(new_n1211), .C1(new_n301), .C2(new_n949), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT58), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(G41), .B1(new_n296), .B2(KEYINPUT3), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1209), .B(new_n1220), .C1(G50), .C2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n781), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n802), .B1(new_n1094), .B2(new_n837), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(KEYINPUT121), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1187), .B2(new_n782), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(KEYINPUT121), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1224), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1195), .B2(new_n795), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1197), .A2(new_n1230), .ZN(G375));
  NAND2_X1  g1031(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1142), .B(new_n1144), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n997), .A3(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1045), .B1(new_n745), .B2(new_n732), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT123), .Z(new_n1236));
  AOI22_X1  g1036(.A1(new_n766), .A2(G116), .B1(G107), .B2(new_n742), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n337), .B1(new_n830), .B2(G77), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1239), .A2(KEYINPUT122), .B1(G303), .B2(new_n749), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1236), .A2(new_n1237), .A3(new_n1240), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n764), .A2(G294), .B1(G97), .B2(new_n755), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(KEYINPUT122), .C2(new_n1239), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n764), .A2(G132), .B1(G159), .B2(new_n755), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n742), .A2(G150), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n766), .A2(new_n1165), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1215), .A2(new_n299), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n734), .A2(new_n377), .B1(new_n748), .B2(new_n1160), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(new_n744), .C2(G137), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .A4(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n814), .B1(new_n1243), .B2(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n872), .A2(new_n783), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n838), .A2(G68), .ZN(new_n1253));
  NOR4_X1   g1053(.A1(new_n1251), .A2(new_n802), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1147), .B2(new_n795), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1234), .A2(new_n1255), .ZN(G381));
  AND3_X1   g1056(.A1(new_n1151), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(new_n1197), .A3(new_n1230), .ZN(new_n1258));
  NOR4_X1   g1058(.A1(new_n1258), .A2(G384), .A3(G387), .A4(G381), .ZN(new_n1259));
  INV_X1    g1059(.A(G390), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(G393), .A2(G396), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(G407));
  OAI211_X1 g1062(.A(G407), .B(G213), .C1(G343), .C2(new_n1258), .ZN(G409));
  NAND2_X1  g1063(.A1(new_n664), .A2(G213), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1194), .A2(new_n997), .A3(new_n1195), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1230), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1264), .B1(G378), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(G378), .B2(G375), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n664), .A2(G213), .A3(G2897), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT60), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1233), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1141), .A2(KEYINPUT60), .A3(new_n1142), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1272), .A2(new_n1273), .A3(new_n1232), .A4(new_n691), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1274), .A2(G384), .A3(new_n1255), .ZN(new_n1275));
  AOI21_X1  g1075(.A(G384), .B1(new_n1274), .B2(new_n1255), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1270), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1274), .A2(new_n1255), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n841), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1274), .A2(G384), .A3(new_n1255), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1279), .A2(new_n1280), .A3(new_n1269), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1277), .A2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(KEYINPUT63), .B1(new_n1268), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G375), .A2(G378), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1265), .A2(new_n1230), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n1257), .A2(new_n1285), .B1(G213), .B2(new_n664), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1284), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1283), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT125), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1025), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n997), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(new_n995), .B2(new_n728), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1020), .B(new_n1016), .C1(new_n1293), .C2(new_n795), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1024), .B1(new_n1294), .B2(new_n962), .ZN(new_n1295));
  OAI211_X1 g1095(.A(KEYINPUT124), .B(new_n1260), .C1(new_n1291), .C2(new_n1295), .ZN(new_n1296));
  AOI22_X1  g1096(.A1(new_n1063), .A2(new_n1066), .B1(new_n803), .B2(new_n798), .ZN(new_n1297));
  OR2_X1    g1097(.A1(new_n1261), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1294), .A2(G390), .A3(new_n962), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(G387), .A2(new_n1260), .B1(KEYINPUT124), .B2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1290), .B1(new_n1299), .B2(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1260), .B1(new_n1291), .B2(new_n1295), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1300), .A2(KEYINPUT124), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1305), .A2(KEYINPUT125), .A3(new_n1298), .A4(new_n1296), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1302), .A2(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1261), .A2(new_n1297), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1300), .ZN(new_n1309));
  AOI21_X1  g1109(.A(G390), .B1(new_n1294), .B2(new_n962), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1308), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT61), .B1(new_n1307), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT63), .ZN(new_n1313));
  OAI21_X1  g1113(.A(KEYINPUT126), .B1(new_n1288), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT126), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1268), .A2(new_n1315), .A3(KEYINPUT63), .A4(new_n1287), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1289), .A2(new_n1312), .A3(new_n1314), .A4(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1288), .A2(KEYINPUT62), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT61), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1257), .B1(new_n1230), .B2(new_n1197), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1281), .B(new_n1277), .C1(new_n1320), .C2(new_n1267), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT62), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1284), .A2(new_n1286), .A3(new_n1322), .A4(new_n1287), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1318), .A2(new_n1319), .A3(new_n1321), .A4(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1306), .ZN(new_n1325));
  AOI21_X1  g1125(.A(G390), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1308), .B1(new_n1326), .B2(KEYINPUT124), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT125), .B1(new_n1327), .B2(new_n1305), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1311), .B1(new_n1325), .B2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1324), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1317), .A2(new_n1331), .ZN(G405));
  NAND2_X1  g1132(.A1(new_n1329), .A2(KEYINPUT127), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1284), .A2(new_n1258), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1334), .B1(new_n1276), .B2(new_n1275), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1284), .A2(new_n1258), .A3(new_n1287), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT127), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1307), .A2(new_n1338), .A3(new_n1311), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1333), .A2(new_n1337), .A3(new_n1339), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1329), .A2(new_n1335), .A3(KEYINPUT127), .A4(new_n1336), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(G402));
endmodule


