

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X2 U550 ( .A(n714), .Z(n516) );
  NAND2_X1 U551 ( .A1(n739), .A2(n740), .ZN(n714) );
  NAND2_X1 U552 ( .A1(n722), .A2(G286), .ZN(n713) );
  INV_X1 U553 ( .A(KEYINPUT93), .ZN(n712) );
  XNOR2_X2 U554 ( .A(n524), .B(KEYINPUT65), .ZN(n588) );
  XOR2_X1 U555 ( .A(n696), .B(KEYINPUT28), .Z(n517) );
  XOR2_X1 U556 ( .A(n710), .B(KEYINPUT31), .Z(n518) );
  OR2_X1 U557 ( .A1(G301), .A2(n707), .ZN(n519) );
  AND2_X1 U558 ( .A1(n688), .A2(G1996), .ZN(n676) );
  OR2_X1 U559 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U560 ( .A1(n982), .A2(n679), .ZN(n685) );
  NAND2_X1 U561 ( .A1(n711), .A2(n518), .ZN(n722) );
  XNOR2_X1 U562 ( .A(n713), .B(n712), .ZN(n719) );
  NAND2_X1 U563 ( .A1(n719), .A2(n718), .ZN(n720) );
  INV_X1 U564 ( .A(KEYINPUT92), .ZN(n728) );
  INV_X1 U565 ( .A(G2105), .ZN(n523) );
  NOR2_X1 U566 ( .A1(G543), .A2(G651), .ZN(n630) );
  XOR2_X1 U567 ( .A(KEYINPUT17), .B(n526), .Z(n882) );
  NOR2_X1 U568 ( .A1(n627), .A2(G651), .ZN(n638) );
  NOR2_X1 U569 ( .A1(n530), .A2(n529), .ZN(G160) );
  AND2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n885) );
  NAND2_X1 U571 ( .A1(G113), .A2(n885), .ZN(n522) );
  NOR2_X1 U572 ( .A1(n523), .A2(G2104), .ZN(n520) );
  XNOR2_X1 U573 ( .A(n520), .B(KEYINPUT64), .ZN(n886) );
  NAND2_X1 U574 ( .A1(G125), .A2(n886), .ZN(n521) );
  NAND2_X1 U575 ( .A1(n522), .A2(n521), .ZN(n530) );
  NAND2_X1 U576 ( .A1(n523), .A2(G2104), .ZN(n524) );
  NAND2_X1 U577 ( .A1(G101), .A2(n588), .ZN(n525) );
  XOR2_X1 U578 ( .A(n525), .B(KEYINPUT23), .Z(n528) );
  NOR2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  NAND2_X1 U580 ( .A1(n882), .A2(G137), .ZN(n527) );
  NAND2_X1 U581 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U582 ( .A1(n630), .A2(G89), .ZN(n531) );
  XNOR2_X1 U583 ( .A(n531), .B(KEYINPUT4), .ZN(n534) );
  INV_X1 U584 ( .A(G651), .ZN(n536) );
  XOR2_X1 U585 ( .A(KEYINPUT0), .B(G543), .Z(n627) );
  OR2_X1 U586 ( .A1(n536), .A2(n627), .ZN(n532) );
  XOR2_X1 U587 ( .A(KEYINPUT66), .B(n532), .Z(n631) );
  NAND2_X1 U588 ( .A1(G76), .A2(n631), .ZN(n533) );
  NAND2_X1 U589 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U590 ( .A(n535), .B(KEYINPUT5), .ZN(n542) );
  NOR2_X1 U591 ( .A1(G543), .A2(n536), .ZN(n537) );
  XOR2_X1 U592 ( .A(KEYINPUT1), .B(n537), .Z(n634) );
  NAND2_X1 U593 ( .A1(G63), .A2(n634), .ZN(n539) );
  NAND2_X1 U594 ( .A1(G51), .A2(n638), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U596 ( .A(KEYINPUT6), .B(n540), .Z(n541) );
  NAND2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U598 ( .A(n543), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U599 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U600 ( .A1(n634), .A2(G64), .ZN(n544) );
  XNOR2_X1 U601 ( .A(n544), .B(KEYINPUT68), .ZN(n546) );
  NAND2_X1 U602 ( .A1(G52), .A2(n638), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U604 ( .A(KEYINPUT69), .B(n547), .Z(n552) );
  NAND2_X1 U605 ( .A1(G77), .A2(n631), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n630), .A2(G90), .ZN(n548) );
  NAND2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U608 ( .A(KEYINPUT9), .B(n550), .Z(n551) );
  NOR2_X1 U609 ( .A1(n552), .A2(n551), .ZN(G171) );
  AND2_X1 U610 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U611 ( .A(G132), .ZN(G219) );
  INV_X1 U612 ( .A(G82), .ZN(G220) );
  INV_X1 U613 ( .A(G120), .ZN(G236) );
  INV_X1 U614 ( .A(G69), .ZN(G235) );
  INV_X1 U615 ( .A(G108), .ZN(G238) );
  NAND2_X1 U616 ( .A1(G7), .A2(G661), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n553), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U618 ( .A(G223), .ZN(n810) );
  NAND2_X1 U619 ( .A1(n810), .A2(G567), .ZN(n554) );
  XOR2_X1 U620 ( .A(KEYINPUT11), .B(n554), .Z(G234) );
  NAND2_X1 U621 ( .A1(n630), .A2(G81), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(KEYINPUT12), .ZN(n557) );
  NAND2_X1 U623 ( .A1(G68), .A2(n631), .ZN(n556) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(KEYINPUT13), .B(n558), .Z(n562) );
  NAND2_X1 U626 ( .A1(G56), .A2(n634), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(KEYINPUT71), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n560), .B(KEYINPUT14), .ZN(n561) );
  NOR2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n564) );
  NAND2_X1 U630 ( .A1(n638), .A2(G43), .ZN(n563) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n982) );
  INV_X1 U632 ( .A(G860), .ZN(n600) );
  OR2_X1 U633 ( .A1(n982), .A2(n600), .ZN(G153) );
  INV_X1 U634 ( .A(G171), .ZN(G301) );
  NAND2_X1 U635 ( .A1(G868), .A2(G301), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n631), .A2(G79), .ZN(n571) );
  NAND2_X1 U637 ( .A1(G66), .A2(n634), .ZN(n566) );
  NAND2_X1 U638 ( .A1(G92), .A2(n630), .ZN(n565) );
  NAND2_X1 U639 ( .A1(n566), .A2(n565), .ZN(n569) );
  NAND2_X1 U640 ( .A1(n638), .A2(G54), .ZN(n567) );
  XOR2_X1 U641 ( .A(KEYINPUT72), .B(n567), .Z(n568) );
  NOR2_X1 U642 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U643 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U644 ( .A(n572), .B(KEYINPUT15), .ZN(n981) );
  OR2_X1 U645 ( .A1(n981), .A2(G868), .ZN(n573) );
  NAND2_X1 U646 ( .A1(n574), .A2(n573), .ZN(G284) );
  NAND2_X1 U647 ( .A1(G65), .A2(n634), .ZN(n576) );
  NAND2_X1 U648 ( .A1(G53), .A2(n638), .ZN(n575) );
  NAND2_X1 U649 ( .A1(n576), .A2(n575), .ZN(n580) );
  NAND2_X1 U650 ( .A1(G91), .A2(n630), .ZN(n578) );
  NAND2_X1 U651 ( .A1(G78), .A2(n631), .ZN(n577) );
  NAND2_X1 U652 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U653 ( .A1(n580), .A2(n579), .ZN(n994) );
  XOR2_X1 U654 ( .A(n994), .B(KEYINPUT70), .Z(G299) );
  NOR2_X1 U655 ( .A1(G299), .A2(G868), .ZN(n582) );
  INV_X1 U656 ( .A(G868), .ZN(n649) );
  NOR2_X1 U657 ( .A1(G286), .A2(n649), .ZN(n581) );
  NOR2_X1 U658 ( .A1(n582), .A2(n581), .ZN(G297) );
  NAND2_X1 U659 ( .A1(n600), .A2(G559), .ZN(n583) );
  NAND2_X1 U660 ( .A1(n583), .A2(n981), .ZN(n584) );
  XNOR2_X1 U661 ( .A(n584), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U662 ( .A1(G868), .A2(n982), .ZN(n587) );
  NAND2_X1 U663 ( .A1(G868), .A2(n981), .ZN(n585) );
  NOR2_X1 U664 ( .A1(G559), .A2(n585), .ZN(n586) );
  NOR2_X1 U665 ( .A1(n587), .A2(n586), .ZN(G282) );
  NAND2_X1 U666 ( .A1(G111), .A2(n885), .ZN(n590) );
  NAND2_X1 U667 ( .A1(G99), .A2(n588), .ZN(n589) );
  NAND2_X1 U668 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U669 ( .A(n591), .B(KEYINPUT73), .ZN(n593) );
  NAND2_X1 U670 ( .A1(G135), .A2(n882), .ZN(n592) );
  NAND2_X1 U671 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n886), .A2(G123), .ZN(n594) );
  XOR2_X1 U673 ( .A(KEYINPUT18), .B(n594), .Z(n595) );
  NOR2_X1 U674 ( .A1(n596), .A2(n595), .ZN(n961) );
  XNOR2_X1 U675 ( .A(G2096), .B(n961), .ZN(n598) );
  INV_X1 U676 ( .A(G2100), .ZN(n597) );
  NAND2_X1 U677 ( .A1(n598), .A2(n597), .ZN(G156) );
  NAND2_X1 U678 ( .A1(G559), .A2(n981), .ZN(n599) );
  XOR2_X1 U679 ( .A(n982), .B(n599), .Z(n646) );
  NAND2_X1 U680 ( .A1(n600), .A2(n646), .ZN(n608) );
  NAND2_X1 U681 ( .A1(G67), .A2(n634), .ZN(n602) );
  NAND2_X1 U682 ( .A1(G55), .A2(n638), .ZN(n601) );
  NAND2_X1 U683 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U684 ( .A(KEYINPUT74), .B(n603), .ZN(n607) );
  NAND2_X1 U685 ( .A1(G93), .A2(n630), .ZN(n605) );
  NAND2_X1 U686 ( .A1(G80), .A2(n631), .ZN(n604) );
  NAND2_X1 U687 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U688 ( .A1(n607), .A2(n606), .ZN(n648) );
  XOR2_X1 U689 ( .A(n608), .B(n648), .Z(G145) );
  NAND2_X1 U690 ( .A1(G88), .A2(n630), .ZN(n610) );
  NAND2_X1 U691 ( .A1(G75), .A2(n631), .ZN(n609) );
  NAND2_X1 U692 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U693 ( .A1(G62), .A2(n634), .ZN(n612) );
  NAND2_X1 U694 ( .A1(G50), .A2(n638), .ZN(n611) );
  NAND2_X1 U695 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U696 ( .A1(n614), .A2(n613), .ZN(G166) );
  XOR2_X1 U697 ( .A(KEYINPUT76), .B(KEYINPUT2), .Z(n616) );
  NAND2_X1 U698 ( .A1(G73), .A2(n631), .ZN(n615) );
  XNOR2_X1 U699 ( .A(n616), .B(n615), .ZN(n620) );
  NAND2_X1 U700 ( .A1(G61), .A2(n634), .ZN(n618) );
  NAND2_X1 U701 ( .A1(G86), .A2(n630), .ZN(n617) );
  NAND2_X1 U702 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U703 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n638), .A2(G48), .ZN(n621) );
  NAND2_X1 U705 ( .A1(n622), .A2(n621), .ZN(G305) );
  NAND2_X1 U706 ( .A1(G49), .A2(n638), .ZN(n624) );
  NAND2_X1 U707 ( .A1(G74), .A2(G651), .ZN(n623) );
  NAND2_X1 U708 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U709 ( .A(KEYINPUT75), .B(n625), .Z(n626) );
  NOR2_X1 U710 ( .A1(n634), .A2(n626), .ZN(n629) );
  NAND2_X1 U711 ( .A1(n627), .A2(G87), .ZN(n628) );
  NAND2_X1 U712 ( .A1(n629), .A2(n628), .ZN(G288) );
  NAND2_X1 U713 ( .A1(G85), .A2(n630), .ZN(n633) );
  NAND2_X1 U714 ( .A1(G72), .A2(n631), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U716 ( .A1(G60), .A2(n634), .ZN(n635) );
  XNOR2_X1 U717 ( .A(KEYINPUT67), .B(n635), .ZN(n636) );
  NOR2_X1 U718 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n638), .A2(G47), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(G290) );
  XNOR2_X1 U721 ( .A(G166), .B(KEYINPUT19), .ZN(n645) );
  XOR2_X1 U722 ( .A(G299), .B(n648), .Z(n641) );
  XNOR2_X1 U723 ( .A(G305), .B(n641), .ZN(n642) );
  XNOR2_X1 U724 ( .A(n642), .B(G288), .ZN(n643) );
  XNOR2_X1 U725 ( .A(n643), .B(G290), .ZN(n644) );
  XNOR2_X1 U726 ( .A(n645), .B(n644), .ZN(n827) );
  XOR2_X1 U727 ( .A(n827), .B(n646), .Z(n647) );
  NOR2_X1 U728 ( .A1(n649), .A2(n647), .ZN(n651) );
  AND2_X1 U729 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U730 ( .A1(n651), .A2(n650), .ZN(G295) );
  NAND2_X1 U731 ( .A1(G2084), .A2(G2078), .ZN(n652) );
  XOR2_X1 U732 ( .A(KEYINPUT20), .B(n652), .Z(n653) );
  NAND2_X1 U733 ( .A1(G2090), .A2(n653), .ZN(n655) );
  XOR2_X1 U734 ( .A(KEYINPUT21), .B(KEYINPUT77), .Z(n654) );
  XNOR2_X1 U735 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n656), .A2(G2072), .ZN(n657) );
  XNOR2_X1 U737 ( .A(n657), .B(KEYINPUT78), .ZN(G158) );
  XNOR2_X1 U738 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U739 ( .A1(G235), .A2(G236), .ZN(n658) );
  XNOR2_X1 U740 ( .A(n658), .B(KEYINPUT79), .ZN(n659) );
  NOR2_X1 U741 ( .A1(G238), .A2(n659), .ZN(n660) );
  NAND2_X1 U742 ( .A1(G57), .A2(n660), .ZN(n814) );
  NAND2_X1 U743 ( .A1(n814), .A2(G567), .ZN(n665) );
  NOR2_X1 U744 ( .A1(G220), .A2(G219), .ZN(n661) );
  XOR2_X1 U745 ( .A(KEYINPUT22), .B(n661), .Z(n662) );
  NOR2_X1 U746 ( .A1(G218), .A2(n662), .ZN(n663) );
  NAND2_X1 U747 ( .A1(G96), .A2(n663), .ZN(n815) );
  NAND2_X1 U748 ( .A1(n815), .A2(G2106), .ZN(n664) );
  NAND2_X1 U749 ( .A1(n665), .A2(n664), .ZN(n832) );
  NAND2_X1 U750 ( .A1(G483), .A2(G661), .ZN(n666) );
  NOR2_X1 U751 ( .A1(n832), .A2(n666), .ZN(n813) );
  NAND2_X1 U752 ( .A1(n813), .A2(G36), .ZN(G176) );
  NAND2_X1 U753 ( .A1(G138), .A2(n882), .ZN(n668) );
  NAND2_X1 U754 ( .A1(G102), .A2(n588), .ZN(n667) );
  NAND2_X1 U755 ( .A1(n668), .A2(n667), .ZN(n674) );
  NAND2_X1 U756 ( .A1(n885), .A2(G114), .ZN(n669) );
  XNOR2_X1 U757 ( .A(n669), .B(KEYINPUT80), .ZN(n671) );
  NAND2_X1 U758 ( .A1(G126), .A2(n886), .ZN(n670) );
  NAND2_X1 U759 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U760 ( .A(KEYINPUT81), .B(n672), .Z(n673) );
  NOR2_X1 U761 ( .A1(n674), .A2(n673), .ZN(G164) );
  INV_X1 U762 ( .A(G166), .ZN(G303) );
  NAND2_X1 U763 ( .A1(G40), .A2(G160), .ZN(n675) );
  XOR2_X1 U764 ( .A(n675), .B(KEYINPUT82), .Z(n739) );
  NOR2_X1 U765 ( .A1(G164), .A2(G1384), .ZN(n740) );
  INV_X1 U766 ( .A(n714), .ZN(n688) );
  XNOR2_X1 U767 ( .A(n676), .B(KEYINPUT26), .ZN(n678) );
  AND2_X1 U768 ( .A1(n516), .A2(G1341), .ZN(n677) );
  INV_X1 U769 ( .A(G2067), .ZN(n680) );
  OR2_X1 U770 ( .A1(n516), .A2(n680), .ZN(n682) );
  NAND2_X1 U771 ( .A1(G1348), .A2(n516), .ZN(n681) );
  NAND2_X1 U772 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U773 ( .A(KEYINPUT90), .B(n683), .Z(n686) );
  OR2_X1 U774 ( .A1(n981), .A2(n686), .ZN(n684) );
  NAND2_X1 U775 ( .A1(n685), .A2(n684), .ZN(n694) );
  AND2_X1 U776 ( .A1(n686), .A2(n981), .ZN(n692) );
  NAND2_X1 U777 ( .A1(n688), .A2(G2072), .ZN(n687) );
  XNOR2_X1 U778 ( .A(n687), .B(KEYINPUT27), .ZN(n690) );
  INV_X1 U779 ( .A(G1956), .ZN(n907) );
  NOR2_X1 U780 ( .A1(n907), .A2(n688), .ZN(n689) );
  NOR2_X1 U781 ( .A1(n690), .A2(n689), .ZN(n695) );
  AND2_X1 U782 ( .A1(n994), .A2(n695), .ZN(n691) );
  NOR2_X1 U783 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U784 ( .A1(n694), .A2(n693), .ZN(n697) );
  NOR2_X1 U785 ( .A1(n695), .A2(n994), .ZN(n696) );
  NAND2_X1 U786 ( .A1(n697), .A2(n517), .ZN(n698) );
  XNOR2_X1 U787 ( .A(n698), .B(KEYINPUT29), .ZN(n699) );
  INV_X1 U788 ( .A(n699), .ZN(n703) );
  XOR2_X1 U789 ( .A(KEYINPUT88), .B(G1961), .Z(n917) );
  NAND2_X1 U790 ( .A1(n917), .A2(n516), .ZN(n700) );
  XNOR2_X1 U791 ( .A(n700), .B(KEYINPUT89), .ZN(n702) );
  XOR2_X1 U792 ( .A(KEYINPUT25), .B(G2078), .Z(n942) );
  NOR2_X1 U793 ( .A1(n516), .A2(n942), .ZN(n701) );
  NOR2_X1 U794 ( .A1(n702), .A2(n701), .ZN(n707) );
  NAND2_X1 U795 ( .A1(n703), .A2(n519), .ZN(n711) );
  NAND2_X1 U796 ( .A1(G8), .A2(n516), .ZN(n771) );
  NOR2_X1 U797 ( .A1(G1966), .A2(n771), .ZN(n727) );
  NOR2_X1 U798 ( .A1(G2084), .A2(n516), .ZN(n723) );
  NOR2_X1 U799 ( .A1(n727), .A2(n723), .ZN(n704) );
  NAND2_X1 U800 ( .A1(G8), .A2(n704), .ZN(n705) );
  XNOR2_X1 U801 ( .A(KEYINPUT30), .B(n705), .ZN(n706) );
  NOR2_X1 U802 ( .A1(G168), .A2(n706), .ZN(n709) );
  AND2_X1 U803 ( .A1(G301), .A2(n707), .ZN(n708) );
  NOR2_X1 U804 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U805 ( .A1(G1971), .A2(n771), .ZN(n716) );
  NOR2_X1 U806 ( .A1(G2090), .A2(n516), .ZN(n715) );
  NOR2_X1 U807 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U808 ( .A1(G303), .A2(n717), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n720), .A2(G8), .ZN(n721) );
  XNOR2_X1 U810 ( .A(n721), .B(KEYINPUT32), .ZN(n731) );
  XOR2_X1 U811 ( .A(n722), .B(KEYINPUT91), .Z(n725) );
  NAND2_X1 U812 ( .A1(n723), .A2(G8), .ZN(n724) );
  NAND2_X1 U813 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U814 ( .A1(n727), .A2(n726), .ZN(n729) );
  XNOR2_X1 U815 ( .A(n729), .B(n728), .ZN(n730) );
  NAND2_X1 U816 ( .A1(n731), .A2(n730), .ZN(n767) );
  NOR2_X1 U817 ( .A1(G1976), .A2(G288), .ZN(n735) );
  NOR2_X1 U818 ( .A1(G1971), .A2(G303), .ZN(n732) );
  NOR2_X1 U819 ( .A1(n735), .A2(n732), .ZN(n1001) );
  NAND2_X1 U820 ( .A1(n767), .A2(n1001), .ZN(n733) );
  XNOR2_X1 U821 ( .A(n733), .B(KEYINPUT94), .ZN(n734) );
  NAND2_X1 U822 ( .A1(G1976), .A2(G288), .ZN(n997) );
  NAND2_X1 U823 ( .A1(n734), .A2(n997), .ZN(n764) );
  NAND2_X1 U824 ( .A1(n735), .A2(KEYINPUT33), .ZN(n736) );
  NOR2_X1 U825 ( .A1(n736), .A2(n771), .ZN(n738) );
  XOR2_X1 U826 ( .A(G1981), .B(G305), .Z(n987) );
  INV_X1 U827 ( .A(n987), .ZN(n737) );
  NOR2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n761) );
  INV_X1 U829 ( .A(n739), .ZN(n741) );
  NOR2_X1 U830 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U831 ( .A(KEYINPUT83), .B(n742), .Z(n805) );
  NAND2_X1 U832 ( .A1(G107), .A2(n885), .ZN(n744) );
  NAND2_X1 U833 ( .A1(G119), .A2(n886), .ZN(n743) );
  NAND2_X1 U834 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U835 ( .A(KEYINPUT85), .B(n745), .ZN(n749) );
  NAND2_X1 U836 ( .A1(n882), .A2(G131), .ZN(n747) );
  NAND2_X1 U837 ( .A1(G95), .A2(n588), .ZN(n746) );
  AND2_X1 U838 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U839 ( .A1(n749), .A2(n748), .ZN(n868) );
  NAND2_X1 U840 ( .A1(G1991), .A2(n868), .ZN(n760) );
  NAND2_X1 U841 ( .A1(G105), .A2(n588), .ZN(n750) );
  XNOR2_X1 U842 ( .A(n750), .B(KEYINPUT86), .ZN(n751) );
  XNOR2_X1 U843 ( .A(n751), .B(KEYINPUT38), .ZN(n753) );
  NAND2_X1 U844 ( .A1(G117), .A2(n885), .ZN(n752) );
  NAND2_X1 U845 ( .A1(n753), .A2(n752), .ZN(n757) );
  NAND2_X1 U846 ( .A1(G141), .A2(n882), .ZN(n755) );
  NAND2_X1 U847 ( .A1(G129), .A2(n886), .ZN(n754) );
  NAND2_X1 U848 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U849 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U850 ( .A(KEYINPUT87), .B(n758), .ZN(n871) );
  NAND2_X1 U851 ( .A1(G1996), .A2(n871), .ZN(n759) );
  NAND2_X1 U852 ( .A1(n760), .A2(n759), .ZN(n973) );
  NAND2_X1 U853 ( .A1(n805), .A2(n973), .ZN(n798) );
  AND2_X1 U854 ( .A1(n761), .A2(n798), .ZN(n775) );
  INV_X1 U855 ( .A(n775), .ZN(n762) );
  OR2_X1 U856 ( .A1(n771), .A2(n762), .ZN(n763) );
  NOR2_X1 U857 ( .A1(n764), .A2(n763), .ZN(n779) );
  NOR2_X1 U858 ( .A1(G2090), .A2(G303), .ZN(n765) );
  NAND2_X1 U859 ( .A1(G8), .A2(n765), .ZN(n766) );
  NAND2_X1 U860 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U861 ( .A1(n768), .A2(n771), .ZN(n773) );
  NOR2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n769) );
  XOR2_X1 U863 ( .A(n769), .B(KEYINPUT24), .Z(n770) );
  OR2_X1 U864 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U865 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U866 ( .A1(n774), .A2(n798), .ZN(n777) );
  NAND2_X1 U867 ( .A1(n775), .A2(KEYINPUT33), .ZN(n776) );
  NAND2_X1 U868 ( .A1(n777), .A2(n776), .ZN(n778) );
  OR2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n792) );
  XOR2_X1 U870 ( .A(G1986), .B(G290), .Z(n998) );
  NAND2_X1 U871 ( .A1(n885), .A2(G116), .ZN(n780) );
  XNOR2_X1 U872 ( .A(n780), .B(KEYINPUT84), .ZN(n782) );
  NAND2_X1 U873 ( .A1(G128), .A2(n886), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U875 ( .A(n783), .B(KEYINPUT35), .ZN(n788) );
  NAND2_X1 U876 ( .A1(G140), .A2(n882), .ZN(n785) );
  NAND2_X1 U877 ( .A1(G104), .A2(n588), .ZN(n784) );
  NAND2_X1 U878 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U879 ( .A(KEYINPUT34), .B(n786), .Z(n787) );
  NAND2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U881 ( .A(n789), .B(KEYINPUT36), .ZN(n893) );
  XOR2_X1 U882 ( .A(G2067), .B(KEYINPUT37), .Z(n793) );
  NAND2_X1 U883 ( .A1(n893), .A2(n793), .ZN(n794) );
  NAND2_X1 U884 ( .A1(n998), .A2(n794), .ZN(n790) );
  NAND2_X1 U885 ( .A1(n790), .A2(n805), .ZN(n791) );
  NAND2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n808) );
  NOR2_X1 U887 ( .A1(n893), .A2(n793), .ZN(n969) );
  INV_X1 U888 ( .A(n794), .ZN(n966) );
  NOR2_X1 U889 ( .A1(n871), .A2(G1996), .ZN(n795) );
  XNOR2_X1 U890 ( .A(n795), .B(KEYINPUT95), .ZN(n958) );
  NOR2_X1 U891 ( .A1(G1986), .A2(G290), .ZN(n796) );
  NOR2_X1 U892 ( .A1(G1991), .A2(n868), .ZN(n962) );
  NOR2_X1 U893 ( .A1(n796), .A2(n962), .ZN(n797) );
  XOR2_X1 U894 ( .A(KEYINPUT96), .B(n797), .Z(n799) );
  NAND2_X1 U895 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U896 ( .A1(n958), .A2(n800), .ZN(n801) );
  XNOR2_X1 U897 ( .A(KEYINPUT39), .B(n801), .ZN(n802) );
  NOR2_X1 U898 ( .A1(n966), .A2(n802), .ZN(n803) );
  NOR2_X1 U899 ( .A1(n969), .A2(n803), .ZN(n804) );
  XNOR2_X1 U900 ( .A(KEYINPUT97), .B(n804), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U903 ( .A(n809), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U904 ( .A1(G2106), .A2(n810), .ZN(G217) );
  AND2_X1 U905 ( .A1(G15), .A2(G2), .ZN(n811) );
  NAND2_X1 U906 ( .A1(G661), .A2(n811), .ZN(G259) );
  NAND2_X1 U907 ( .A1(G3), .A2(G1), .ZN(n812) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(G188) );
  NOR2_X1 U909 ( .A1(n815), .A2(n814), .ZN(G325) );
  XNOR2_X1 U910 ( .A(KEYINPUT101), .B(G325), .ZN(G261) );
  INV_X1 U912 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U913 ( .A(G2454), .B(G2446), .ZN(n824) );
  XNOR2_X1 U914 ( .A(G2430), .B(G2443), .ZN(n822) );
  XOR2_X1 U915 ( .A(G2435), .B(KEYINPUT98), .Z(n817) );
  XNOR2_X1 U916 ( .A(G2451), .B(G2438), .ZN(n816) );
  XNOR2_X1 U917 ( .A(n817), .B(n816), .ZN(n818) );
  XOR2_X1 U918 ( .A(n818), .B(G2427), .Z(n820) );
  XNOR2_X1 U919 ( .A(G1341), .B(G1348), .ZN(n819) );
  XNOR2_X1 U920 ( .A(n820), .B(n819), .ZN(n821) );
  XNOR2_X1 U921 ( .A(n822), .B(n821), .ZN(n823) );
  XNOR2_X1 U922 ( .A(n824), .B(n823), .ZN(n825) );
  NAND2_X1 U923 ( .A1(n825), .A2(G14), .ZN(n826) );
  XOR2_X1 U924 ( .A(KEYINPUT99), .B(n826), .Z(n903) );
  XOR2_X1 U925 ( .A(KEYINPUT100), .B(n903), .Z(G401) );
  XNOR2_X1 U926 ( .A(n982), .B(n827), .ZN(n829) );
  XNOR2_X1 U927 ( .A(G171), .B(n981), .ZN(n828) );
  XNOR2_X1 U928 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U929 ( .A(G286), .B(n830), .Z(n831) );
  NOR2_X1 U930 ( .A1(G37), .A2(n831), .ZN(G397) );
  INV_X1 U931 ( .A(n832), .ZN(G319) );
  XOR2_X1 U932 ( .A(G2096), .B(KEYINPUT43), .Z(n834) );
  XNOR2_X1 U933 ( .A(G2090), .B(KEYINPUT102), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U935 ( .A(n835), .B(G2678), .Z(n837) );
  XNOR2_X1 U936 ( .A(G2072), .B(G2067), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U938 ( .A(KEYINPUT42), .B(G2100), .Z(n839) );
  XNOR2_X1 U939 ( .A(G2084), .B(G2078), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(G227) );
  XOR2_X1 U942 ( .A(G1986), .B(G1991), .Z(n843) );
  XNOR2_X1 U943 ( .A(G1966), .B(G1996), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n855) );
  XOR2_X1 U945 ( .A(G1976), .B(G1981), .Z(n845) );
  XNOR2_X1 U946 ( .A(G1956), .B(G1971), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U948 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n847) );
  XNOR2_X1 U949 ( .A(G1961), .B(KEYINPUT41), .ZN(n846) );
  XNOR2_X1 U950 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U952 ( .A(KEYINPUT104), .B(G2474), .Z(n851) );
  XNOR2_X1 U953 ( .A(KEYINPUT103), .B(KEYINPUT105), .ZN(n850) );
  XNOR2_X1 U954 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(G229) );
  NAND2_X1 U957 ( .A1(G112), .A2(n885), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n856), .B(KEYINPUT108), .ZN(n863) );
  NAND2_X1 U959 ( .A1(G136), .A2(n882), .ZN(n858) );
  NAND2_X1 U960 ( .A1(G100), .A2(n588), .ZN(n857) );
  NAND2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n861) );
  NAND2_X1 U962 ( .A1(n886), .A2(G124), .ZN(n859) );
  XOR2_X1 U963 ( .A(KEYINPUT44), .B(n859), .Z(n860) );
  NOR2_X1 U964 ( .A1(n861), .A2(n860), .ZN(n862) );
  NAND2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U966 ( .A(KEYINPUT109), .B(n864), .ZN(G162) );
  XOR2_X1 U967 ( .A(KEYINPUT48), .B(KEYINPUT112), .Z(n866) );
  XNOR2_X1 U968 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n865) );
  XNOR2_X1 U969 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U970 ( .A(G160), .B(n961), .Z(n867) );
  XNOR2_X1 U971 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n871), .B(G162), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n897) );
  NAND2_X1 U975 ( .A1(G118), .A2(n885), .ZN(n875) );
  NAND2_X1 U976 ( .A1(G130), .A2(n886), .ZN(n874) );
  NAND2_X1 U977 ( .A1(n875), .A2(n874), .ZN(n881) );
  NAND2_X1 U978 ( .A1(n882), .A2(G142), .ZN(n876) );
  XNOR2_X1 U979 ( .A(n876), .B(KEYINPUT110), .ZN(n878) );
  NAND2_X1 U980 ( .A1(G106), .A2(n588), .ZN(n877) );
  NAND2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U982 ( .A(KEYINPUT45), .B(n879), .Z(n880) );
  NOR2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n892) );
  NAND2_X1 U984 ( .A1(G139), .A2(n882), .ZN(n884) );
  NAND2_X1 U985 ( .A1(G103), .A2(n588), .ZN(n883) );
  NAND2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G115), .A2(n885), .ZN(n888) );
  NAND2_X1 U988 ( .A1(G127), .A2(n886), .ZN(n887) );
  NAND2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U990 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U991 ( .A1(n891), .A2(n890), .ZN(n954) );
  XOR2_X1 U992 ( .A(n892), .B(n954), .Z(n895) );
  XNOR2_X1 U993 ( .A(G164), .B(n893), .ZN(n894) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U995 ( .A(n897), .B(n896), .Z(n898) );
  NOR2_X1 U996 ( .A1(G37), .A2(n898), .ZN(G395) );
  NOR2_X1 U997 ( .A1(G227), .A2(G229), .ZN(n900) );
  XNOR2_X1 U998 ( .A(KEYINPUT113), .B(KEYINPUT49), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n900), .B(n899), .ZN(n901) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n901), .ZN(n902) );
  NOR2_X1 U1001 ( .A1(G397), .A2(n902), .ZN(n904) );
  NAND2_X1 U1002 ( .A1(n904), .A2(n903), .ZN(n905) );
  NOR2_X1 U1003 ( .A1(n905), .A2(G395), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n906), .B(KEYINPUT114), .ZN(G308) );
  INV_X1 U1005 ( .A(G308), .ZN(G225) );
  INV_X1 U1006 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1007 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n1014) );
  XNOR2_X1 U1008 ( .A(G20), .B(n907), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(G1341), .B(G19), .ZN(n909) );
  XNOR2_X1 U1010 ( .A(G6), .B(G1981), .ZN(n908) );
  NOR2_X1 U1011 ( .A1(n909), .A2(n908), .ZN(n910) );
  NAND2_X1 U1012 ( .A1(n911), .A2(n910), .ZN(n914) );
  XOR2_X1 U1013 ( .A(KEYINPUT59), .B(G1348), .Z(n912) );
  XNOR2_X1 U1014 ( .A(G4), .B(n912), .ZN(n913) );
  NOR2_X1 U1015 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(KEYINPUT124), .B(n915), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(n916), .B(KEYINPUT60), .ZN(n921) );
  XOR2_X1 U1018 ( .A(n917), .B(G5), .Z(n919) );
  XNOR2_X1 U1019 ( .A(G21), .B(G1966), .ZN(n918) );
  NOR2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n929) );
  XNOR2_X1 U1022 ( .A(G1971), .B(G22), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(G23), .B(G1976), .ZN(n922) );
  NOR2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(G1986), .B(KEYINPUT125), .ZN(n924) );
  XNOR2_X1 U1026 ( .A(n924), .B(G24), .ZN(n925) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(KEYINPUT58), .B(n927), .ZN(n928) );
  NOR2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1030 ( .A(KEYINPUT61), .B(n930), .Z(n931) );
  NOR2_X1 U1031 ( .A1(G16), .A2(n931), .ZN(n1012) );
  XNOR2_X1 U1032 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n932) );
  XNOR2_X1 U1033 ( .A(n932), .B(G34), .ZN(n933) );
  XNOR2_X1 U1034 ( .A(G2084), .B(n933), .ZN(n951) );
  XNOR2_X1 U1035 ( .A(G2067), .B(G26), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(G1991), .B(G25), .ZN(n934) );
  NOR2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n941) );
  XOR2_X1 U1038 ( .A(G2072), .B(G33), .Z(n936) );
  NAND2_X1 U1039 ( .A1(n936), .A2(G28), .ZN(n939) );
  XOR2_X1 U1040 ( .A(G32), .B(G1996), .Z(n937) );
  XNOR2_X1 U1041 ( .A(KEYINPUT117), .B(n937), .ZN(n938) );
  NOR2_X1 U1042 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1043 ( .A1(n941), .A2(n940), .ZN(n944) );
  XNOR2_X1 U1044 ( .A(G27), .B(n942), .ZN(n943) );
  NOR2_X1 U1045 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1046 ( .A(n945), .B(KEYINPUT53), .ZN(n946) );
  XNOR2_X1 U1047 ( .A(n946), .B(KEYINPUT118), .ZN(n948) );
  XNOR2_X1 U1048 ( .A(G35), .B(G2090), .ZN(n947) );
  NOR2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1050 ( .A(KEYINPUT119), .B(n949), .ZN(n950) );
  NOR2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1052 ( .A1(G29), .A2(n952), .ZN(n953) );
  XNOR2_X1 U1053 ( .A(n953), .B(KEYINPUT55), .ZN(n980) );
  XOR2_X1 U1054 ( .A(G2072), .B(n954), .Z(n956) );
  XOR2_X1 U1055 ( .A(G164), .B(G2078), .Z(n955) );
  NOR2_X1 U1056 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1057 ( .A(KEYINPUT50), .B(n957), .ZN(n976) );
  XNOR2_X1 U1058 ( .A(G2090), .B(G162), .ZN(n959) );
  NAND2_X1 U1059 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1060 ( .A(n960), .B(KEYINPUT51), .ZN(n971) );
  XNOR2_X1 U1061 ( .A(G160), .B(G2084), .ZN(n964) );
  NOR2_X1 U1062 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1063 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1064 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1065 ( .A(KEYINPUT115), .B(n967), .ZN(n968) );
  NOR2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(KEYINPUT116), .B(n974), .ZN(n975) );
  NAND2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(KEYINPUT52), .B(n977), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(G29), .A2(n978), .ZN(n979) );
  NAND2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n1009) );
  XOR2_X1 U1074 ( .A(G16), .B(KEYINPUT56), .Z(n1006) );
  XNOR2_X1 U1075 ( .A(G171), .B(G1961), .ZN(n993) );
  XNOR2_X1 U1076 ( .A(n981), .B(G1348), .ZN(n984) );
  XOR2_X1 U1077 ( .A(G1341), .B(n982), .Z(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n991) );
  XOR2_X1 U1079 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n989) );
  XOR2_X1 U1080 ( .A(G1966), .B(G168), .Z(n985) );
  XNOR2_X1 U1081 ( .A(KEYINPUT121), .B(n985), .ZN(n986) );
  NAND2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1083 ( .A(n989), .B(n988), .ZN(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n1004) );
  XNOR2_X1 U1086 ( .A(n994), .B(G1956), .ZN(n996) );
  NAND2_X1 U1087 ( .A1(G1971), .A2(G303), .ZN(n995) );
  NAND2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1094 ( .A(KEYINPUT123), .B(n1007), .Z(n1008) );
  NOR2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(G11), .ZN(n1011) );
  NOR2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(n1014), .B(n1013), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(KEYINPUT62), .B(n1015), .ZN(G150) );
  INV_X1 U1100 ( .A(G150), .ZN(G311) );
endmodule

