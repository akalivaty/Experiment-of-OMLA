//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  NAND2_X1  g005(.A1(G229gat), .A2(G233gat), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n207), .B(KEYINPUT13), .Z(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  AND2_X1   g008(.A1(KEYINPUT88), .A2(G29gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(KEYINPUT88), .A2(G29gat), .ZN(new_n211));
  OAI21_X1  g010(.A(G36gat), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT89), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT88), .B(G29gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT89), .A3(G36gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT14), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n214), .A2(new_n216), .A3(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G43gat), .B(G50gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT90), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT15), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226));
  INV_X1    g025(.A(G43gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(G50gat), .ZN(new_n228));
  INV_X1    g027(.A(G50gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(G43gat), .ZN(new_n230));
  OAI211_X1 g029(.A(KEYINPUT90), .B(new_n226), .C1(new_n228), .C2(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT91), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n222), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n214), .A2(new_n216), .A3(new_n221), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n225), .A2(new_n231), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT91), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT92), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n235), .A2(KEYINPUT15), .A3(new_n223), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n239), .B1(new_n238), .B2(new_n240), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G15gat), .B(G22gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT16), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n244), .B1(new_n245), .B2(G1gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(G1gat), .B2(new_n244), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(G8gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n233), .B1(new_n222), .B2(new_n232), .ZN(new_n250));
  NOR3_X1   g049(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT91), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n240), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT92), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n248), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n209), .B1(new_n249), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT17), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n259), .B1(new_n238), .B2(new_n240), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n260), .B1(new_n255), .B2(new_n259), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n207), .B(new_n249), .C1(new_n261), .C2(new_n248), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT18), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n258), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n259), .B1(new_n241), .B2(new_n242), .ZN(new_n265));
  INV_X1    g064(.A(new_n260), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n256), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n268), .A2(KEYINPUT18), .A3(new_n207), .A4(new_n249), .ZN(new_n269));
  AOI211_X1 g068(.A(KEYINPUT87), .B(new_n206), .C1(new_n264), .C2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n206), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n262), .A2(new_n263), .ZN(new_n272));
  INV_X1    g071(.A(new_n258), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT87), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n271), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT27), .B(G183gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G190gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT28), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n279), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n280), .A2(KEYINPUT68), .A3(KEYINPUT28), .A4(new_n282), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT27), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT67), .B1(new_n286), .B2(G183gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n282), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n288), .B1(new_n281), .B2(new_n289), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n284), .B(new_n285), .C1(new_n290), .C2(KEYINPUT28), .ZN(new_n291));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT26), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G169gat), .ZN(new_n296));
  INV_X1    g095(.A(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT69), .B1(new_n298), .B2(KEYINPUT26), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n293), .A2(new_n300), .A3(new_n294), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n295), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(KEYINPUT70), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT70), .ZN(new_n307));
  NOR3_X1   g106(.A1(new_n302), .A2(new_n307), .A3(new_n304), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n291), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT66), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(new_n303), .ZN(new_n312));
  NAND4_X1  g111(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT64), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n312), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n296), .A2(new_n297), .A3(KEYINPUT23), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT23), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n319), .B1(G169gat), .B2(G176gat), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT25), .A4(new_n292), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT65), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n318), .A2(new_n320), .A3(new_n292), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n312), .A2(new_n313), .A3(new_n316), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT65), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .A4(KEYINPUT25), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n314), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT25), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n310), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  AOI211_X1 g130(.A(KEYINPUT66), .B(new_n329), .C1(new_n322), .C2(new_n326), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n309), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT29), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n309), .B(KEYINPUT75), .C1(new_n331), .C2(new_n332), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G226gat), .A2(G233gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT76), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n338), .A2(new_n342), .A3(new_n339), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n330), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n339), .B1(new_n309), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n341), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G197gat), .B(G204gat), .ZN(new_n348));
  AND2_X1   g147(.A1(G211gat), .A2(G218gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n348), .B1(KEYINPUT22), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G211gat), .B(G218gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n337), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(G226gat), .A3(G233gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n309), .A2(new_n344), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n356), .A2(new_n336), .A3(new_n339), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n352), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(G8gat), .B(G36gat), .Z(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT77), .ZN(new_n361));
  XNOR2_X1  g160(.A(G64gat), .B(G92gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n353), .A2(KEYINPUT30), .A3(new_n359), .A4(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n351), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n350), .B(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n345), .B1(new_n340), .B2(KEYINPUT76), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n367), .B1(new_n368), .B2(new_n343), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n363), .B1(new_n369), .B2(new_n358), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n358), .B1(new_n347), .B2(new_n352), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT30), .B1(new_n372), .B2(new_n364), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT5), .ZN(new_n375));
  INV_X1    g174(.A(G113gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(G120gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT72), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(G120gat), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(new_n378), .B2(new_n379), .ZN(new_n381));
  XOR2_X1   g180(.A(G127gat), .B(G134gat), .Z(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(KEYINPUT1), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G120gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(G113gat), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT71), .B1(new_n377), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT1), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n385), .A2(G113gat), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT71), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n379), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n387), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n382), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n384), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(G155gat), .ZN(new_n395));
  INV_X1    g194(.A(G162gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G155gat), .A2(G162gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT78), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n397), .A2(KEYINPUT78), .A3(new_n398), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n398), .A2(KEYINPUT2), .ZN(new_n403));
  OR2_X1    g202(.A1(G141gat), .A2(G148gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(G141gat), .A2(G148gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n401), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n397), .A2(new_n398), .ZN(new_n408));
  XOR2_X1   g207(.A(G141gat), .B(G148gat), .Z(new_n409));
  NAND4_X1  g208(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT78), .A4(new_n403), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n394), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n384), .A3(new_n393), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G225gat), .A2(G233gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n375), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n411), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT3), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n420), .B(new_n394), .C1(new_n421), .C2(new_n411), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n381), .A2(new_n383), .B1(new_n392), .B2(new_n382), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(KEYINPUT4), .A3(new_n411), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n422), .A2(new_n416), .A3(new_n424), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n418), .A2(new_n427), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n424), .A2(new_n426), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n429), .A2(new_n375), .A3(new_n416), .A4(new_n422), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT80), .ZN(new_n432));
  XOR2_X1   g231(.A(G1gat), .B(G29gat), .Z(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G57gat), .B(G85gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT80), .B1(new_n418), .B2(new_n427), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n432), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT6), .ZN(new_n441));
  INV_X1    g240(.A(new_n437), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT80), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n443), .B1(new_n428), .B2(new_n430), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n442), .B1(new_n444), .B2(new_n438), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n440), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT6), .B(new_n442), .C1(new_n444), .C2(new_n438), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT86), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n333), .A2(new_n425), .ZN(new_n450));
  INV_X1    g249(.A(G227gat), .ZN(new_n451));
  INV_X1    g250(.A(G233gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n309), .B(new_n394), .C1(new_n331), .C2(new_n332), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n450), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  XOR2_X1   g254(.A(G71gat), .B(G99gat), .Z(new_n456));
  XNOR2_X1  g255(.A(G15gat), .B(G43gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT33), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n455), .A2(KEYINPUT32), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT73), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n455), .A2(KEYINPUT73), .A3(KEYINPUT32), .A4(new_n459), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n453), .B1(new_n450), .B2(new_n454), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(KEYINPUT34), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n455), .A2(KEYINPUT32), .ZN(new_n467));
  INV_X1    g266(.A(new_n455), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n467), .B(new_n458), .C1(new_n468), .C2(KEYINPUT33), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n464), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n466), .B1(new_n464), .B2(new_n469), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G78gat), .B(G106gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(G22gat), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(G228gat), .A2(G233gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n352), .A2(KEYINPUT29), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT82), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n421), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n367), .A2(new_n336), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(KEYINPUT82), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n412), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n367), .B1(new_n420), .B2(new_n336), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n476), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n419), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n412), .B1(new_n477), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n487), .A2(new_n484), .A3(new_n476), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT31), .B(G50gat), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n485), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n490), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT3), .B1(new_n480), .B2(KEYINPUT82), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n411), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(G228gat), .B(G233gat), .C1(new_n495), .C2(new_n483), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n492), .B1(new_n496), .B2(new_n488), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n475), .B1(new_n491), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n490), .B1(new_n485), .B2(new_n489), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n488), .A3(new_n492), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n474), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n449), .B1(new_n472), .B2(new_n503), .ZN(new_n504));
  NOR4_X1   g303(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT86), .A4(new_n502), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n374), .B(new_n448), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT35), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n472), .A2(new_n503), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT85), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(KEYINPUT35), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n369), .A2(new_n358), .A3(new_n363), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n448), .B1(new_n511), .B2(KEYINPUT30), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n512), .A2(new_n371), .A3(KEYINPUT85), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n510), .B1(new_n513), .B2(KEYINPUT35), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n507), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT83), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n365), .A2(new_n370), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n446), .A2(new_n447), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n353), .A2(new_n359), .A3(new_n364), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT30), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n503), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT74), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(new_n470), .B2(new_n471), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n523), .B(KEYINPUT36), .C1(new_n470), .C2(new_n471), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n516), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n502), .B1(new_n512), .B2(new_n371), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n530), .A2(KEYINPUT83), .A3(new_n526), .A4(new_n527), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n422), .A2(new_n424), .A3(new_n426), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n417), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n533), .B(KEYINPUT84), .Z(new_n534));
  INV_X1    g333(.A(KEYINPUT39), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n442), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n533), .B(KEYINPUT84), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n537), .B(KEYINPUT39), .C1(new_n417), .C2(new_n415), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(KEYINPUT40), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n445), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT40), .B1(new_n536), .B2(new_n538), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n542), .B1(new_n371), .B2(new_n373), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT37), .ZN(new_n544));
  INV_X1    g343(.A(new_n343), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n342), .B1(new_n338), .B2(new_n339), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n545), .A2(new_n546), .A3(new_n345), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n544), .B(new_n359), .C1(new_n547), .C2(new_n367), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n355), .A2(new_n357), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n544), .B1(new_n549), .B2(new_n352), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(new_n547), .B2(new_n352), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT38), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n548), .A2(new_n551), .A3(new_n552), .A4(new_n363), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n448), .B1(new_n372), .B2(new_n364), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n364), .B1(new_n372), .B2(new_n544), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT37), .B1(new_n369), .B2(new_n358), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n552), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n543), .B(new_n503), .C1(new_n555), .C2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n529), .A2(new_n531), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n278), .B1(new_n515), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT9), .ZN(new_n562));
  INV_X1    g361(.A(G71gat), .ZN(new_n563));
  INV_X1    g362(.A(G78gat), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT94), .ZN(new_n566));
  XOR2_X1   g365(.A(G57gat), .B(G64gat), .Z(new_n567));
  INV_X1    g366(.A(KEYINPUT94), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n568), .B(new_n562), .C1(new_n563), .C2(new_n564), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G71gat), .B(G78gat), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n571), .A2(KEYINPUT93), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(KEYINPUT93), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n574), .A2(KEYINPUT95), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n566), .A2(new_n567), .A3(new_n569), .A4(new_n571), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n576), .B1(new_n574), .B2(KEYINPUT95), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT21), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G127gat), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n256), .B1(new_n578), .B2(new_n579), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT96), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n585), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(new_n395), .ZN(new_n590));
  XNOR2_X1  g389(.A(G183gat), .B(G211gat), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n590), .B(new_n591), .Z(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n586), .A2(new_n587), .A3(new_n592), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT101), .ZN(new_n599));
  NAND3_X1  g398(.A1(KEYINPUT98), .A2(G85gat), .A3(G92gat), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT97), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(KEYINPUT7), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G99gat), .A2(G106gat), .ZN(new_n605));
  INV_X1    g404(.A(G85gat), .ZN(new_n606));
  INV_X1    g405(.A(G92gat), .ZN(new_n607));
  AOI22_X1  g406(.A1(KEYINPUT8), .A2(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n604), .B(new_n608), .C1(KEYINPUT7), .C2(new_n602), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT99), .ZN(new_n610));
  XOR2_X1   g409(.A(G99gat), .B(G106gat), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  OR3_X1    g411(.A1(new_n609), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(KEYINPUT99), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n611), .A2(KEYINPUT99), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n609), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n613), .A2(KEYINPUT100), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT100), .B1(new_n613), .B2(new_n616), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n261), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n243), .A2(new_n619), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT41), .ZN(new_n622));
  NAND2_X1  g421(.A1(G232gat), .A2(G233gat), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n599), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n598), .A2(KEYINPUT101), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n623), .A2(new_n622), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n628), .B(new_n629), .Z(new_n630));
  INV_X1    g429(.A(new_n626), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n599), .B(new_n631), .C1(new_n620), .C2(new_n624), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n627), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n630), .B1(new_n627), .B2(new_n632), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G230gat), .A2(G233gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT103), .Z(new_n637));
  NOR2_X1   g436(.A1(new_n575), .A2(new_n577), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n612), .A2(KEYINPUT102), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n609), .B(new_n639), .Z(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT10), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n616), .B(new_n613), .C1(new_n575), .C2(new_n577), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  OAI211_X1 g443(.A(KEYINPUT10), .B(new_n638), .C1(new_n617), .C2(new_n618), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n637), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n641), .A2(new_n643), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n646), .B1(new_n637), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G120gat), .B(G148gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(G176gat), .B(G204gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  OR2_X1    g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n644), .A2(new_n645), .ZN(new_n653));
  INV_X1    g452(.A(new_n637), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n647), .A2(new_n637), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(new_n656), .A3(new_n651), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n596), .A2(new_n635), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n561), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(new_n448), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n661), .B(G1gat), .Z(G1324gat));
  INV_X1    g461(.A(new_n374), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n561), .A2(new_n663), .A3(new_n659), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT16), .B(G8gat), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(KEYINPUT42), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT104), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n664), .A2(G8gat), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n669), .A2(KEYINPUT105), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(KEYINPUT105), .ZN(new_n671));
  AOI22_X1  g470(.A1(new_n670), .A2(new_n671), .B1(KEYINPUT42), .B2(new_n666), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(G1325gat));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n528), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n526), .A2(KEYINPUT106), .A3(new_n527), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G15gat), .B1(new_n660), .B2(new_n678), .ZN(new_n679));
  OR3_X1    g478(.A1(new_n470), .A2(new_n471), .A3(G15gat), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n679), .B1(new_n660), .B2(new_n680), .ZN(G1326gat));
  NOR2_X1   g480(.A1(new_n660), .A2(new_n503), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT43), .B(G22gat), .Z(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  INV_X1    g483(.A(new_n658), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n596), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n635), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT107), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n561), .A2(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n690), .A2(new_n448), .A3(new_n215), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n691), .B(KEYINPUT45), .Z(new_n692));
  NAND2_X1  g491(.A1(new_n635), .A2(KEYINPUT44), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n693), .B1(new_n515), .B2(new_n560), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n559), .A2(new_n530), .A3(new_n675), .A4(new_n676), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n515), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n635), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n694), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n686), .A2(new_n278), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n215), .B1(new_n701), .B2(new_n448), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n692), .A2(new_n702), .ZN(G1328gat));
  NOR3_X1   g502(.A1(new_n690), .A2(G36gat), .A3(new_n374), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT46), .ZN(new_n705));
  OAI21_X1  g504(.A(G36gat), .B1(new_n701), .B2(new_n374), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1329gat));
  AND3_X1   g506(.A1(new_n526), .A2(KEYINPUT106), .A3(new_n527), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT106), .B1(new_n526), .B2(new_n527), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n708), .A2(new_n709), .A3(new_n522), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n710), .A2(new_n559), .B1(new_n507), .B2(new_n514), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n698), .B1(new_n711), .B2(new_n687), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n515), .A2(new_n560), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n713), .A2(KEYINPUT44), .A3(new_n635), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n712), .A2(new_n714), .A3(new_n677), .A4(new_n700), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n699), .A2(KEYINPUT108), .A3(new_n677), .A4(new_n700), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n717), .A2(new_n718), .A3(G43gat), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n561), .A2(new_n227), .A3(new_n472), .A4(new_n689), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT47), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n715), .A2(G43gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n720), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT47), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n723), .A2(new_n724), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n227), .B1(new_n715), .B2(new_n716), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n721), .B1(new_n730), .B2(new_n718), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT47), .B1(new_n725), .B2(new_n720), .ZN(new_n732));
  OAI21_X1  g531(.A(KEYINPUT109), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n729), .A2(new_n733), .ZN(G1330gat));
  NAND4_X1  g533(.A1(new_n712), .A2(new_n714), .A3(new_n502), .A4(new_n700), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G50gat), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n561), .A2(new_n229), .A3(new_n502), .A4(new_n689), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT48), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT110), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n736), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n741), .B1(new_n736), .B2(new_n740), .ZN(new_n744));
  OAI22_X1  g543(.A1(new_n743), .A2(new_n744), .B1(KEYINPUT110), .B2(new_n738), .ZN(new_n745));
  INV_X1    g544(.A(new_n744), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n738), .A2(KEYINPUT110), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n746), .A2(new_n747), .A3(new_n742), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(G1331gat));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750));
  INV_X1    g549(.A(new_n596), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n277), .A2(new_n685), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n751), .A2(new_n752), .A3(new_n687), .ZN(new_n753));
  OR3_X1    g552(.A1(new_n711), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n750), .B1(new_n711), .B2(new_n753), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n518), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g558(.A1(new_n756), .A2(new_n374), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  AND2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n760), .B2(new_n761), .ZN(G1333gat));
  NAND3_X1  g563(.A1(new_n757), .A2(new_n563), .A3(new_n472), .ZN(new_n765));
  OAI21_X1  g564(.A(G71gat), .B1(new_n756), .B2(new_n678), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n765), .A2(KEYINPUT50), .A3(new_n766), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1334gat));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n503), .ZN(new_n772));
  XOR2_X1   g571(.A(KEYINPUT113), .B(G78gat), .Z(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1335gat));
  NAND2_X1  g573(.A1(new_n596), .A2(new_n278), .ZN(new_n775));
  AOI211_X1 g574(.A(new_n687), .B(new_n775), .C1(new_n515), .C2(new_n695), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n685), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n779), .A2(new_n606), .A3(new_n518), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n752), .A2(new_n596), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n699), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(G85gat), .B1(new_n783), .B2(new_n448), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n780), .A2(new_n784), .ZN(G1336gat));
  NAND4_X1  g584(.A1(new_n712), .A2(new_n714), .A3(new_n663), .A4(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G92gat), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n374), .A2(G92gat), .A3(new_n685), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n787), .B(new_n788), .C1(new_n778), .C2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT114), .B1(new_n793), .B2(KEYINPUT51), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n687), .B1(new_n515), .B2(new_n695), .ZN(new_n795));
  INV_X1    g594(.A(new_n775), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT115), .B1(new_n776), .B2(new_n799), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n798), .B(new_n789), .C1(new_n800), .C2(KEYINPUT51), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n787), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n792), .B1(new_n802), .B2(KEYINPUT52), .ZN(new_n803));
  AOI211_X1 g602(.A(KEYINPUT116), .B(new_n788), .C1(new_n801), .C2(new_n787), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n791), .B1(new_n803), .B2(new_n804), .ZN(G1337gat));
  INV_X1    g604(.A(G99gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n779), .A2(new_n806), .A3(new_n472), .ZN(new_n807));
  OAI21_X1  g606(.A(G99gat), .B1(new_n783), .B2(new_n678), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(G1338gat));
  NAND4_X1  g608(.A1(new_n712), .A2(new_n714), .A3(new_n502), .A4(new_n782), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G106gat), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n685), .A2(G106gat), .A3(new_n503), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n811), .B(new_n812), .C1(new_n778), .C2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n696), .A2(new_n799), .A3(new_n635), .A4(new_n796), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n793), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n797), .B1(new_n817), .B2(new_n777), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT117), .B1(new_n818), .B2(new_n813), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT51), .B1(new_n816), .B2(new_n793), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821));
  NOR4_X1   g620(.A1(new_n820), .A2(new_n821), .A3(new_n797), .A4(new_n814), .ZN(new_n822));
  INV_X1    g621(.A(new_n811), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n819), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n815), .B1(new_n824), .B2(new_n812), .ZN(G1339gat));
  NAND3_X1  g624(.A1(new_n644), .A2(new_n645), .A3(new_n637), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n655), .A2(KEYINPUT54), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n651), .B1(new_n646), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n827), .A2(KEYINPUT55), .A3(new_n829), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n832), .A2(new_n657), .A3(new_n833), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n270), .A2(new_n276), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n264), .A2(new_n269), .A3(new_n271), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n207), .B1(new_n268), .B2(new_n249), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n249), .A2(new_n257), .A3(new_n209), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n205), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n658), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n687), .B1(new_n835), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n834), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n635), .A2(new_n836), .A3(new_n839), .A4(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n751), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  NOR4_X1   g643(.A1(new_n596), .A2(new_n635), .A3(new_n277), .A4(new_n658), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n448), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n504), .A2(new_n505), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n847), .A2(new_n374), .A3(new_n848), .ZN(new_n849));
  XOR2_X1   g648(.A(new_n849), .B(KEYINPUT118), .Z(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n376), .A3(new_n277), .ZN(new_n851));
  INV_X1    g650(.A(new_n846), .ZN(new_n852));
  INV_X1    g651(.A(new_n508), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n663), .A2(new_n448), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(G113gat), .B1(new_n855), .B2(new_n278), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n851), .A2(new_n856), .ZN(G1340gat));
  NAND3_X1  g656(.A1(new_n850), .A2(new_n385), .A3(new_n658), .ZN(new_n858));
  OAI21_X1  g657(.A(G120gat), .B1(new_n855), .B2(new_n685), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1341gat));
  OAI21_X1  g659(.A(G127gat), .B1(new_n855), .B2(new_n596), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n596), .A2(G127gat), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n849), .B2(new_n862), .ZN(G1342gat));
  NOR3_X1   g662(.A1(new_n849), .A2(G134gat), .A3(new_n687), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n855), .B2(new_n687), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(G1343gat));
  NOR3_X1   g668(.A1(new_n677), .A2(new_n663), .A3(new_n503), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n847), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(G141gat), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n277), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n878), .B1(new_n835), .B2(new_n840), .ZN(new_n879));
  INV_X1    g678(.A(new_n276), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n274), .A2(new_n275), .A3(new_n271), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(new_n842), .A3(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n840), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n883), .A3(KEYINPUT120), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n879), .A2(new_n687), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n751), .B1(new_n885), .B2(new_n843), .ZN(new_n886));
  OAI211_X1 g685(.A(KEYINPUT57), .B(new_n502), .C1(new_n886), .C2(new_n845), .ZN(new_n887));
  XOR2_X1   g686(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n846), .B2(new_n503), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n678), .A2(new_n854), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n890), .A2(new_n277), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n872), .B1(new_n893), .B2(KEYINPUT121), .ZN(new_n894));
  AOI211_X1 g693(.A(new_n278), .B(new_n891), .C1(new_n887), .C2(new_n889), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n877), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n893), .A2(G141gat), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n876), .B1(new_n899), .B2(new_n875), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT122), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n874), .A2(KEYINPUT58), .ZN(new_n902));
  OAI21_X1  g701(.A(G141gat), .B1(new_n895), .B2(new_n896), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n893), .A2(KEYINPUT121), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n895), .A2(new_n872), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT58), .B1(new_n907), .B2(new_n874), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n901), .A2(new_n909), .ZN(G1344gat));
  NOR2_X1   g709(.A1(new_n886), .A2(new_n845), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n911), .A2(new_n503), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n852), .A2(new_n502), .ZN(new_n913));
  OAI22_X1  g712(.A1(new_n912), .A2(KEYINPUT57), .B1(new_n913), .B2(new_n888), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n658), .A3(new_n892), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n891), .B1(new_n887), .B2(new_n889), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(new_n918), .A3(new_n658), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n871), .A2(new_n685), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(new_n918), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n916), .B(new_n919), .C1(G148gat), .C2(new_n921), .ZN(G1345gat));
  AND2_X1   g721(.A1(new_n917), .A2(new_n751), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n751), .A2(new_n395), .ZN(new_n924));
  OAI22_X1  g723(.A1(new_n923), .A2(new_n395), .B1(new_n871), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT123), .ZN(G1346gat));
  NOR2_X1   g725(.A1(new_n687), .A2(new_n396), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n847), .A2(new_n635), .A3(new_n870), .ZN(new_n928));
  AOI22_X1  g727(.A1(new_n917), .A2(new_n927), .B1(new_n396), .B2(new_n928), .ZN(G1347gat));
  NOR3_X1   g728(.A1(new_n846), .A2(new_n518), .A3(new_n374), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n853), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n931), .A2(new_n296), .A3(new_n278), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n848), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n277), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n932), .B1(new_n296), .B2(new_n935), .ZN(G1348gat));
  NOR3_X1   g735(.A1(new_n931), .A2(new_n297), .A3(new_n685), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n297), .B1(new_n933), .B2(new_n685), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n939), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(G1349gat));
  OAI21_X1  g741(.A(G183gat), .B1(new_n931), .B2(new_n596), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n751), .A2(new_n280), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n933), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g744(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n945), .B(new_n946), .ZN(G1350gat));
  OAI21_X1  g746(.A(G190gat), .B1(new_n931), .B2(new_n687), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT61), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n934), .A2(new_n282), .A3(new_n635), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1351gat));
  INV_X1    g750(.A(G197gat), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n374), .A2(new_n518), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n678), .A2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n914), .A2(new_n277), .A3(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n952), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n958), .B1(new_n957), .B2(new_n956), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n677), .A2(new_n503), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n930), .A2(new_n960), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n961), .A2(G197gat), .A3(new_n278), .ZN(new_n962));
  XOR2_X1   g761(.A(new_n962), .B(KEYINPUT126), .Z(new_n963));
  NAND2_X1  g762(.A1(new_n959), .A2(new_n963), .ZN(G1352gat));
  NOR3_X1   g763(.A1(new_n961), .A2(G204gat), .A3(new_n685), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT62), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n914), .A2(new_n658), .A3(new_n955), .ZN(new_n967));
  INV_X1    g766(.A(G204gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(G1353gat));
  OR3_X1    g768(.A1(new_n961), .A2(G211gat), .A3(new_n596), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n914), .A2(new_n751), .A3(new_n955), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n971), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT63), .B1(new_n971), .B2(G211gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(G1354gat));
  NAND3_X1  g773(.A1(new_n914), .A2(new_n635), .A3(new_n955), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(G218gat), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n687), .A2(G218gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n976), .B1(new_n961), .B2(new_n977), .ZN(G1355gat));
endmodule


