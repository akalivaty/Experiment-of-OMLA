//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT90), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(G8gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  AND2_X1   g005(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G1gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n205), .B(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G29gat), .A2(G36gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G43gat), .B(G50gat), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n215), .A2(KEYINPUT15), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT87), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n214), .A2(KEYINPUT87), .A3(new_n216), .ZN(new_n220));
  XOR2_X1   g019(.A(new_n213), .B(KEYINPUT88), .Z(new_n221));
  AND2_X1   g020(.A1(new_n221), .A2(new_n212), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n215), .A2(KEYINPUT15), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n216), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n219), .A2(new_n220), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n209), .B1(KEYINPUT17), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n219), .A2(new_n220), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n222), .A2(new_n224), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT17), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT89), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT89), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n225), .A2(new_n232), .A3(KEYINPUT17), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n226), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n229), .A2(new_n209), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT18), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n207), .A2(G1gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n205), .B(new_n239), .ZN(new_n240));
  OR3_X1    g039(.A1(new_n240), .A2(new_n225), .A3(KEYINPUT91), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n236), .A2(KEYINPUT91), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT92), .B1(new_n240), .B2(new_n225), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n240), .A2(KEYINPUT92), .A3(new_n225), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n241), .B(new_n242), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n235), .B(KEYINPUT13), .Z(new_n246));
  AOI22_X1  g045(.A1(new_n237), .A2(new_n238), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n234), .A2(KEYINPUT18), .A3(new_n235), .A4(new_n236), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G141gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(G197gat), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT11), .B(G169gat), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n253), .B(KEYINPUT12), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n238), .ZN(new_n256));
  INV_X1    g055(.A(new_n254), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n245), .A2(new_n246), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n256), .A2(new_n257), .A3(new_n248), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G228gat), .ZN(new_n262));
  INV_X1    g061(.A(G233gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT75), .B(G148gat), .Z(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268));
  INV_X1    g067(.A(G155gat), .ZN(new_n269));
  INV_X1    g068(.A(G162gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n268), .B1(new_n271), .B2(KEYINPUT2), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT75), .B(G148gat), .ZN(new_n273));
  INV_X1    g072(.A(G141gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT76), .ZN(new_n276));
  INV_X1    g075(.A(G148gat), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n276), .B1(new_n277), .B2(G141gat), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n267), .B(new_n272), .C1(new_n275), .C2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT3), .ZN(new_n280));
  XNOR2_X1  g079(.A(G141gat), .B(G148gat), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n268), .B(new_n271), .C1(new_n281), .C2(KEYINPUT2), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT29), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n286));
  NAND2_X1  g085(.A1(G211gat), .A2(G218gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(G211gat), .A2(G218gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G211gat), .ZN(new_n292));
  INV_X1    g091(.A(G218gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT72), .B1(new_n294), .B2(new_n287), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n286), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n290), .B1(new_n288), .B2(new_n289), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n294), .A2(KEYINPUT72), .A3(new_n287), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT73), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT22), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n287), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n287), .A2(KEYINPUT71), .A3(new_n300), .ZN(new_n304));
  OR2_X1    g103(.A1(G197gat), .A2(G204gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(G197gat), .A2(G204gat), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n303), .A2(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n296), .A2(new_n299), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n305), .A2(new_n306), .ZN(new_n309));
  INV_X1    g108(.A(new_n304), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT71), .B1(new_n287), .B2(new_n300), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n298), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n312), .A2(new_n286), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n285), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n279), .A2(new_n282), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n308), .A2(new_n284), .A3(new_n314), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT3), .B1(new_n319), .B2(KEYINPUT81), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT81), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n308), .A2(new_n314), .A3(new_n321), .A4(new_n284), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n318), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n316), .B1(new_n323), .B2(KEYINPUT82), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT82), .ZN(new_n325));
  AOI211_X1 g124(.A(new_n325), .B(new_n318), .C1(new_n320), .C2(new_n322), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n265), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G22gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n315), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(new_n284), .A3(new_n317), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n265), .B1(new_n317), .B2(KEYINPUT3), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n327), .A2(new_n328), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n328), .B1(new_n327), .B2(new_n332), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT83), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n319), .A2(KEYINPUT81), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(new_n280), .A3(new_n322), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n317), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n338), .A2(new_n325), .B1(new_n315), .B2(new_n285), .ZN(new_n339));
  INV_X1    g138(.A(new_n326), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n264), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n332), .ZN(new_n342));
  OAI21_X1  g141(.A(G22gat), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT83), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n328), .A3(new_n332), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G78gat), .B(G106gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT31), .B(G50gat), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n347), .B(new_n348), .Z(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n346), .A3(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n343), .A2(new_n344), .A3(new_n345), .A4(new_n349), .ZN(new_n352));
  NAND2_X1  g151(.A1(G227gat), .A2(G233gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT26), .ZN(new_n355));
  NAND2_X1  g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356));
  INV_X1    g155(.A(G169gat), .ZN(new_n357));
  INV_X1    g156(.A(G176gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT26), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(G169gat), .B2(G176gat), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n355), .B(new_n356), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT27), .B(G183gat), .ZN(new_n363));
  INV_X1    g162(.A(G190gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT28), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n363), .A2(KEYINPUT28), .A3(new_n364), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n362), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OR2_X1    g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n370), .A2(KEYINPUT24), .A3(new_n356), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT64), .ZN(new_n372));
  OR2_X1    g171(.A1(new_n356), .A2(KEYINPUT24), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT23), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(G169gat), .B2(G176gat), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n371), .A2(new_n372), .A3(new_n373), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT25), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n359), .B1(KEYINPUT23), .B2(new_n354), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n378), .A2(new_n371), .A3(new_n375), .A4(new_n373), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n371), .A2(new_n375), .A3(new_n373), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n381), .A2(KEYINPUT64), .A3(KEYINPUT25), .A4(new_n378), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n369), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G113gat), .B(G120gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(KEYINPUT1), .ZN(new_n385));
  XNOR2_X1  g184(.A(G127gat), .B(G134gat), .ZN(new_n386));
  OR2_X1    g185(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n386), .B(new_n387), .C1(new_n384), .C2(KEYINPUT1), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n383), .A2(new_n392), .ZN(new_n393));
  AOI211_X1 g192(.A(new_n391), .B(new_n369), .C1(new_n380), .C2(new_n382), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n353), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(KEYINPUT67), .A2(KEYINPUT34), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(KEYINPUT67), .A2(KEYINPUT34), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n382), .ZN(new_n399));
  INV_X1    g198(.A(new_n369), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n391), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n392), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n402), .A2(KEYINPUT68), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n353), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n402), .A2(new_n403), .B1(KEYINPUT68), .B2(KEYINPUT34), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n397), .B(new_n398), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n393), .A2(new_n394), .A3(new_n353), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT32), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT66), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G15gat), .B(G43gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(G71gat), .B(G99gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n402), .A2(G227gat), .A3(G233gat), .A4(new_n403), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT33), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT66), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n414), .A2(new_n417), .A3(KEYINPUT32), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n410), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n414), .B(KEYINPUT32), .C1(new_n415), .C2(new_n413), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n407), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n420), .A3(new_n407), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT69), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT69), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n419), .A2(new_n420), .A3(new_n424), .A4(new_n407), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n421), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n317), .A2(KEYINPUT3), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT77), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n391), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n389), .A2(KEYINPUT77), .A3(new_n390), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n427), .A2(new_n431), .A3(new_n283), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n279), .A2(new_n391), .A3(new_n282), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT4), .ZN(new_n435));
  NAND2_X1  g234(.A1(G225gat), .A2(G233gat), .ZN(new_n436));
  XOR2_X1   g235(.A(new_n436), .B(KEYINPUT78), .Z(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT4), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n432), .A2(new_n435), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  OR2_X1    g240(.A1(new_n441), .A2(KEYINPUT5), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n429), .A2(new_n430), .B1(new_n279), .B2(new_n282), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n437), .B1(new_n443), .B2(new_n434), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT79), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT79), .B(new_n437), .C1(new_n443), .C2(new_n434), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n446), .A2(new_n441), .A3(KEYINPUT5), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(G1gat), .B(G29gat), .Z(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(G57gat), .B(G85gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n456));
  INV_X1    g255(.A(new_n454), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n448), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n455), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n449), .A2(KEYINPUT6), .A3(new_n454), .ZN(new_n460));
  XNOR2_X1  g259(.A(G8gat), .B(G36gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(G64gat), .B(G92gat), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n461), .B(new_n462), .Z(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n401), .A2(KEYINPUT74), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT74), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n383), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n465), .A2(G226gat), .A3(G233gat), .A4(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n401), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n468), .A2(new_n315), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n383), .A2(new_n466), .ZN(new_n472));
  AOI211_X1 g271(.A(KEYINPUT74), .B(new_n369), .C1(new_n380), .C2(new_n382), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n383), .A2(G226gat), .A3(G233gat), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n315), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n464), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n468), .A2(new_n315), .A3(new_n470), .ZN(new_n478));
  INV_X1    g277(.A(new_n475), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n465), .A2(new_n467), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(new_n469), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n478), .B(new_n463), .C1(new_n481), .C2(new_n315), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n477), .A2(KEYINPUT30), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n476), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT30), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n484), .A2(new_n485), .A3(new_n478), .A4(new_n463), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n459), .A2(new_n460), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n351), .A2(new_n352), .A3(new_n426), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT35), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT86), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n488), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n492));
  INV_X1    g291(.A(new_n460), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT84), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n494), .B1(new_n449), .B2(new_n454), .ZN(new_n495));
  AOI211_X1 g294(.A(KEYINPUT84), .B(new_n457), .C1(new_n442), .C2(new_n448), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n458), .A2(new_n456), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n493), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n486), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n499), .A2(KEYINPUT35), .A3(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n351), .A2(new_n352), .ZN(new_n503));
  INV_X1    g302(.A(new_n421), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n423), .A2(new_n425), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT70), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n423), .A2(KEYINPUT70), .A3(new_n425), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n502), .A2(new_n503), .A3(new_n504), .A4(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n491), .A2(new_n492), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n482), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n478), .B1(new_n481), .B2(new_n315), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n464), .B1(new_n513), .B2(KEYINPUT37), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n514), .A2(KEYINPUT38), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n481), .A2(new_n329), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n468), .A2(new_n329), .A3(new_n470), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n516), .A2(KEYINPUT85), .A3(KEYINPUT37), .A4(new_n517), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n517), .B(KEYINPUT37), .C1(new_n481), .C2(new_n329), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT85), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n512), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n513), .A2(KEYINPUT37), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT38), .B1(new_n524), .B2(new_n514), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n499), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n435), .A2(new_n440), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n438), .B1(new_n527), .B2(new_n432), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT39), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n454), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n443), .A2(new_n434), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT39), .B1(new_n531), .B2(new_n437), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n530), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT40), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(new_n501), .A3(new_n497), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n503), .A2(new_n526), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n351), .A2(new_n352), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n459), .A2(new_n460), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n537), .B1(new_n539), .B2(new_n501), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT36), .B1(new_n509), .B2(new_n504), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n426), .A2(KEYINPUT36), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n536), .B(new_n540), .C1(new_n541), .C2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n261), .B1(new_n511), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n546));
  INV_X1    g345(.A(G57gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(G64gat), .ZN(new_n548));
  INV_X1    g347(.A(G64gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(G57gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT93), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n546), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(new_n552), .B2(new_n551), .ZN(new_n554));
  XOR2_X1   g353(.A(G71gat), .B(G78gat), .Z(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n546), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT94), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n548), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n548), .A2(new_n558), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n550), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n557), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n563), .A2(KEYINPUT21), .ZN(new_n564));
  XNOR2_X1  g363(.A(G127gat), .B(G155gat), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n564), .B(new_n565), .Z(new_n566));
  AOI21_X1  g365(.A(new_n209), .B1(KEYINPUT21), .B2(new_n563), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT95), .ZN(new_n570));
  XOR2_X1   g369(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G183gat), .B(G211gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n568), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G232gat), .A2(G233gat), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(KEYINPUT41), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT96), .ZN(new_n580));
  XNOR2_X1  g379(.A(G190gat), .B(G218gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT97), .B(KEYINPUT7), .ZN(new_n584));
  NAND2_X1  g383(.A1(G85gat), .A2(G92gat), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  NAND2_X1  g386(.A1(G99gat), .A2(G106gat), .ZN(new_n588));
  INV_X1    g387(.A(G85gat), .ZN(new_n589));
  INV_X1    g388(.A(G92gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(KEYINPUT8), .A2(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G99gat), .B(G106gat), .Z(new_n593));
  OR2_X1    g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(new_n229), .B2(new_n230), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n232), .B1(new_n225), .B2(KEYINPUT17), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n229), .A2(KEYINPUT89), .A3(new_n230), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n594), .A2(new_n595), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n601), .A2(new_n229), .B1(KEYINPUT41), .B2(new_n578), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT98), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n601), .B1(KEYINPUT17), .B2(new_n225), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n605), .B1(new_n231), .B2(new_n233), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT98), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n606), .A2(new_n607), .A3(new_n602), .ZN(new_n608));
  XNOR2_X1  g407(.A(G134gat), .B(G162gat), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n604), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n610), .B1(new_n604), .B2(new_n608), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n583), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NOR3_X1   g412(.A1(new_n600), .A2(KEYINPUT98), .A3(new_n603), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n607), .B1(new_n606), .B2(new_n602), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n609), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n604), .A2(new_n608), .A3(new_n610), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n582), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n556), .A2(new_n562), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n596), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n563), .A2(new_n594), .A3(new_n595), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n601), .A2(KEYINPUT10), .A3(new_n563), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n621), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n623), .A2(new_n624), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n628), .B1(new_n629), .B2(new_n621), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  OR2_X1    g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n626), .A2(new_n627), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n620), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n629), .A2(new_n621), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(new_n637), .A3(new_n633), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n576), .A2(new_n619), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n545), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n539), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G1gat), .ZN(G1324gat));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n644), .A2(new_n647), .A3(new_n501), .ZN(new_n648));
  OAI21_X1  g447(.A(KEYINPUT99), .B1(new_n643), .B2(new_n500), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(G8gat), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT16), .B(G8gat), .Z(new_n651));
  NAND4_X1  g450(.A1(new_n644), .A2(KEYINPUT42), .A3(new_n501), .A4(new_n651), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n648), .A2(new_n649), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n651), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AOI211_X1 g457(.A(KEYINPUT100), .B(KEYINPUT42), .C1(new_n655), .C2(new_n651), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n653), .B1(new_n658), .B2(new_n659), .ZN(G1325gat));
  NOR2_X1   g459(.A1(new_n541), .A2(new_n543), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n644), .A2(G15gat), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n509), .A2(new_n504), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n643), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(G15gat), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n665), .A2(KEYINPUT101), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(KEYINPUT101), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(G1326gat));
  NOR2_X1   g467(.A1(new_n643), .A2(new_n503), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT43), .B(G22gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  NOR3_X1   g470(.A1(new_n611), .A2(new_n612), .A3(new_n583), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n582), .B1(new_n616), .B2(new_n617), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n576), .A2(new_n639), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n545), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n676), .A2(G29gat), .A3(new_n538), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(KEYINPUT45), .Z(new_n678));
  INV_X1    g477(.A(new_n675), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(new_n261), .ZN(new_n680));
  AND2_X1   g479(.A1(KEYINPUT102), .A2(KEYINPUT44), .ZN(new_n681));
  NOR2_X1   g480(.A1(KEYINPUT102), .A2(KEYINPUT44), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n511), .A2(new_n544), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n684), .B2(new_n674), .ZN(new_n685));
  AOI211_X1 g484(.A(new_n619), .B(new_n681), .C1(new_n511), .C2(new_n544), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n680), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(G29gat), .B1(new_n687), .B2(new_n538), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n678), .A2(new_n688), .ZN(G1328gat));
  NOR3_X1   g488(.A1(new_n676), .A2(G36gat), .A3(new_n500), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT46), .ZN(new_n691));
  OAI21_X1  g490(.A(G36gat), .B1(new_n687), .B2(new_n500), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(G1329gat));
  NAND2_X1  g492(.A1(new_n661), .A2(G43gat), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n676), .A2(new_n663), .ZN(new_n695));
  OAI22_X1  g494(.A1(new_n687), .A2(new_n694), .B1(new_n695), .B2(G43gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g496(.A(KEYINPUT48), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n676), .A2(G50gat), .A3(new_n503), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n537), .B(new_n680), .C1(new_n685), .C2(new_n686), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n699), .B1(new_n700), .B2(G50gat), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n698), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n700), .A2(G50gat), .ZN(new_n704));
  OAI211_X1 g503(.A(KEYINPUT103), .B(KEYINPUT48), .C1(new_n704), .C2(new_n699), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n703), .A2(new_n705), .ZN(G1331gat));
  NOR2_X1   g505(.A1(new_n674), .A2(new_n575), .ZN(new_n707));
  AND4_X1   g506(.A1(new_n261), .A2(new_n684), .A3(new_n707), .A4(new_n639), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n539), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT104), .B(G57gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1332gat));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n500), .B(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n708), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT106), .ZN(new_n717));
  OR2_X1    g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1333gat));
  INV_X1    g518(.A(G71gat), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n708), .B2(new_n661), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n509), .A2(new_n720), .A3(new_n504), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n721), .B1(new_n708), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n537), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g526(.A(new_n619), .B1(new_n511), .B2(new_n544), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n576), .A2(new_n260), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT51), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n684), .A2(KEYINPUT51), .A3(new_n674), .A4(new_n729), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n728), .A2(KEYINPUT108), .A3(KEYINPUT51), .A4(new_n729), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n730), .B1(new_n735), .B2(KEYINPUT109), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n733), .A2(new_n737), .A3(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n539), .A2(new_n589), .A3(new_n639), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n260), .A2(new_n576), .A3(new_n640), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n685), .B2(new_n686), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI211_X1 g544(.A(KEYINPUT107), .B(new_n742), .C1(new_n685), .C2(new_n686), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n745), .A2(new_n539), .A3(new_n746), .ZN(new_n747));
  OAI22_X1  g546(.A1(new_n740), .A2(new_n741), .B1(new_n589), .B2(new_n747), .ZN(G1336gat));
  NAND3_X1  g547(.A1(new_n713), .A2(new_n590), .A3(new_n639), .ZN(new_n749));
  INV_X1    g548(.A(new_n730), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n749), .B1(new_n735), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n745), .A2(new_n501), .A3(new_n746), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n752), .B2(G92gat), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n749), .B1(new_n736), .B2(new_n738), .ZN(new_n755));
  OAI21_X1  g554(.A(G92gat), .B1(new_n743), .B2(new_n714), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n754), .ZN(new_n757));
  OAI22_X1  g556(.A1(new_n753), .A2(new_n754), .B1(new_n755), .B2(new_n757), .ZN(G1337gat));
  NAND3_X1  g557(.A1(new_n745), .A2(new_n661), .A3(new_n746), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT110), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n745), .A2(new_n761), .A3(new_n661), .A4(new_n746), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(G99gat), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n640), .A2(G99gat), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n739), .A2(new_n504), .A3(new_n509), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(G1338gat));
  OR3_X1    g565(.A1(new_n503), .A2(G106gat), .A3(new_n640), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n767), .B1(new_n735), .B2(new_n750), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n745), .A2(new_n537), .A3(new_n746), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n768), .B1(new_n769), .B2(G106gat), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n767), .B1(new_n736), .B2(new_n738), .ZN(new_n772));
  OAI21_X1  g571(.A(G106gat), .B1(new_n743), .B2(new_n503), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n771), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n770), .A2(new_n771), .B1(new_n772), .B2(new_n774), .ZN(G1339gat));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n626), .A2(new_n627), .A3(new_n621), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n636), .A2(KEYINPUT54), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n633), .B1(new_n628), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n778), .A2(KEYINPUT55), .A3(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n781), .A2(new_n638), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n778), .A2(new_n780), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n259), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n257), .B1(new_n247), .B2(new_n248), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n782), .B(new_n785), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n245), .A2(new_n246), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n235), .B1(new_n234), .B2(new_n236), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n253), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n259), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n639), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n674), .B1(new_n788), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n785), .A2(new_n638), .A3(new_n781), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n619), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n776), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n785), .A2(new_n638), .A3(new_n781), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n674), .A2(new_n793), .A3(new_n799), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n799), .A2(new_n260), .B1(new_n793), .B2(new_n639), .ZN(new_n801));
  OAI211_X1 g600(.A(KEYINPUT112), .B(new_n800), .C1(new_n801), .C2(new_n674), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n798), .A2(new_n575), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT111), .B1(new_n641), .B2(new_n260), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n707), .A2(new_n261), .A3(new_n805), .A4(new_n640), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n537), .B1(new_n803), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n713), .A2(new_n538), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n808), .A2(new_n504), .A3(new_n509), .A4(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(G113gat), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n810), .A2(new_n811), .A3(new_n261), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n800), .B1(new_n801), .B2(new_n674), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n576), .B1(new_n813), .B2(new_n776), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n814), .A2(new_n802), .B1(new_n804), .B2(new_n806), .ZN(new_n815));
  INV_X1    g614(.A(new_n426), .ZN(new_n816));
  NOR4_X1   g615(.A1(new_n815), .A2(new_n538), .A3(new_n537), .A4(new_n816), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(new_n714), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n260), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n812), .B1(new_n819), .B2(new_n811), .ZN(G1340gat));
  INV_X1    g619(.A(G120gat), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n810), .A2(new_n821), .A3(new_n640), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n818), .A2(new_n639), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(new_n821), .ZN(G1341gat));
  INV_X1    g623(.A(G127gat), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n818), .A2(new_n825), .A3(new_n576), .ZN(new_n826));
  OAI21_X1  g625(.A(G127gat), .B1(new_n810), .B2(new_n575), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1342gat));
  NOR2_X1   g627(.A1(new_n619), .A2(new_n501), .ZN(new_n829));
  AOI21_X1  g628(.A(G134gat), .B1(KEYINPUT113), .B2(KEYINPUT56), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n817), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(KEYINPUT113), .A2(KEYINPUT56), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n831), .B(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(G134gat), .B1(new_n810), .B2(new_n619), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT114), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(G1343gat));
  NAND2_X1  g635(.A1(new_n803), .A2(new_n807), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n537), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(KEYINPUT57), .ZN(new_n839));
  INV_X1    g638(.A(new_n661), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n813), .A2(new_n575), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n503), .B1(new_n807), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n840), .B(new_n809), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(G141gat), .B1(new_n845), .B2(new_n261), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n661), .A2(new_n503), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n837), .A2(new_n539), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n713), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n260), .A2(new_n274), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT115), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n846), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT58), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n846), .A2(new_n855), .A3(new_n852), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(G1344gat));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n858), .B(new_n273), .C1(new_n845), .C2(new_n640), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n838), .A2(KEYINPUT57), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n841), .B1(new_n260), .B2(new_n641), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(new_n843), .A3(new_n537), .ZN(new_n862));
  NOR4_X1   g661(.A1(new_n661), .A2(new_n538), .A3(new_n640), .A4(new_n713), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(G148gat), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT116), .B1(new_n865), .B2(KEYINPUT59), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n867));
  AOI211_X1 g666(.A(new_n867), .B(new_n858), .C1(new_n864), .C2(G148gat), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n859), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n849), .A2(new_n266), .A3(new_n639), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(G1345gat));
  OAI21_X1  g670(.A(G155gat), .B1(new_n845), .B2(new_n575), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n849), .A2(new_n269), .A3(new_n576), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT117), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n872), .A2(new_n876), .A3(new_n873), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(G1346gat));
  OAI21_X1  g677(.A(G162gat), .B1(new_n845), .B2(new_n619), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n829), .A2(new_n270), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n879), .B1(new_n848), .B2(new_n880), .ZN(G1347gat));
  NAND2_X1  g680(.A1(new_n501), .A2(new_n538), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n663), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n837), .A2(new_n503), .A3(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n808), .A2(KEYINPUT118), .A3(new_n884), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n889), .A2(new_n357), .A3(new_n261), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n815), .A2(new_n539), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n714), .A2(new_n537), .A3(new_n816), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(G169gat), .B1(new_n893), .B2(new_n260), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n890), .A2(new_n894), .ZN(G1348gat));
  OAI21_X1  g694(.A(G176gat), .B1(new_n889), .B2(new_n640), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n893), .A2(new_n358), .A3(new_n639), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1349gat));
  NAND3_X1  g697(.A1(new_n887), .A2(new_n576), .A3(new_n888), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(G183gat), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n576), .A2(new_n363), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n837), .A2(new_n538), .A3(new_n892), .A4(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n904), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n900), .A2(KEYINPUT121), .A3(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT60), .ZN(new_n910));
  AOI22_X1  g709(.A1(new_n899), .A2(G183gat), .B1(new_n905), .B2(new_n906), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT120), .B1(new_n911), .B2(KEYINPUT121), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n913), .B1(new_n911), .B2(KEYINPUT120), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n910), .B1(new_n912), .B2(new_n914), .ZN(G1350gat));
  NAND3_X1  g714(.A1(new_n893), .A2(new_n364), .A3(new_n674), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT122), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n364), .B1(KEYINPUT123), .B2(KEYINPUT61), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n918), .B1(new_n889), .B2(new_n619), .ZN(new_n919));
  NOR2_X1   g718(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n917), .A2(new_n921), .A3(new_n922), .ZN(G1351gat));
  NOR3_X1   g722(.A1(new_n661), .A2(new_n503), .A3(new_n714), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n891), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(KEYINPUT124), .B(G197gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n260), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n661), .A2(new_n882), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n860), .A2(new_n862), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n261), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n927), .B1(new_n930), .B2(new_n926), .ZN(G1352gat));
  OAI21_X1  g730(.A(G204gat), .B1(new_n929), .B2(new_n640), .ZN(new_n932));
  INV_X1    g731(.A(G204gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n925), .A2(new_n933), .A3(new_n639), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n934), .A2(KEYINPUT62), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n934), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT125), .B1(new_n934), .B2(KEYINPUT62), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n932), .B(new_n935), .C1(new_n936), .C2(new_n937), .ZN(G1353gat));
  NAND4_X1  g737(.A1(new_n891), .A2(new_n292), .A3(new_n576), .A4(new_n924), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT126), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n860), .A2(new_n576), .A3(new_n862), .A4(new_n928), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT63), .B1(new_n942), .B2(G211gat), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n940), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(new_n941), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n942), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n944), .A2(new_n947), .ZN(G1354gat));
  OAI21_X1  g747(.A(G218gat), .B1(new_n929), .B2(new_n619), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n925), .A2(new_n293), .A3(new_n674), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1355gat));
endmodule


