//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n444, new_n445, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n554, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  INV_X1    g017(.A(G2072), .ZN(new_n443));
  INV_X1    g018(.A(G2078), .ZN(new_n444));
  NOR2_X1   g019(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g020(.A1(new_n445), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g022(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n463), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n470), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT66), .ZN(G160));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n467), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n473), .A2(G136), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n477), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  AND2_X1   g059(.A1(new_n464), .A2(new_n466), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(new_n477), .ZN(new_n486));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  OAI21_X1  g062(.A(KEYINPUT4), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n473), .A2(new_n489), .A3(G138), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT67), .B(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n478), .A2(G126), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n485), .A2(G126), .A3(G2105), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n492), .B2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT68), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n491), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT5), .B(G543), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT69), .B(G88), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n504), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n509), .A2(G50), .A3(G543), .ZN(new_n513));
  AND3_X1   g088(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n512), .B1(new_n511), .B2(new_n513), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n508), .B1(new_n514), .B2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND3_X1  g092(.A1(new_n504), .A2(new_n509), .A3(G89), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n509), .A2(G51), .A3(G543), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT5), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G543), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n521), .A2(new_n523), .A3(G63), .A4(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT7), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n527), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n518), .A2(new_n519), .A3(new_n524), .A4(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  NAND2_X1  g106(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT6), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G651), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n532), .A2(new_n534), .A3(G52), .A4(G543), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n521), .A2(new_n523), .A3(new_n532), .A4(new_n534), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n521), .A2(new_n523), .A3(G64), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n506), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n521), .A2(new_n523), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G651), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n532), .A2(new_n534), .A3(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G43), .ZN(new_n549));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  OAI211_X1 g125(.A(new_n547), .B(new_n549), .C1(new_n550), .C2(new_n536), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G188));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT71), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT71), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G65), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n559), .B1(new_n544), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n532), .A2(new_n534), .A3(G53), .A4(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n509), .A2(new_n569), .A3(G53), .A4(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n536), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G91), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n566), .A2(new_n571), .A3(new_n573), .ZN(G299));
  NAND2_X1  g149(.A1(new_n539), .A2(new_n540), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G651), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n504), .A2(new_n509), .A3(G90), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n576), .A2(KEYINPUT72), .A3(new_n535), .A4(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT72), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n579), .B1(new_n538), .B2(new_n541), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(G301));
  NAND2_X1  g156(.A1(new_n548), .A2(G49), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n504), .A2(new_n509), .A3(G87), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  NAND2_X1  g160(.A1(new_n548), .A2(G48), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n588));
  OAI221_X1 g163(.A(new_n586), .B1(new_n587), .B2(new_n536), .C1(new_n588), .C2(new_n506), .ZN(G305));
  NAND2_X1  g164(.A1(new_n548), .A2(G47), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n504), .A2(new_n509), .A3(G85), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OAI211_X1 g167(.A(new_n590), .B(new_n591), .C1(new_n592), .C2(new_n506), .ZN(G290));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  OAI21_X1  g169(.A(KEYINPUT10), .B1(new_n536), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n504), .A2(new_n509), .A3(new_n596), .A4(G92), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g173(.A(KEYINPUT74), .B(G66), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n504), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(G54), .B2(new_n548), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT73), .B1(new_n605), .B2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  MUX2_X1   g182(.A(KEYINPUT73), .B(new_n606), .S(new_n607), .Z(G321));
  XNOR2_X1  g183(.A(G321), .B(KEYINPUT75), .ZN(G284));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G299), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G297));
  XOR2_X1   g187(.A(G297), .B(KEYINPUT76), .Z(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n605), .B1(new_n614), .B2(G860), .ZN(G148));
  OAI21_X1  g190(.A(KEYINPUT78), .B1(new_n552), .B2(G868), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n604), .A2(G559), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT77), .ZN(new_n618));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  MUX2_X1   g195(.A(new_n616), .B(KEYINPUT78), .S(new_n620), .Z(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n485), .A2(new_n471), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2100), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n478), .A2(G123), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT80), .ZN(new_n629));
  INV_X1    g204(.A(G135), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n486), .B2(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(G99), .A2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n632), .B(G2104), .C1(G111), .C2(new_n477), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n473), .A2(KEYINPUT80), .A3(G135), .ZN(new_n634));
  AND4_X1   g209(.A1(new_n628), .A2(new_n631), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2096), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n627), .A2(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(G2427), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT82), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT83), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT84), .Z(new_n653));
  INV_X1    g228(.A(G14), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(new_n649), .B2(new_n651), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2067), .B(G2678), .Z(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(KEYINPUT85), .B2(KEYINPUT17), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n662), .B(new_n663), .C1(KEYINPUT85), .C2(KEYINPUT17), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(G2072), .A2(G2078), .ZN(new_n667));
  OAI22_X1  g242(.A1(new_n661), .A2(new_n665), .B1(new_n445), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n669), .B(new_n670), .Z(G227));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n672), .A2(new_n673), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n675), .A2(new_n677), .A3(new_n679), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n682), .B(new_n683), .C1(new_n681), .C2(new_n680), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  INV_X1    g260(.A(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1991), .B(G1996), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1981), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT86), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(G229));
  AND2_X1   g267(.A1(KEYINPUT87), .A2(G29), .ZN(new_n693));
  NOR2_X1   g268(.A1(KEYINPUT87), .A2(G29), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT24), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n697), .A2(G34), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(G34), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI22_X1  g275(.A1(G160), .A2(G29), .B1(new_n696), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G2084), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n696), .A2(G27), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G164), .B2(new_n696), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT99), .B(G2078), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G4), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n605), .B2(new_n707), .ZN(new_n709));
  INV_X1    g284(.A(G1348), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G11), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n713), .A2(KEYINPUT31), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT88), .B(G16), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G19), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n552), .B2(new_n716), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G1341), .ZN(new_n719));
  OR2_X1    g294(.A1(G29), .A2(G33), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n471), .A2(G103), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT25), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n473), .A2(G139), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n485), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n722), .B(new_n723), .C1(new_n477), .C2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n720), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT96), .B(G28), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(G29), .B1(new_n729), .B2(KEYINPUT30), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(KEYINPUT30), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT97), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n727), .A2(new_n443), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n635), .A2(new_n695), .B1(KEYINPUT31), .B2(new_n713), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR4_X1   g310(.A1(new_n712), .A2(new_n714), .A3(new_n719), .A4(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(KEYINPUT28), .B1(new_n696), .B2(G26), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n696), .A2(KEYINPUT28), .A3(G26), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n478), .A2(G128), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n473), .A2(G140), .ZN(new_n741));
  OAI21_X1  g316(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n477), .A2(G116), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n740), .B(new_n741), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT91), .ZN(new_n745));
  AOI211_X1 g320(.A(new_n737), .B(new_n739), .C1(new_n745), .C2(G29), .ZN(new_n746));
  INV_X1    g321(.A(G2067), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G1966), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n707), .A2(G21), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G168), .B2(new_n707), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT95), .Z(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n748), .B1(new_n749), .B2(new_n753), .ZN(new_n754));
  OAI22_X1  g329(.A1(new_n753), .A2(new_n749), .B1(G2084), .B2(new_n701), .ZN(new_n755));
  OAI21_X1  g330(.A(KEYINPUT98), .B1(G5), .B2(G16), .ZN(new_n756));
  OR3_X1    g331(.A1(KEYINPUT98), .A2(G5), .A3(G16), .ZN(new_n757));
  INV_X1    g332(.A(G171), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n756), .B(new_n757), .C1(new_n758), .C2(new_n707), .ZN(new_n759));
  INV_X1    g334(.A(G1961), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n727), .A2(new_n443), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n716), .A2(KEYINPUT23), .A3(G20), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT23), .ZN(new_n764));
  INV_X1    g339(.A(G20), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n715), .B2(new_n765), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n763), .B(new_n766), .C1(new_n611), .C2(new_n707), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1956), .ZN(new_n768));
  NOR4_X1   g343(.A1(new_n755), .A2(new_n761), .A3(new_n762), .A4(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n736), .A2(new_n754), .A3(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n716), .A2(G24), .ZN(new_n772));
  INV_X1    g347(.A(G290), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n716), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(G1986), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(G1986), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n716), .A2(G22), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G166), .B2(new_n716), .ZN(new_n778));
  INV_X1    g353(.A(G1971), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n707), .A2(G23), .ZN(new_n781));
  INV_X1    g356(.A(G288), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n707), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT89), .B(KEYINPUT33), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1976), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n783), .B(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G6), .A2(G16), .ZN(new_n787));
  INV_X1    g362(.A(G305), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(G16), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT32), .B(G1981), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n780), .A2(new_n786), .A3(new_n791), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n775), .B(new_n776), .C1(new_n792), .C2(KEYINPUT34), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n478), .A2(G119), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n473), .A2(G131), .ZN(new_n795));
  OAI21_X1  g370(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n477), .A2(G107), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n794), .B(new_n795), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  MUX2_X1   g373(.A(G25), .B(new_n798), .S(new_n695), .Z(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT35), .B(G1991), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n793), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT90), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT36), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n792), .A2(KEYINPUT34), .ZN(new_n806));
  AND3_X1   g381(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n805), .B1(new_n804), .B2(new_n806), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n702), .B(new_n771), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n726), .A2(G32), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT92), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n477), .A2(G2104), .ZN(new_n812));
  INV_X1    g387(.A(G105), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n471), .A2(KEYINPUT92), .A3(G105), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n473), .A2(G141), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n478), .A2(G129), .ZN(new_n817));
  NAND3_X1  g392(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT26), .Z(new_n819));
  NAND3_X1  g394(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT93), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n810), .B1(new_n825), .B2(new_n726), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT94), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT27), .B(G1996), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n696), .A2(G35), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(G162), .B2(new_n696), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT29), .B(G2090), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n809), .A2(new_n829), .A3(new_n833), .ZN(G311));
  INV_X1    g409(.A(G311), .ZN(G150));
  NAND3_X1  g410(.A1(new_n504), .A2(new_n509), .A3(G93), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n509), .A2(G55), .A3(G543), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n836), .A2(new_n837), .A3(KEYINPUT101), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(KEYINPUT101), .B1(new_n836), .B2(new_n837), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n521), .A2(new_n523), .A3(G67), .ZN(new_n841));
  NAND2_X1  g416(.A1(G80), .A2(G543), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(KEYINPUT100), .B1(new_n843), .B2(G651), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n845));
  AOI211_X1 g420(.A(new_n845), .B(new_n506), .C1(new_n841), .C2(new_n842), .ZN(new_n846));
  OAI22_X1  g421(.A1(new_n839), .A2(new_n840), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(G860), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT37), .Z(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n552), .ZN(new_n850));
  INV_X1    g425(.A(new_n840), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(new_n838), .ZN(new_n852));
  INV_X1    g427(.A(new_n844), .ZN(new_n853));
  INV_X1    g428(.A(new_n846), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n852), .A2(new_n855), .A3(new_n551), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n850), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT39), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n605), .A2(G559), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT38), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n858), .B(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n849), .B1(new_n861), .B2(G860), .ZN(G145));
  AND2_X1   g437(.A1(new_n824), .A2(new_n725), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n824), .A2(new_n725), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n745), .ZN(new_n866));
  INV_X1    g441(.A(new_n745), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n863), .B2(new_n864), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n491), .A2(new_n496), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n866), .A2(new_n491), .A3(new_n496), .A4(new_n868), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n473), .A2(G142), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n477), .A2(G118), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(G130), .B2(new_n478), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n624), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(new_n798), .Z(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n873), .A2(KEYINPUT103), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT103), .B1(new_n873), .B2(new_n881), .ZN(new_n883));
  OAI22_X1  g458(.A1(new_n882), .A2(new_n883), .B1(new_n873), .B2(new_n881), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n483), .B(KEYINPUT102), .Z(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(G160), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(new_n635), .Z(new_n887));
  AOI21_X1  g462(.A(G37), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n873), .A2(KEYINPUT104), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n873), .A2(KEYINPUT104), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n880), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n887), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n891), .B(new_n892), .C1(new_n883), .C2(new_n882), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g470(.A1(new_n847), .A2(new_n619), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n898));
  NAND3_X1  g473(.A1(G299), .A2(new_n598), .A3(new_n603), .ZN(new_n899));
  AOI22_X1  g474(.A1(new_n565), .A2(G651), .B1(new_n572), .B2(G91), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n595), .A2(new_n597), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n548), .A2(G54), .ZN(new_n902));
  INV_X1    g477(.A(new_n601), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(new_n504), .B2(new_n599), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n902), .B1(new_n904), .B2(new_n506), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n900), .B(new_n571), .C1(new_n901), .C2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n898), .B1(new_n899), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT105), .B1(new_n604), .B2(new_n611), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n897), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n899), .A2(new_n906), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT41), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n618), .B(new_n857), .ZN(new_n914));
  MUX2_X1   g489(.A(new_n913), .B(new_n910), .S(new_n914), .Z(new_n915));
  XNOR2_X1  g490(.A(G290), .B(G288), .ZN(new_n916));
  NAND2_X1  g491(.A1(G303), .A2(new_n788), .ZN(new_n917));
  OAI211_X1 g492(.A(G305), .B(new_n508), .C1(new_n515), .C2(new_n514), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n916), .B1(new_n918), .B2(new_n917), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n922), .A2(KEYINPUT42), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n920), .B2(new_n921), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n917), .A2(new_n918), .ZN(new_n926));
  INV_X1    g501(.A(new_n916), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n928), .A2(KEYINPUT106), .A3(new_n919), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n923), .B1(KEYINPUT42), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n915), .B(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n896), .B1(new_n932), .B2(new_n619), .ZN(G295));
  OAI21_X1  g508(.A(new_n896), .B1(new_n932), .B2(new_n619), .ZN(G331));
  NAND2_X1  g509(.A1(G301), .A2(G168), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n758), .B2(G168), .ZN(new_n937));
  NAND3_X1  g512(.A1(G171), .A2(KEYINPUT107), .A3(G286), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n857), .ZN(new_n940));
  AOI21_X1  g515(.A(G286), .B1(new_n578), .B2(new_n580), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n577), .A2(new_n535), .ZN(new_n942));
  AND4_X1   g517(.A1(KEYINPUT107), .A2(new_n942), .A3(G286), .A4(new_n576), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n944), .A2(new_n850), .A3(new_n856), .A4(new_n937), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n940), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n913), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT108), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n913), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n930), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n940), .A2(new_n945), .A3(new_n910), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n951), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n946), .A2(KEYINPUT41), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n957), .A2(new_n911), .B1(new_n925), .B2(new_n929), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n946), .B(KEYINPUT41), .C1(new_n907), .C2(new_n908), .ZN(new_n959));
  AOI21_X1  g534(.A(G37), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n913), .A2(new_n946), .A3(new_n949), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n949), .B1(new_n913), .B2(new_n946), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n953), .B(KEYINPUT109), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n930), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G37), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n968), .A3(new_n956), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n962), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT43), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n956), .A2(new_n960), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n956), .A2(new_n973), .A3(new_n960), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT110), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n971), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n978), .B1(new_n977), .B2(new_n979), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n970), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT112), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT112), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n984), .B(new_n970), .C1(new_n980), .C2(new_n981), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(G397));
  INV_X1    g561(.A(KEYINPUT126), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n988), .B1(new_n502), .B2(new_n989), .ZN(new_n990));
  AOI211_X1 g565(.A(KEYINPUT50), .B(G1384), .C1(new_n491), .C2(new_n496), .ZN(new_n991));
  INV_X1    g566(.A(G40), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n475), .A2(new_n992), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n990), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n987), .B1(new_n994), .B2(G1961), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n502), .A2(new_n989), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT50), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n475), .A2(new_n992), .ZN(new_n998));
  INV_X1    g573(.A(new_n991), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(KEYINPUT126), .A3(new_n760), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n996), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n491), .B2(new_n496), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n993), .B1(new_n1006), .B2(KEYINPUT45), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1007), .A3(new_n444), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT53), .B(new_n998), .C1(new_n1006), .C2(KEYINPUT45), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(G2078), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1006), .A2(KEYINPUT45), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n1003), .A2(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n758), .B1(new_n1002), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1010), .B1(new_n1004), .B2(new_n996), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1008), .A2(new_n1003), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1000), .A2(new_n760), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G301), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1013), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT125), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1017), .A2(KEYINPUT125), .A3(new_n1018), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1002), .A2(G301), .A3(new_n1012), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1021), .B1(new_n1027), .B2(new_n1020), .ZN(new_n1028));
  INV_X1    g603(.A(G1956), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n502), .A2(new_n988), .A3(new_n989), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n998), .B1(new_n1006), .B2(new_n988), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT56), .B(G2072), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1005), .A2(new_n1007), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n1036));
  XNOR2_X1  g611(.A(G299), .B(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1033), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n870), .A2(new_n989), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1039), .A2(G2067), .A3(new_n993), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1040), .B1(new_n1000), .B2(new_n710), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(new_n604), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1037), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1038), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT121), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT121), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1046), .B(new_n1038), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT60), .ZN(new_n1048));
  AOI211_X1 g623(.A(new_n1048), .B(new_n1040), .C1(new_n1000), .C2(new_n710), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1011), .A2(new_n998), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT45), .B1(new_n502), .B2(new_n989), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1050), .A2(new_n1051), .A3(G1996), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT58), .B(G1341), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(new_n1006), .B2(new_n998), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n552), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT122), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(KEYINPUT59), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1049), .A2(new_n604), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n994), .A2(G1348), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1048), .B1(new_n1059), .B2(new_n1040), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1041), .A2(KEYINPUT60), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n605), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1063));
  OR2_X1    g638(.A1(new_n1055), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT123), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(KEYINPUT61), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1038), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1066), .B1(new_n1067), .B2(new_n1043), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1058), .A2(new_n1062), .A3(new_n1064), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1065), .A2(KEYINPUT61), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1043), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n1038), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1072), .B2(new_n1066), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1045), .B(new_n1047), .C1(new_n1069), .C2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n588), .A2(new_n506), .ZN(new_n1075));
  OAI21_X1  g650(.A(G1981), .B1(new_n1075), .B2(KEYINPUT116), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1076), .A2(G305), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(G305), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(KEYINPUT117), .A3(new_n1078), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1079), .A2(KEYINPUT49), .ZN(new_n1080));
  INV_X1    g655(.A(G8), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(new_n1006), .B2(new_n998), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1079), .A2(KEYINPUT49), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n782), .A2(G1976), .ZN(new_n1086));
  INV_X1    g661(.A(G1976), .ZN(new_n1087));
  NAND2_X1  g662(.A1(G288), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1082), .A2(new_n1085), .A3(new_n1086), .A4(new_n1088), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1089), .A2(KEYINPUT115), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1085), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1089), .B1(new_n1091), .B2(KEYINPUT115), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1084), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(G303), .A2(G8), .ZN(new_n1095));
  XOR2_X1   g670(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n1096));
  OR2_X1    g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1000), .A2(G2090), .ZN(new_n1101));
  AOI21_X1  g676(.A(G1971), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1100), .B(G8), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n779), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n993), .B1(new_n1039), .B2(KEYINPUT50), .ZN(new_n1105));
  INV_X1    g680(.A(G2090), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(new_n1030), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1081), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1108), .A2(new_n1100), .A3(KEYINPUT119), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1031), .A2(new_n1032), .A3(G2090), .ZN(new_n1111));
  OAI21_X1  g686(.A(G8), .B1(new_n1111), .B2(new_n1102), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1100), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1110), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1094), .B(new_n1103), .C1(new_n1109), .C2(new_n1114), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n989), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n998), .B1(new_n1006), .B2(KEYINPUT45), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n749), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G2084), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n994), .A2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g697(.A(KEYINPUT120), .B(new_n749), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1120), .A2(new_n1122), .A3(G168), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT51), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1081), .A2(KEYINPUT124), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1125), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1120), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1131), .A2(G8), .A3(G286), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1115), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1028), .A2(new_n1074), .A3(new_n1133), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1131), .A2(G8), .A3(G168), .ZN(new_n1135));
  OAI21_X1  g710(.A(G8), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n1113), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1135), .A2(new_n1094), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT63), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1084), .A2(new_n1087), .A3(new_n782), .ZN(new_n1140));
  NOR2_X1   g715(.A1(G305), .A2(G1981), .ZN(new_n1141));
  XOR2_X1   g716(.A(new_n1141), .B(KEYINPUT118), .Z(new_n1142));
  OAI21_X1  g717(.A(new_n1082), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT119), .B1(new_n1108), .B2(new_n1100), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1112), .A2(new_n1110), .A3(new_n1113), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT63), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1147), .A2(new_n1135), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1093), .B1(new_n1149), .B2(new_n1103), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1144), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1129), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1152), .A2(new_n1132), .A3(new_n1127), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT62), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1115), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1152), .A2(new_n1157), .A3(new_n1132), .A4(new_n1127), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1134), .A2(new_n1151), .A3(new_n1159), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1006), .A2(new_n993), .A3(KEYINPUT45), .ZN(new_n1161));
  INV_X1    g736(.A(G1996), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1163), .A2(new_n824), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n745), .B(G2067), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n825), .A2(new_n1162), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT113), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1161), .B(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1164), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1169), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n798), .B(new_n800), .Z(new_n1172));
  OAI21_X1  g747(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(G290), .B(G1986), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1173), .B1(new_n1161), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1160), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1169), .B1(new_n824), .B2(new_n1165), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1163), .B(KEYINPUT46), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT47), .Z(new_n1180));
  NAND3_X1  g755(.A1(new_n1161), .A2(new_n686), .A3(new_n773), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT48), .Z(new_n1182));
  NOR2_X1   g757(.A1(new_n1173), .A2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n798), .A2(new_n800), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1170), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n867), .A2(new_n747), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1171), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1180), .A2(new_n1183), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1176), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(KEYINPUT127), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1176), .A2(new_n1191), .A3(new_n1188), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1190), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g768(.A(G229), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n656), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g770(.A(new_n1196), .B1(new_n888), .B2(new_n893), .ZN(new_n1197));
  INV_X1    g771(.A(G227), .ZN(new_n1198));
  NAND4_X1  g772(.A1(new_n1197), .A2(G319), .A3(new_n1198), .A4(new_n977), .ZN(G225));
  INV_X1    g773(.A(G225), .ZN(G308));
endmodule


