//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  AND2_X1   g001(.A1(new_n187), .A2(G952), .ZN(new_n188));
  NAND2_X1  g002(.A1(G234), .A2(G237), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(G902), .A3(G953), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT21), .B(G898), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n191), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(G214), .B1(G237), .B2(G902), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G113), .B(G122), .ZN(new_n200));
  INV_X1    g014(.A(G104), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n200), .B(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT75), .ZN(new_n203));
  INV_X1    g017(.A(G140), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G125), .ZN(new_n205));
  INV_X1    g019(.A(G125), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n203), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n208), .A2(KEYINPUT75), .A3(G146), .ZN(new_n212));
  OAI22_X1  g026(.A1(new_n211), .A2(new_n212), .B1(new_n210), .B2(new_n209), .ZN(new_n213));
  NOR2_X1   g027(.A1(G237), .A2(G953), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT88), .ZN(new_n216));
  INV_X1    g030(.A(G143), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n214), .B(G214), .C1(KEYINPUT88), .C2(G143), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT18), .A2(G131), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n220), .A2(KEYINPUT18), .A3(G131), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n213), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT16), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n204), .A3(G125), .ZN(new_n227));
  OAI211_X1 g041(.A(G146), .B(new_n227), .C1(new_n208), .C2(new_n226), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT19), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT19), .B1(new_n205), .B2(new_n207), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g045(.A(KEYINPUT65), .B(G131), .Z(new_n232));
  AND3_X1   g046(.A1(new_n218), .A2(new_n232), .A3(new_n219), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(new_n218), .B2(new_n219), .ZN(new_n234));
  OAI221_X1 g048(.A(new_n228), .B1(new_n231), .B2(G146), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n202), .B1(new_n225), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n234), .A2(KEYINPUT17), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n227), .B1(new_n208), .B2(new_n226), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n210), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n228), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  OR3_X1    g055(.A1(new_n233), .A2(new_n234), .A3(KEYINPUT17), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n220), .B(new_n222), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n241), .A2(new_n242), .B1(new_n213), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n236), .B1(new_n244), .B2(new_n202), .ZN(new_n245));
  NOR2_X1   g059(.A1(G475), .A2(G902), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT20), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT20), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n241), .A2(new_n242), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n250), .A2(new_n202), .A3(new_n225), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n249), .B(new_n246), .C1(new_n251), .C2(new_n236), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n217), .A2(G128), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT13), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(KEYINPUT90), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G128), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G143), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n256), .B(new_n258), .C1(new_n255), .C2(new_n254), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT90), .B1(new_n254), .B2(new_n255), .ZN(new_n260));
  OAI21_X1  g074(.A(G134), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n254), .A2(new_n258), .ZN(new_n262));
  INV_X1    g076(.A(G134), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G122), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G116), .ZN(new_n266));
  INV_X1    g080(.A(G116), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G122), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT89), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n266), .A2(new_n268), .A3(KEYINPUT89), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G107), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(G107), .B1(new_n271), .B2(new_n272), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n261), .B(new_n264), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n276), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n262), .B(new_n263), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n267), .A2(KEYINPUT14), .A3(G122), .ZN(new_n280));
  OAI211_X1 g094(.A(G107), .B(new_n280), .C1(new_n269), .C2(KEYINPUT14), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g097(.A(KEYINPUT71), .B(G217), .Z(new_n284));
  XOR2_X1   g098(.A(KEYINPUT9), .B(G234), .Z(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n187), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n286), .B(KEYINPUT91), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT92), .ZN(new_n289));
  INV_X1    g103(.A(new_n287), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(new_n277), .A3(new_n282), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n288), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n283), .A2(KEYINPUT92), .A3(new_n287), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G478), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(KEYINPUT15), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n297), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n292), .A2(new_n293), .A3(new_n294), .A4(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n202), .B1(new_n250), .B2(new_n225), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n293), .B1(new_n251), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G475), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n253), .A2(new_n298), .A3(new_n300), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n210), .A2(G143), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n217), .A2(G146), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT0), .A4(G128), .ZN(new_n307));
  XNOR2_X1  g121(.A(G143), .B(G146), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT0), .B(G128), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G125), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT1), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n308), .A2(new_n313), .A3(G128), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT67), .ZN(new_n315));
  AOI21_X1  g129(.A(G128), .B1(new_n305), .B2(new_n306), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n313), .A2(new_n210), .A3(G143), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n210), .A2(G143), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT1), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n320), .B(KEYINPUT67), .C1(new_n308), .C2(G128), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n314), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n312), .B1(new_n322), .B2(G125), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n187), .A2(G224), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT79), .B(G104), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(new_n274), .ZN(new_n328));
  OR2_X1    g142(.A1(KEYINPUT79), .A2(G104), .ZN(new_n329));
  NAND2_X1  g143(.A1(KEYINPUT79), .A2(G104), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(G107), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n326), .A2(new_n274), .A3(G104), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(G101), .B1(new_n328), .B2(new_n333), .ZN(new_n334));
  AND2_X1   g148(.A1(KEYINPUT79), .A2(G104), .ZN(new_n335));
  NOR2_X1   g149(.A1(KEYINPUT79), .A2(G104), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n274), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT3), .ZN(new_n338));
  INV_X1    g152(.A(G101), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n338), .A2(new_n339), .A3(new_n331), .A4(new_n332), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n334), .A2(KEYINPUT4), .A3(new_n340), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT2), .B(G113), .Z(new_n342));
  XNOR2_X1  g156(.A(G116), .B(G119), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n342), .B(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n345), .B(G101), .C1(new_n328), .C2(new_n333), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n341), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n201), .A2(G107), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n339), .B1(new_n337), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n343), .A2(KEYINPUT5), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n267), .A2(KEYINPUT5), .A3(G119), .ZN(new_n352));
  INV_X1    g166(.A(G113), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n351), .A2(new_n354), .B1(new_n342), .B2(new_n343), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n340), .A2(new_n350), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(G110), .B(G122), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n347), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n347), .A2(new_n357), .ZN(new_n360));
  XOR2_X1   g174(.A(new_n358), .B(KEYINPUT83), .Z(new_n361));
  AOI22_X1  g175(.A1(new_n359), .A2(KEYINPUT6), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n360), .A2(KEYINPUT6), .A3(new_n361), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n325), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n308), .A2(new_n313), .A3(G128), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n217), .A2(G146), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n257), .B1(new_n366), .B2(new_n319), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT67), .B1(new_n367), .B2(new_n320), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n316), .A2(new_n315), .A3(new_n317), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n365), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n206), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n324), .A2(KEYINPUT7), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n312), .A4(new_n373), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n312), .B(new_n373), .C1(new_n322), .C2(G125), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT85), .ZN(new_n376));
  INV_X1    g190(.A(new_n373), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n323), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT84), .B(KEYINPUT8), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n358), .B(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n355), .B1(new_n340), .B2(new_n350), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n380), .B1(new_n356), .B2(new_n381), .ZN(new_n382));
  AND4_X1   g196(.A1(new_n374), .A2(new_n376), .A3(new_n378), .A4(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(G902), .B1(new_n383), .B2(new_n359), .ZN(new_n384));
  OAI21_X1  g198(.A(G210), .B1(G237), .B2(G902), .ZN(new_n385));
  XOR2_X1   g199(.A(new_n385), .B(KEYINPUT86), .Z(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n364), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n364), .A2(new_n384), .ZN(new_n390));
  XOR2_X1   g204(.A(new_n386), .B(KEYINPUT87), .Z(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  AOI211_X1 g207(.A(new_n199), .B(new_n304), .C1(new_n389), .C2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n365), .A2(new_n367), .A3(new_n320), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n340), .A2(new_n350), .A3(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n328), .A2(new_n333), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n349), .B1(new_n397), .B2(new_n339), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n396), .B1(new_n398), .B2(new_n370), .ZN(new_n399));
  INV_X1    g213(.A(G137), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT66), .B1(new_n400), .B2(G134), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT66), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(new_n263), .A3(G137), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(G134), .ZN(new_n404));
  NOR2_X1   g218(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n401), .A2(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n263), .B2(G137), .ZN(new_n408));
  INV_X1    g222(.A(new_n405), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n406), .A2(new_n410), .A3(new_n232), .ZN(new_n411));
  INV_X1    g225(.A(G131), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n406), .B2(new_n410), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n399), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT12), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(KEYINPUT80), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT80), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n340), .A2(new_n350), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n322), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n414), .B1(new_n421), .B2(new_n396), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n419), .B1(new_n422), .B2(KEYINPUT12), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(KEYINPUT12), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n418), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n341), .A2(new_n311), .A3(new_n346), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n370), .A2(KEYINPUT10), .A3(new_n340), .A4(new_n350), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT10), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n396), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n426), .A2(new_n427), .A3(new_n414), .A4(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(G110), .B(G140), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT78), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n187), .A2(G227), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n432), .B(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT81), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n430), .A2(KEYINPUT81), .A3(new_n434), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n425), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT82), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n425), .A2(new_n437), .A3(KEYINPUT82), .A4(new_n438), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n415), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n444), .A2(new_n430), .ZN(new_n445));
  OR2_X1    g259(.A1(new_n445), .A2(new_n434), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n441), .A2(new_n442), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G469), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n448), .A3(new_n293), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n448), .A2(new_n293), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n434), .B1(new_n425), .B2(new_n430), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n435), .B1(new_n415), .B2(new_n443), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G469), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n449), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G221), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(new_n285), .B2(new_n293), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n394), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT22), .B(G137), .ZN(new_n461));
  INV_X1    g275(.A(G234), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n457), .A2(new_n462), .A3(G953), .ZN(new_n463));
  XOR2_X1   g277(.A(new_n461), .B(new_n463), .Z(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n257), .A2(KEYINPUT23), .A3(G119), .ZN(new_n466));
  INV_X1    g280(.A(G119), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G128), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n468), .A2(KEYINPUT23), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n257), .A2(G119), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n466), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G110), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT24), .B(G110), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n468), .B(KEYINPUT73), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT72), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n470), .B(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n240), .B(new_n473), .C1(new_n474), .C2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n228), .B1(new_n211), .B2(new_n212), .ZN(new_n480));
  INV_X1    g294(.A(G110), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n481), .B(new_n466), .C1(new_n469), .C2(new_n471), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n474), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n475), .B2(new_n477), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT74), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n478), .A2(new_n474), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT74), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n480), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n479), .B1(new_n490), .B2(KEYINPUT76), .ZN(new_n491));
  INV_X1    g305(.A(new_n480), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n478), .A2(new_n486), .A3(new_n474), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n482), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n485), .A2(new_n486), .ZN(new_n495));
  OAI211_X1 g309(.A(KEYINPUT76), .B(new_n492), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n465), .B1(new_n491), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT76), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n501), .A2(new_n496), .A3(new_n479), .A4(new_n464), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n284), .B1(new_n462), .B2(G902), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n505), .A2(G902), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n498), .A2(new_n293), .A3(new_n502), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT25), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n508), .B1(new_n511), .B2(new_n505), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT70), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT68), .ZN(new_n514));
  INV_X1    g328(.A(new_n344), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n401), .A2(new_n403), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n404), .A2(new_n405), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n410), .A2(new_n232), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n404), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n400), .A2(G134), .ZN(new_n520));
  OAI21_X1  g334(.A(G131), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n322), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n516), .A2(new_n517), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n405), .B1(new_n404), .B2(new_n407), .ZN(new_n525));
  OAI21_X1  g339(.A(G131), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n310), .B1(new_n526), .B2(new_n518), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT30), .B1(new_n523), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n311), .B1(new_n411), .B2(new_n413), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n529), .B(new_n530), .C1(new_n322), .C2(new_n522), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n515), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n214), .A2(G210), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(KEYINPUT27), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT26), .B(G101), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n534), .B(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n523), .A2(new_n527), .A3(new_n344), .ZN(new_n538));
  NOR4_X1   g352(.A1(new_n532), .A2(KEYINPUT31), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n344), .B1(new_n523), .B2(new_n527), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n529), .B(new_n515), .C1(new_n322), .C2(new_n522), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT28), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT28), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT31), .B1(new_n547), .B2(new_n537), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n532), .A2(new_n537), .A3(new_n538), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n514), .B(new_n540), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n545), .B1(new_n541), .B2(new_n542), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n523), .A2(new_n527), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT28), .B1(new_n552), .B2(new_n515), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n537), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT31), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n528), .A2(new_n531), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n538), .B1(new_n556), .B2(new_n344), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n554), .A2(new_n555), .B1(new_n557), .B2(new_n536), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT68), .B1(new_n558), .B2(new_n539), .ZN(new_n559));
  NOR2_X1   g373(.A1(G472), .A2(G902), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n550), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT32), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT32), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n550), .A2(new_n559), .A3(new_n563), .A4(new_n560), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G472), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n544), .A2(new_n536), .A3(new_n546), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n537), .B1(new_n532), .B2(new_n538), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT29), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n570), .A2(KEYINPUT69), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n544), .A2(KEYINPUT29), .A3(new_n536), .A4(new_n546), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n293), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(KEYINPUT69), .B2(new_n570), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n566), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n513), .B1(new_n565), .B2(new_n576), .ZN(new_n577));
  AOI211_X1 g391(.A(KEYINPUT70), .B(new_n575), .C1(new_n562), .C2(new_n564), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n512), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT77), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g395(.A(KEYINPUT77), .B(new_n512), .C1(new_n577), .C2(new_n578), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n460), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(new_n339), .ZN(G3));
  NAND2_X1  g398(.A1(new_n456), .A2(new_n459), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n550), .A2(new_n559), .A3(new_n293), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(G472), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(new_n561), .A3(new_n512), .ZN(new_n588));
  OR2_X1    g402(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n248), .A2(new_n252), .B1(new_n302), .B2(G475), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n292), .A2(new_n591), .A3(new_n294), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT93), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n288), .A2(KEYINPUT94), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n291), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n290), .A2(new_n277), .A3(KEYINPUT94), .A4(new_n282), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(KEYINPUT33), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT93), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n292), .A2(new_n598), .A3(new_n591), .A4(new_n294), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n296), .A2(G902), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n593), .A2(new_n597), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n295), .A2(new_n296), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n590), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n195), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n387), .B1(new_n364), .B2(new_n384), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n196), .B(new_n605), .C1(new_n388), .C2(new_n606), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n589), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT34), .B(G104), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G6));
  NAND2_X1  g424(.A1(new_n298), .A2(new_n300), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n590), .A2(new_n611), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n589), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT35), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT95), .B(G107), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  AND2_X1   g430(.A1(new_n509), .A2(new_n510), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n509), .A2(new_n510), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n505), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n491), .A2(new_n497), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n465), .A2(KEYINPUT36), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT96), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n620), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n506), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n587), .A2(new_n561), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n460), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT97), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT37), .B(G110), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G12));
  INV_X1    g444(.A(new_n625), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n196), .B1(new_n388), .B2(new_n606), .ZN(new_n632));
  INV_X1    g446(.A(G900), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n191), .B1(new_n193), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n612), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n631), .A2(new_n632), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n585), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n637), .B(new_n638), .C1(new_n577), .C2(new_n578), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G128), .ZN(G30));
  NAND2_X1  g454(.A1(new_n389), .A2(new_n393), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n641), .B(KEYINPUT38), .Z(new_n642));
  INV_X1    g456(.A(new_n590), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n611), .ZN(new_n644));
  NOR4_X1   g458(.A1(new_n642), .A2(new_n197), .A3(new_n625), .A4(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n557), .A2(new_n537), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n293), .B1(new_n543), .B2(new_n536), .ZN(new_n647));
  OAI21_X1  g461(.A(G472), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n565), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n634), .B(KEYINPUT39), .Z(new_n650));
  NAND2_X1  g464(.A1(new_n638), .A2(new_n650), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n645), .B(new_n649), .C1(KEYINPUT40), .C2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(KEYINPUT40), .B2(new_n651), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(new_n217), .ZN(G45));
  INV_X1    g468(.A(new_n634), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n603), .A2(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n631), .A2(new_n632), .A3(new_n656), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n638), .B(new_n657), .C1(new_n577), .C2(new_n578), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G146), .ZN(G48));
  NOR2_X1   g473(.A1(new_n604), .A2(new_n607), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n448), .A2(KEYINPUT98), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n447), .A2(new_n293), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n447), .A2(new_n293), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n661), .ZN(new_n665));
  AND4_X1   g479(.A1(new_n459), .A2(new_n660), .A3(new_n663), .A4(new_n665), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n666), .B(new_n512), .C1(new_n577), .C2(new_n578), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT99), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT41), .B(G113), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G15));
  NOR2_X1   g484(.A1(new_n577), .A2(new_n578), .ZN(new_n671));
  INV_X1    g485(.A(new_n663), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n662), .B1(new_n447), .B2(new_n293), .ZN(new_n673));
  NOR4_X1   g487(.A1(new_n672), .A2(new_n673), .A3(new_n458), .A4(new_n632), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n619), .B1(new_n503), .B2(new_n507), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n677), .A2(new_n195), .A3(new_n612), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G116), .ZN(G18));
  AOI211_X1 g494(.A(new_n304), .B(new_n195), .C1(new_n619), .C2(new_n624), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G119), .ZN(G21));
  NOR2_X1   g497(.A1(new_n607), .A2(new_n644), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n684), .A2(new_n665), .A3(new_n459), .A4(new_n663), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT100), .B(G472), .Z(new_n686));
  NAND2_X1  g500(.A1(new_n586), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n560), .B1(new_n558), .B2(new_n539), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(new_n688), .A3(new_n512), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n265), .ZN(G24));
  INV_X1    g505(.A(new_n656), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n687), .A2(new_n625), .A3(new_n688), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n674), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G125), .ZN(G27));
  AOI21_X1  g509(.A(new_n575), .B1(new_n565), .B2(KEYINPUT102), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n562), .A2(new_n697), .A3(new_n564), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n677), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n452), .A2(KEYINPUT101), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n453), .B1(new_n452), .B2(KEYINPUT101), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(G469), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n449), .A2(new_n702), .A3(new_n451), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n389), .A2(new_n393), .A3(new_n196), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n703), .A2(new_n459), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT42), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n706), .A2(new_n707), .A3(new_n656), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n699), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT103), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n703), .A2(new_n459), .A3(new_n705), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n711), .B(new_n512), .C1(new_n577), .C2(new_n578), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n707), .B1(new_n712), .B2(new_n656), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT103), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n699), .A2(new_n714), .A3(new_n708), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n710), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G131), .ZN(G33));
  NOR2_X1   g531(.A1(new_n712), .A2(new_n636), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n263), .ZN(G36));
  AOI21_X1  g533(.A(new_n643), .B1(new_n601), .B2(new_n602), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n724));
  OAI21_X1  g538(.A(new_n723), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n631), .B1(new_n561), .B2(new_n587), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT44), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n725), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g545(.A(new_n704), .B(KEYINPUT106), .Z(new_n732));
  AND3_X1   g546(.A1(new_n731), .A2(KEYINPUT107), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT107), .B1(new_n731), .B2(new_n732), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n454), .A2(KEYINPUT45), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n448), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n700), .A2(KEYINPUT45), .A3(new_n701), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n450), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n739), .A2(KEYINPUT46), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n449), .B1(new_n739), .B2(KEYINPUT46), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n459), .B(new_n650), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(new_n742), .B(KEYINPUT104), .Z(new_n743));
  NAND2_X1  g557(.A1(new_n735), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G137), .ZN(G39));
  OAI21_X1  g559(.A(new_n459), .B1(new_n740), .B2(new_n741), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n747), .A2(KEYINPUT108), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(KEYINPUT108), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n746), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n750), .B1(new_n746), .B2(new_n749), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n671), .A2(new_n677), .A3(new_n692), .A4(new_n705), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n204), .ZN(G42));
  NOR2_X1   g568(.A1(new_n672), .A2(new_n673), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n755), .B(KEYINPUT49), .Z(new_n756));
  INV_X1    g570(.A(new_n642), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n512), .A2(new_n459), .A3(new_n196), .A4(new_n720), .ZN(new_n758));
  OR4_X1    g572(.A1(new_n649), .A2(new_n756), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT99), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n667), .B(new_n760), .ZN(new_n761));
  OAI221_X1 g575(.A(new_n674), .B1(new_n678), .B2(new_n681), .C1(new_n577), .C2(new_n578), .ZN(new_n762));
  OAI22_X1  g576(.A1(new_n460), .A2(new_n626), .B1(new_n685), .B2(new_n689), .ZN(new_n763));
  INV_X1    g577(.A(new_n612), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n641), .B(new_n198), .C1(new_n603), .C2(new_n764), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n585), .A2(new_n588), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n761), .A2(new_n583), .A3(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n304), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n705), .A2(KEYINPUT109), .A3(new_n770), .A4(new_n655), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n655), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n772), .B1(new_n773), .B2(new_n704), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n631), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n775), .B(new_n638), .C1(new_n578), .C2(new_n577), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n711), .A2(new_n692), .A3(new_n693), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n776), .B(new_n777), .C1(new_n712), .C2(new_n636), .ZN(new_n778));
  INV_X1    g592(.A(new_n715), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n714), .B1(new_n699), .B2(new_n708), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n778), .B1(new_n781), .B2(new_n713), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n632), .A2(new_n644), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n784), .A2(new_n625), .A3(new_n634), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(new_n649), .A3(new_n459), .A4(new_n703), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n639), .A2(new_n658), .A3(new_n694), .A4(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n787), .A2(new_n783), .A3(new_n788), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n769), .B(new_n782), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n581), .A2(new_n582), .ZN(new_n796));
  INV_X1    g610(.A(new_n460), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n768), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n778), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n668), .A3(new_n716), .A4(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n787), .B(KEYINPUT52), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n800), .A2(new_n794), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT54), .B1(new_n795), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n794), .B1(new_n800), .B2(new_n801), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n804), .B1(new_n793), .B2(new_n794), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n803), .B1(KEYINPUT54), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT111), .B1(new_n725), .B2(new_n191), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n725), .A2(KEYINPUT111), .A3(new_n191), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n689), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n757), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n755), .A2(new_n459), .A3(new_n197), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT113), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT114), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n816), .A2(KEYINPUT50), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(KEYINPUT50), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n755), .A2(new_n459), .A3(new_n705), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n808), .B2(new_n809), .ZN(new_n820));
  NOR4_X1   g634(.A1(new_n819), .A2(new_n649), .A3(new_n677), .A4(new_n190), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n601), .A2(new_n590), .A3(new_n602), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n820), .A2(new_n693), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n817), .A2(new_n818), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n812), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n751), .A2(KEYINPUT112), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n755), .A2(new_n458), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n829), .B1(new_n751), .B2(KEYINPUT112), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n732), .B(new_n827), .C1(new_n828), .C2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT51), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n821), .A2(new_n603), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n188), .B(new_n833), .C1(new_n812), .C2(new_n675), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n820), .A2(new_n699), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n835), .A2(KEYINPUT48), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(KEYINPUT48), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n834), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n751), .A2(new_n829), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n827), .A2(KEYINPUT51), .A3(new_n732), .ZN(new_n840));
  OAI22_X1  g654(.A1(new_n839), .A2(new_n840), .B1(KEYINPUT115), .B2(KEYINPUT51), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n838), .B1(new_n824), .B2(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n806), .A2(new_n832), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(G952), .A2(G953), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n759), .B1(new_n843), .B2(new_n844), .ZN(G75));
  NOR2_X1   g659(.A1(new_n187), .A2(G952), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n805), .A2(G902), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT56), .B1(new_n848), .B2(new_n386), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n362), .A2(new_n363), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(new_n325), .ZN(new_n851));
  XOR2_X1   g665(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n852));
  XNOR2_X1  g666(.A(new_n851), .B(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n847), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT56), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n805), .A2(new_n857), .A3(G902), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n857), .B1(new_n805), .B2(G902), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n858), .A2(new_n859), .A3(new_n391), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n856), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n805), .A2(G902), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT117), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n805), .A2(new_n857), .A3(G902), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n392), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT118), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n854), .B1(new_n862), .B2(new_n867), .ZN(G51));
  XNOR2_X1  g682(.A(new_n805), .B(KEYINPUT54), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n450), .B(KEYINPUT57), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n447), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n864), .A2(new_n738), .A3(new_n737), .A4(new_n865), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n846), .B1(new_n872), .B2(new_n873), .ZN(G54));
  AND2_X1   g688(.A1(KEYINPUT58), .A2(G475), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n864), .A2(new_n865), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n245), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n847), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n876), .A2(new_n245), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(G60));
  AND3_X1   g694(.A1(new_n593), .A2(new_n599), .A3(new_n597), .ZN(new_n881));
  NAND2_X1  g695(.A1(G478), .A2(G902), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT59), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n869), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n881), .B1(new_n806), .B2(new_n883), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n884), .A2(new_n885), .A3(new_n846), .ZN(G63));
  NAND2_X1  g700(.A1(G217), .A2(G902), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT119), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT60), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n805), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n846), .B1(new_n890), .B2(new_n503), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n623), .B(KEYINPUT120), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n891), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n893), .B(new_n894), .ZN(G66));
  INV_X1    g709(.A(G224), .ZN(new_n896));
  OAI21_X1  g710(.A(G953), .B1(new_n194), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(new_n769), .B2(G953), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n850), .B1(G898), .B2(new_n187), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT121), .Z(new_n900));
  XNOR2_X1  g714(.A(new_n898), .B(new_n900), .ZN(G69));
  XNOR2_X1  g715(.A(new_n556), .B(KEYINPUT122), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n231), .ZN(new_n903));
  NAND2_X1  g717(.A1(G900), .A2(G953), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n677), .B(new_n784), .C1(new_n696), .C2(new_n698), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n743), .B1(new_n735), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n639), .A2(new_n658), .A3(new_n694), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n753), .A2(new_n718), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n906), .A2(new_n716), .A3(new_n908), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n903), .B(new_n904), .C1(new_n909), .C2(G953), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n911), .A2(KEYINPUT123), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(KEYINPUT123), .ZN(new_n913));
  OR4_X1    g727(.A1(new_n653), .A2(new_n907), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  OAI211_X1 g728(.A(KEYINPUT123), .B(new_n911), .C1(new_n653), .C2(new_n907), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n753), .B1(new_n735), .B2(new_n743), .ZN(new_n918));
  AOI211_X1 g732(.A(new_n704), .B(new_n651), .C1(new_n604), .C2(new_n612), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n796), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT124), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT125), .B1(new_n917), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n916), .A2(new_n924), .A3(new_n921), .A4(new_n918), .ZN(new_n925));
  AOI21_X1  g739(.A(G953), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n910), .B1(new_n926), .B2(new_n903), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n928), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n930), .B(new_n910), .C1(new_n926), .C2(new_n903), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(G72));
  INV_X1    g746(.A(new_n646), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n923), .A2(new_n769), .A3(new_n925), .ZN(new_n934));
  XNOR2_X1  g748(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n935));
  NAND2_X1  g749(.A1(G472), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n935), .B(new_n936), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT127), .Z(new_n938));
  AOI21_X1  g752(.A(new_n933), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n933), .A2(new_n937), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n795), .A2(new_n802), .ZN(new_n941));
  AOI211_X1 g755(.A(new_n940), .B(new_n941), .C1(new_n537), .C2(new_n557), .ZN(new_n942));
  INV_X1    g756(.A(new_n769), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n938), .B1(new_n909), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n944), .A2(new_n537), .A3(new_n557), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n847), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n939), .A2(new_n942), .A3(new_n946), .ZN(G57));
endmodule


