//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n187));
  XNOR2_X1  g001(.A(G125), .B(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT16), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G125), .ZN(new_n192));
  AND3_X1   g006(.A1(new_n189), .A2(G146), .A3(new_n192), .ZN(new_n193));
  AOI21_X1  g007(.A(G146), .B1(new_n189), .B2(new_n192), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(G128), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(new_n199), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G110), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT74), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n204), .B1(new_n197), .B2(G128), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(KEYINPUT74), .A3(G119), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(new_n199), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT24), .B(G110), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n203), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n195), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n189), .A2(G146), .A3(new_n192), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT64), .B(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n188), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n207), .A2(new_n208), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n202), .A2(G110), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n211), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n187), .B1(new_n210), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT22), .B(G137), .ZN(new_n219));
  INV_X1    g033(.A(G221), .ZN(new_n220));
  INV_X1    g034(.A(G234), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n220), .A2(new_n221), .A3(G953), .ZN(new_n222));
  XOR2_X1   g036(.A(new_n219), .B(new_n222), .Z(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  OAI221_X1 g038(.A(new_n203), .B1(new_n207), .B2(new_n208), .C1(new_n193), .C2(new_n194), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(KEYINPUT75), .A3(new_n216), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n218), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  XOR2_X1   g041(.A(KEYINPUT71), .B(G902), .Z(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n225), .A2(new_n216), .A3(new_n223), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT76), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(KEYINPUT25), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(G217), .B1(new_n228), .B2(new_n221), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n236), .B(KEYINPUT73), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n227), .A2(new_n229), .A3(new_n230), .A4(new_n233), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n227), .A2(new_n230), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n237), .A2(G902), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(KEYINPUT77), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n239), .A2(KEYINPUT78), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT78), .B1(new_n239), .B2(new_n244), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G146), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT64), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G146), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n252), .A3(G143), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n249), .A2(G143), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n200), .B1(new_n253), .B2(KEYINPUT1), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n249), .A2(G143), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n250), .A2(new_n252), .ZN(new_n261));
  INV_X1    g075(.A(G143), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n257), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT11), .ZN(new_n265));
  INV_X1    g079(.A(G134), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(G137), .ZN(new_n267));
  INV_X1    g081(.A(G137), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(KEYINPUT11), .A3(G134), .ZN(new_n269));
  INV_X1    g083(.A(G131), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n266), .A2(G137), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n267), .A2(new_n269), .A3(new_n270), .A4(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n268), .A2(G134), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n266), .A2(G137), .ZN(new_n274));
  OAI21_X1  g088(.A(G131), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT66), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n272), .A2(new_n275), .A3(KEYINPUT66), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n264), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT67), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT30), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n267), .A2(new_n271), .A3(new_n269), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G131), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n272), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n259), .B1(new_n212), .B2(G143), .ZN(new_n284));
  AND2_X1   g098(.A1(KEYINPUT0), .A2(G128), .ZN(new_n285));
  NOR2_X1   g099(.A1(KEYINPUT0), .A2(G128), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n254), .B1(new_n212), .B2(G143), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT65), .B1(new_n289), .B2(new_n285), .ZN(new_n290));
  AND4_X1   g104(.A1(KEYINPUT65), .A2(new_n253), .A3(new_n255), .A4(new_n285), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n283), .B(new_n288), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT67), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n264), .B(new_n293), .C1(new_n276), .C2(new_n277), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n279), .A2(new_n280), .A3(new_n292), .A4(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n264), .A2(new_n275), .A3(new_n272), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT30), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(G116), .B(G119), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(KEYINPUT68), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT2), .B(G113), .Z(new_n302));
  XOR2_X1   g116(.A(new_n301), .B(new_n302), .Z(new_n303));
  NAND2_X1  g117(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(G237), .A2(G953), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G210), .ZN(new_n306));
  XOR2_X1   g120(.A(new_n306), .B(KEYINPUT27), .Z(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT26), .B(G101), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n303), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(new_n296), .A3(new_n292), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n304), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT31), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n297), .A2(new_n303), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n316), .B1(new_n299), .B2(new_n303), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(KEYINPUT31), .A3(new_n310), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT69), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n294), .A2(new_n292), .ZN(new_n320));
  INV_X1    g134(.A(new_n276), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n272), .A2(new_n275), .A3(KEYINPUT66), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n293), .B1(new_n323), .B2(new_n264), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n319), .B(new_n303), .C1(new_n320), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n312), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n279), .A2(new_n292), .A3(new_n294), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n319), .B1(new_n327), .B2(new_n303), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT28), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n297), .A2(KEYINPUT70), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT70), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n292), .A2(new_n296), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n303), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  OR2_X1    g147(.A1(new_n333), .A2(KEYINPUT28), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n315), .A2(new_n318), .B1(new_n335), .B2(new_n309), .ZN(new_n336));
  NOR2_X1   g150(.A1(G472), .A2(G902), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT32), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n333), .A2(KEYINPUT28), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n303), .B1(new_n320), .B2(new_n324), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT69), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(new_n325), .A3(new_n312), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n340), .B1(new_n343), .B2(KEYINPUT28), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT31), .B1(new_n317), .B2(new_n310), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n311), .B1(new_n295), .B2(new_n298), .ZN(new_n346));
  NOR4_X1   g160(.A1(new_n346), .A2(new_n314), .A3(new_n309), .A4(new_n316), .ZN(new_n347));
  OAI22_X1  g161(.A1(new_n344), .A2(new_n310), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT32), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n349), .A3(new_n337), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n339), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT72), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n311), .B1(new_n292), .B2(new_n296), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT28), .B1(new_n316), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n309), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n354), .B(new_n356), .C1(new_n333), .C2(KEYINPUT28), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n352), .B1(new_n358), .B2(new_n228), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(KEYINPUT72), .A3(new_n229), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n355), .B1(new_n317), .B2(new_n310), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(new_n344), .B2(new_n310), .ZN(new_n363));
  OAI21_X1  g177(.A(G472), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n248), .B1(new_n351), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G214), .B1(G237), .B2(G902), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n368));
  INV_X1    g182(.A(G107), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(G104), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(G104), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G104), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(KEYINPUT3), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n369), .A2(KEYINPUT80), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT80), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G107), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G101), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n372), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT81), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n372), .A2(new_n378), .A3(new_n382), .A4(new_n379), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n372), .A2(new_n378), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n385), .B1(new_n386), .B2(G101), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT80), .B(G107), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n389), .A2(new_n374), .B1(new_n370), .B2(new_n371), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n390), .A2(KEYINPUT4), .A3(new_n379), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n388), .A2(new_n303), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n375), .A2(new_n377), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n373), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT82), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n371), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n369), .A2(KEYINPUT82), .A3(G104), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G101), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n300), .A2(KEYINPUT5), .ZN(new_n402));
  INV_X1    g216(.A(G116), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n403), .A2(KEYINPUT5), .A3(G119), .ZN(new_n404));
  INV_X1    g218(.A(G113), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n402), .A2(new_n406), .B1(new_n302), .B2(new_n300), .ZN(new_n407));
  AND4_X1   g221(.A1(KEYINPUT87), .A2(new_n384), .A3(new_n401), .A4(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n379), .B1(new_n395), .B2(new_n399), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(new_n381), .B2(new_n383), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT87), .B1(new_n410), .B2(new_n407), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n393), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G110), .B(G122), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n393), .B(new_n413), .C1(new_n408), .C2(new_n411), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(KEYINPUT6), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n288), .B1(new_n290), .B2(new_n291), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G125), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT88), .B1(new_n264), .B2(G125), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G224), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(G953), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  OR3_X1    g238(.A1(new_n264), .A2(KEYINPUT88), .A3(G125), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n421), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n419), .A3(new_n420), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n423), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n412), .A2(new_n430), .A3(new_n414), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n417), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT89), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n417), .A2(KEYINPUT89), .A3(new_n429), .A4(new_n431), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n421), .A2(KEYINPUT7), .A3(new_n424), .A4(new_n425), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT7), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n427), .B1(new_n438), .B2(new_n423), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n413), .B(KEYINPUT8), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n410), .A2(new_n407), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n410), .A2(new_n407), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n437), .A2(new_n416), .A3(new_n439), .A4(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G902), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n436), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G210), .B1(G237), .B2(G902), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n436), .A2(new_n449), .A3(new_n447), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n367), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(G143), .B1(new_n305), .B2(G214), .ZN(new_n454));
  INV_X1    g268(.A(G237), .ZN(new_n455));
  INV_X1    g269(.A(G953), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n455), .A2(new_n456), .A3(G143), .A4(G214), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT90), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT90), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n305), .A2(new_n459), .A3(G143), .A4(G214), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n454), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT91), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT18), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n461), .A2(new_n270), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT93), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(KEYINPUT18), .A3(G131), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT92), .ZN(new_n469));
  INV_X1    g283(.A(G125), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(G140), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n191), .A2(G125), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n469), .B(G146), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT92), .B1(new_n212), .B2(new_n188), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n188), .A2(new_n249), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n465), .A2(new_n466), .A3(new_n468), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n468), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT93), .B1(new_n478), .B2(new_n464), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G113), .B(G122), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(new_n373), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n461), .A2(new_n270), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT17), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n461), .B(new_n270), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n195), .B(new_n484), .C1(new_n485), .C2(KEYINPUT17), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n480), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n482), .B1(new_n480), .B2(new_n486), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n445), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G475), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n188), .B(KEYINPUT19), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n193), .B1(new_n212), .B2(new_n492), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n477), .A2(new_n479), .B1(new_n485), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n487), .B1(new_n482), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT20), .ZN(new_n496));
  NOR2_X1   g310(.A1(G475), .A2(G902), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n496), .B1(new_n495), .B2(new_n497), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n491), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n200), .A2(G143), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n262), .A2(G128), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n501), .A2(new_n502), .A3(G134), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n403), .A2(G122), .ZN(new_n504));
  INV_X1    g318(.A(G122), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n505), .A2(G116), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n394), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G116), .B(G122), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n389), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n503), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n200), .A2(G143), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n501), .B1(KEYINPUT13), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n501), .A2(KEYINPUT13), .ZN(new_n513));
  OAI21_X1  g327(.A(G134), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT94), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT94), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n510), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n509), .B(KEYINPUT95), .ZN(new_n520));
  INV_X1    g334(.A(new_n501), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n266), .B1(new_n521), .B2(new_n511), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n504), .A2(KEYINPUT14), .ZN(new_n523));
  MUX2_X1   g337(.A(new_n523), .B(KEYINPUT14), .S(new_n506), .Z(new_n524));
  OAI221_X1 g338(.A(new_n520), .B1(new_n503), .B2(new_n522), .C1(new_n369), .C2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT9), .B(G234), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(KEYINPUT79), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(G217), .A3(new_n456), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n519), .A2(new_n525), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n530), .B1(new_n519), .B2(new_n525), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n229), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G478), .ZN(new_n535));
  NOR2_X1   g349(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n534), .B(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n456), .A2(G952), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(G234), .B2(G237), .ZN(new_n542));
  AOI211_X1 g356(.A(new_n456), .B(new_n229), .C1(G234), .C2(G237), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT21), .B(G898), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n500), .A2(new_n540), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n220), .B1(new_n528), .B2(new_n445), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(G110), .B(G140), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n456), .A2(G227), .ZN(new_n550));
  XOR2_X1   g364(.A(new_n549), .B(new_n550), .Z(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n418), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n391), .B1(new_n384), .B2(new_n387), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n253), .A2(new_n255), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT1), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(G143), .B2(new_n249), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT83), .ZN(new_n558));
  OAI21_X1  g372(.A(G128), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n259), .A2(new_n558), .A3(KEYINPUT1), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n555), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n257), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n384), .A2(new_n563), .A3(new_n401), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT10), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n553), .A2(new_n554), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT84), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n382), .B1(new_n390), .B2(new_n379), .ZN(new_n568));
  INV_X1    g382(.A(new_n383), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n401), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n264), .A2(KEYINPUT10), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n410), .A2(KEYINPUT84), .A3(KEYINPUT10), .A4(new_n264), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n283), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n566), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n575), .B1(new_n566), .B2(new_n574), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n552), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT86), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n576), .A2(new_n580), .A3(new_n551), .ZN(new_n581));
  INV_X1    g395(.A(new_n264), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n570), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n575), .B1(new_n583), .B2(new_n564), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT12), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n580), .B1(new_n576), .B2(new_n551), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n579), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(G469), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n588), .A2(new_n589), .A3(new_n229), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n583), .A2(new_n564), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n591), .A2(KEYINPUT12), .A3(new_n283), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT12), .B1(new_n591), .B2(new_n283), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n576), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n552), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT85), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n576), .A2(new_n596), .A3(new_n551), .ZN(new_n597));
  INV_X1    g411(.A(new_n578), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n596), .B1(new_n576), .B2(new_n551), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n595), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n589), .B1(new_n601), .B2(new_n445), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n546), .B(new_n548), .C1(new_n590), .C2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n365), .A2(new_n453), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G101), .ZN(G3));
  NOR2_X1   g420(.A1(new_n228), .A2(new_n535), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT33), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n519), .A2(new_n525), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n529), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n609), .B1(new_n611), .B2(new_n531), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n607), .B1(new_n608), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n228), .B1(new_n611), .B2(new_n531), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT98), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT97), .B(G478), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n616), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT98), .B1(new_n534), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n613), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n500), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n545), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n453), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n247), .B(new_n548), .C1(new_n590), .C2(new_n602), .ZN(new_n625));
  OAI21_X1  g439(.A(G472), .B1(new_n336), .B2(new_n228), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n348), .A2(new_n337), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT99), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT34), .B(G104), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  XOR2_X1   g447(.A(new_n545), .B(KEYINPUT100), .Z(new_n634));
  AOI21_X1  g448(.A(new_n449), .B1(new_n436), .B2(new_n447), .ZN(new_n635));
  AOI211_X1 g449(.A(new_n450), .B(new_n446), .C1(new_n434), .C2(new_n435), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n366), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n500), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n540), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n629), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT101), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  AND2_X1   g458(.A1(new_n218), .A2(new_n226), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n224), .A2(KEYINPUT36), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  OR2_X1    g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n645), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n648), .A2(new_n649), .A3(new_n243), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n239), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n628), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n604), .A3(new_n453), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT37), .B(G110), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  OAI21_X1  g470(.A(new_n548), .B1(new_n590), .B2(new_n602), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n351), .B2(new_n364), .ZN(new_n658));
  INV_X1    g472(.A(G900), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n542), .B1(new_n543), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT102), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n639), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n658), .A2(new_n453), .A3(new_n651), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  OAI21_X1  g478(.A(new_n309), .B1(new_n316), .B2(new_n353), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n313), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n666), .B2(G902), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n351), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT103), .Z(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n601), .A2(new_n445), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(G469), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n588), .A2(new_n589), .A3(new_n229), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n547), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n661), .B(KEYINPUT39), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT40), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n635), .A2(new_n636), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT38), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n500), .A2(new_n540), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n366), .A3(new_n652), .ZN(new_n683));
  NOR4_X1   g497(.A1(new_n670), .A2(new_n678), .A3(new_n680), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n262), .ZN(G45));
  INV_X1    g499(.A(new_n661), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n500), .A2(new_n620), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n453), .A2(KEYINPUT104), .A3(new_n687), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n687), .B(new_n366), .C1(new_n635), .C2(new_n636), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n688), .A2(new_n651), .A3(new_n658), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  NAND2_X1  g507(.A1(new_n588), .A2(new_n229), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G469), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n548), .A3(new_n673), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT105), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n348), .A2(new_n349), .A3(new_n337), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n349), .B1(new_n348), .B2(new_n337), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n364), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n695), .A2(new_n701), .A3(new_n548), .A4(new_n673), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n697), .A2(new_n700), .A3(new_n247), .A4(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n623), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT106), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n704), .B(new_n706), .ZN(G15));
  INV_X1    g521(.A(new_n639), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n453), .A2(new_n708), .A3(new_n634), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n703), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n403), .ZN(G18));
  NAND2_X1  g525(.A1(new_n697), .A2(new_n702), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n546), .A2(new_n651), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n700), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n713), .A2(new_n716), .A3(new_n453), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  INV_X1    g532(.A(G472), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n348), .B2(new_n229), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n239), .A2(new_n244), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n315), .A2(new_n318), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n334), .A2(new_n354), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n309), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n338), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n720), .A2(new_n721), .A3(new_n725), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n697), .A2(new_n702), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n637), .A2(new_n681), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  INV_X1    g544(.A(new_n725), .ZN(new_n731));
  AND4_X1   g545(.A1(new_n626), .A2(new_n687), .A3(new_n731), .A4(new_n651), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n453), .A3(new_n697), .A4(new_n702), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  NAND4_X1  g548(.A1(new_n679), .A2(new_n674), .A3(new_n366), .A4(new_n687), .ZN(new_n735));
  INV_X1    g549(.A(new_n721), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n700), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT42), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n635), .A2(new_n636), .A3(new_n367), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n621), .A2(KEYINPUT42), .A3(new_n661), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n365), .A2(new_n674), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  NAND4_X1  g557(.A1(new_n739), .A2(new_n700), .A3(new_n247), .A4(new_n674), .ZN(new_n744));
  INV_X1    g558(.A(new_n662), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT107), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n679), .A2(new_n674), .A3(new_n366), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n365), .A4(new_n662), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  NAND2_X1  g566(.A1(new_n638), .A2(new_n620), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT109), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n753), .A2(KEYINPUT109), .A3(KEYINPUT43), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n628), .A3(new_n651), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n739), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n601), .B(KEYINPUT45), .ZN(new_n764));
  OAI21_X1  g578(.A(G469), .B1(new_n764), .B2(G902), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n766), .A3(KEYINPUT46), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n767), .B(new_n673), .C1(KEYINPUT46), .C2(new_n765), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n766), .B1(new_n765), .B2(KEYINPUT46), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n548), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n770), .A2(new_n675), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n763), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(new_n268), .ZN(G39));
  NAND2_X1  g587(.A1(new_n679), .A2(new_n366), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n248), .A2(new_n687), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n774), .A2(new_n700), .A3(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT47), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n770), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  OAI211_X1 g593(.A(KEYINPUT47), .B(new_n548), .C1(new_n768), .C2(new_n769), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n776), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  OR2_X1    g597(.A1(G952), .A2(G953), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n758), .A2(new_n542), .A3(new_n726), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n774), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n778), .A2(KEYINPUT114), .A3(new_n780), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n695), .A2(new_n673), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n547), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT114), .B1(new_n778), .B2(new_n780), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n786), .B(new_n788), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n720), .A2(new_n652), .A3(new_n725), .ZN(new_n795));
  INV_X1    g609(.A(new_n542), .ZN(new_n796));
  OR3_X1    g610(.A1(new_n712), .A2(KEYINPUT116), .A3(new_n774), .ZN(new_n797));
  OAI21_X1  g611(.A(KEYINPUT116), .B1(new_n712), .B2(new_n774), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n800), .A3(new_n758), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n800), .B1(new_n799), .B2(new_n758), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n795), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n799), .A2(new_n247), .A3(new_n670), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n500), .A2(new_n620), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n680), .A2(new_n367), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n713), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n807), .B1(new_n809), .B2(new_n787), .ZN(new_n810));
  INV_X1    g624(.A(new_n787), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(new_n808), .A3(KEYINPUT50), .A4(new_n713), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n805), .A2(new_n806), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n794), .A2(new_n804), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n793), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n791), .A3(new_n789), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n786), .B1(new_n816), .B2(new_n788), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n785), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n778), .A2(new_n780), .A3(new_n791), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n785), .B1(new_n819), .B2(new_n788), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n804), .A2(new_n813), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n453), .A2(new_n697), .A3(new_n702), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n787), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n621), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n541), .B(new_n823), .C1(new_n805), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n799), .A2(new_n758), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT117), .ZN(new_n827));
  AOI211_X1 g641(.A(KEYINPUT48), .B(new_n737), .C1(new_n827), .C2(new_n801), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT48), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n827), .A2(new_n801), .ZN(new_n830));
  INV_X1    g644(.A(new_n737), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n821), .B(new_n825), .C1(new_n828), .C2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n818), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n651), .A2(KEYINPUT112), .A3(new_n661), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT112), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n652), .B2(new_n686), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n657), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(new_n453), .A3(new_n668), .A4(new_n682), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n692), .A2(new_n663), .A3(new_n733), .A4(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT52), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n540), .B(KEYINPUT110), .ZN(new_n844));
  NOR4_X1   g658(.A1(new_n844), .A2(new_n652), .A3(new_n500), .A4(new_n661), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n658), .A2(new_n739), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n738), .A2(new_n741), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT111), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n626), .A2(new_n687), .A3(new_n731), .A4(new_n651), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n747), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n732), .A2(KEYINPUT111), .A3(new_n674), .A4(new_n739), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n697), .A2(new_n702), .A3(new_n726), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n451), .A2(new_n452), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(new_n366), .A3(new_n634), .A4(new_n682), .ZN(new_n856));
  OAI22_X1  g670(.A1(new_n822), .A2(new_n715), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n857), .A2(new_n710), .A3(new_n704), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n844), .A2(new_n638), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n621), .ZN(new_n860));
  INV_X1    g674(.A(new_n637), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n629), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n862), .A2(new_n605), .A3(new_n654), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n853), .A2(new_n858), .A3(new_n751), .A4(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n836), .B1(new_n843), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n850), .A2(new_n851), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n742), .A2(new_n751), .A3(new_n867), .A4(new_n846), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n663), .A2(new_n733), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(KEYINPUT52), .A3(new_n692), .A4(new_n841), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT52), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n842), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n862), .A2(new_n605), .A3(new_n654), .A4(KEYINPUT53), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n624), .A2(new_n713), .A3(new_n365), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n713), .A2(new_n640), .A3(new_n365), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n876), .A2(new_n877), .A3(new_n717), .A4(new_n729), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT113), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n875), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n858), .A2(KEYINPUT113), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n869), .A2(new_n874), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n865), .A2(new_n866), .A3(new_n882), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n843), .A2(new_n864), .A3(new_n836), .ZN(new_n884));
  INV_X1    g698(.A(new_n857), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n863), .A2(new_n885), .A3(new_n876), .A4(new_n877), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n868), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT53), .B1(new_n887), .B2(new_n874), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n883), .B1(new_n889), .B2(new_n866), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n784), .B1(new_n835), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n790), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n892), .A2(KEYINPUT49), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(KEYINPUT49), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n736), .A2(new_n366), .A3(new_n548), .ZN(new_n895));
  NOR4_X1   g709(.A1(new_n893), .A2(new_n894), .A3(new_n753), .A4(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n670), .A2(new_n896), .A3(new_n680), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n891), .A2(new_n897), .ZN(G75));
  NAND2_X1  g712(.A1(new_n865), .A2(new_n882), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(new_n228), .A3(new_n450), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT56), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n417), .A2(new_n431), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n429), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(KEYINPUT55), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(KEYINPUT118), .B2(new_n901), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n903), .A2(KEYINPUT55), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n900), .A2(new_n901), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n907), .B1(new_n900), .B2(new_n901), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n456), .A2(G952), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(G51));
  NAND2_X1  g725(.A1(new_n764), .A2(G469), .ZN(new_n912));
  AOI211_X1 g726(.A(new_n229), .B(new_n912), .C1(new_n865), .C2(new_n882), .ZN(new_n913));
  NAND2_X1  g727(.A1(G469), .A2(G902), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT57), .Z(new_n915));
  AND3_X1   g729(.A1(new_n865), .A2(new_n866), .A3(new_n882), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n866), .B1(new_n865), .B2(new_n882), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n913), .B1(new_n918), .B2(new_n588), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT119), .B1(new_n919), .B2(new_n910), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT119), .ZN(new_n921));
  INV_X1    g735(.A(new_n910), .ZN(new_n922));
  INV_X1    g736(.A(new_n588), .ZN(new_n923));
  AND4_X1   g737(.A1(new_n874), .A2(new_n869), .A3(new_n880), .A4(new_n881), .ZN(new_n924));
  OAI21_X1  g738(.A(KEYINPUT54), .B1(new_n924), .B2(new_n888), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n883), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n923), .B1(new_n926), .B2(new_n915), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n921), .B(new_n922), .C1(new_n927), .C2(new_n913), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n920), .A2(new_n928), .ZN(G54));
  NAND4_X1  g743(.A1(new_n899), .A2(KEYINPUT58), .A3(G475), .A4(new_n228), .ZN(new_n930));
  INV_X1    g744(.A(new_n495), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n930), .A2(KEYINPUT120), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n922), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT120), .B1(new_n930), .B2(new_n931), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(G60));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT59), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n608), .A2(new_n612), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT121), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n926), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n939), .B1(new_n890), .B2(new_n937), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n940), .A2(new_n941), .A3(new_n910), .ZN(G63));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT60), .Z(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n865), .B2(new_n882), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n922), .B1(new_n946), .B2(new_n241), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n648), .A2(new_n649), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n948), .A2(new_n950), .A3(KEYINPUT122), .A4(new_n951), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n951), .A2(KEYINPUT122), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(KEYINPUT122), .ZN(new_n954));
  INV_X1    g768(.A(new_n950), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n953), .B(new_n954), .C1(new_n955), .C2(new_n947), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n952), .A2(new_n956), .ZN(G66));
  NOR3_X1   g771(.A1(new_n544), .A2(new_n422), .A3(new_n456), .ZN(new_n958));
  INV_X1    g772(.A(new_n886), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(new_n456), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n902), .B1(G898), .B2(new_n456), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(G69));
  XNOR2_X1  g776(.A(new_n492), .B(KEYINPUT123), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n299), .B(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(G900), .B2(G953), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n870), .A2(new_n692), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n772), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n771), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n968), .A2(new_n453), .A3(new_n682), .A4(new_n831), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n742), .A2(new_n751), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n967), .A2(new_n969), .A3(new_n782), .A4(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n965), .B1(new_n971), .B2(G953), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n684), .A2(new_n966), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT62), .ZN(new_n974));
  INV_X1    g788(.A(new_n772), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n860), .B(KEYINPUT125), .ZN(new_n976));
  INV_X1    g790(.A(new_n677), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n976), .A2(new_n365), .A3(new_n977), .A4(new_n739), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n975), .A2(new_n782), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(G953), .B1(new_n974), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n964), .B(KEYINPUT124), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n972), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n456), .B1(G227), .B2(G900), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n983), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n972), .B(new_n985), .C1(new_n980), .C2(new_n981), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n984), .A2(new_n986), .ZN(G72));
  NAND2_X1  g801(.A1(new_n317), .A2(new_n309), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n310), .B1(new_n346), .B2(new_n316), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g804(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n991));
  NOR2_X1   g805(.A1(new_n719), .A2(new_n445), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT127), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n922), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n889), .A2(new_n993), .A3(new_n990), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n974), .A2(new_n979), .ZN(new_n998));
  OAI22_X1  g812(.A1(new_n998), .A2(new_n989), .B1(new_n971), .B2(new_n988), .ZN(new_n999));
  AOI211_X1 g813(.A(new_n996), .B(new_n997), .C1(new_n999), .C2(new_n959), .ZN(G57));
endmodule


