

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735;

  NOR2_X1 U367 ( .A1(G953), .A2(G237), .ZN(n439) );
  XNOR2_X1 U368 ( .A(G902), .B(KEYINPUT15), .ZN(n641) );
  NAND2_X2 U369 ( .A1(n547), .A2(n533), .ZN(n612) );
  NOR2_X2 U370 ( .A1(n582), .A2(n573), .ZN(n567) );
  AND2_X1 U371 ( .A1(n364), .A2(n351), .ZN(n363) );
  NOR2_X1 U372 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U373 ( .A(n506), .B(KEYINPUT40), .ZN(n401) );
  XNOR2_X1 U374 ( .A(n513), .B(KEYINPUT19), .ZN(n556) );
  OR2_X1 U375 ( .A1(n562), .A2(n614), .ZN(n454) );
  XNOR2_X1 U376 ( .A(n531), .B(n530), .ZN(n596) );
  XNOR2_X1 U377 ( .A(n435), .B(n434), .ZN(n531) );
  XNOR2_X1 U378 ( .A(n356), .B(G110), .ZN(n466) );
  XOR2_X1 U379 ( .A(G146), .B(G125), .Z(n469) );
  XNOR2_X2 U380 ( .A(n716), .B(G146), .ZN(n448) );
  INV_X1 U381 ( .A(KEYINPUT87), .ZN(n366) );
  NOR2_X1 U382 ( .A1(n615), .A2(n614), .ZN(n613) );
  INV_X1 U383 ( .A(G469), .ZN(n434) );
  NOR2_X1 U384 ( .A1(G902), .A2(n682), .ZN(n435) );
  INV_X1 U385 ( .A(KEYINPUT72), .ZN(n356) );
  AND2_X1 U386 ( .A1(n616), .A2(n395), .ZN(n381) );
  XNOR2_X1 U387 ( .A(n382), .B(n541), .ZN(n369) );
  NAND2_X1 U388 ( .A1(n367), .A2(n366), .ZN(n365) );
  INV_X1 U389 ( .A(n731), .ZN(n367) );
  XNOR2_X1 U390 ( .A(n379), .B(n378), .ZN(n377) );
  INV_X1 U391 ( .A(KEYINPUT44), .ZN(n378) );
  XNOR2_X1 U392 ( .A(n469), .B(n414), .ZN(n482) );
  XNOR2_X1 U393 ( .A(KEYINPUT10), .B(KEYINPUT66), .ZN(n414) );
  XNOR2_X1 U394 ( .A(G143), .B(G140), .ZN(n487) );
  INV_X1 U395 ( .A(KEYINPUT12), .ZN(n486) );
  XNOR2_X1 U396 ( .A(n482), .B(n354), .ZN(n485) );
  INV_X1 U397 ( .A(KEYINPUT11), .ZN(n354) );
  XNOR2_X1 U398 ( .A(n512), .B(n479), .ZN(n615) );
  AND2_X1 U399 ( .A1(n534), .A2(n394), .ZN(n392) );
  XNOR2_X1 U400 ( .A(n492), .B(n491), .ZN(n524) );
  OR2_X1 U401 ( .A1(n698), .A2(G902), .ZN(n396) );
  XNOR2_X1 U402 ( .A(G101), .B(KEYINPUT3), .ZN(n440) );
  XOR2_X1 U403 ( .A(G116), .B(G107), .Z(n497) );
  XNOR2_X1 U404 ( .A(n464), .B(G122), .ZN(n483) );
  XNOR2_X1 U405 ( .A(G113), .B(G104), .ZN(n464) );
  INV_X1 U406 ( .A(KEYINPUT16), .ZN(n355) );
  INV_X1 U407 ( .A(n596), .ZN(n561) );
  INV_X1 U408 ( .A(KEYINPUT34), .ZN(n359) );
  XNOR2_X1 U409 ( .A(n557), .B(KEYINPUT0), .ZN(n583) );
  NOR2_X1 U410 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U411 ( .A(n463), .B(n399), .ZN(n398) );
  INV_X1 U412 ( .A(KEYINPUT74), .ZN(n399) );
  XNOR2_X1 U413 ( .A(n583), .B(KEYINPUT94), .ZN(n580) );
  INV_X1 U414 ( .A(n550), .ZN(n601) );
  XNOR2_X1 U415 ( .A(n430), .B(n429), .ZN(n433) );
  AND2_X1 U416 ( .A1(n647), .A2(G953), .ZN(n701) );
  XNOR2_X1 U417 ( .A(n520), .B(n518), .ZN(n521) );
  XNOR2_X1 U418 ( .A(n384), .B(n511), .ZN(n383) );
  NAND2_X1 U419 ( .A1(n400), .A2(n401), .ZN(n384) );
  NAND2_X1 U420 ( .A1(G234), .A2(G237), .ZN(n455) );
  XNOR2_X1 U421 ( .A(G116), .B(G113), .ZN(n442) );
  XNOR2_X1 U422 ( .A(KEYINPUT5), .B(G137), .ZN(n443) );
  OR2_X1 U423 ( .A1(G237), .A2(G902), .ZN(n476) );
  NAND2_X1 U424 ( .A1(n362), .A2(n366), .ZN(n361) );
  INV_X1 U425 ( .A(n369), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n376), .B(n352), .ZN(n710) );
  INV_X1 U427 ( .A(KEYINPUT96), .ZN(n406) );
  XNOR2_X1 U428 ( .A(KEYINPUT8), .B(KEYINPUT65), .ZN(n410) );
  XNOR2_X1 U429 ( .A(n489), .B(n353), .ZN(n686) );
  XNOR2_X1 U430 ( .A(n490), .B(n488), .ZN(n353) );
  XNOR2_X1 U431 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U432 ( .A(n466), .B(n402), .ZN(n424) );
  XNOR2_X1 U433 ( .A(n375), .B(n374), .ZN(n626) );
  INV_X1 U434 ( .A(KEYINPUT41), .ZN(n374) );
  NAND2_X1 U435 ( .A1(n398), .A2(n397), .ZN(n480) );
  NAND2_X1 U436 ( .A1(n388), .A2(n387), .ZN(n389) );
  NOR2_X1 U437 ( .A1(n392), .A2(n391), .ZN(n390) );
  NOR2_X1 U438 ( .A1(n512), .A2(n614), .ZN(n513) );
  XNOR2_X1 U439 ( .A(n437), .B(n436), .ZN(n578) );
  INV_X1 U440 ( .A(G953), .ZN(n725) );
  XNOR2_X1 U441 ( .A(n465), .B(n497), .ZN(n370) );
  XNOR2_X1 U442 ( .A(n467), .B(n483), .ZN(n371) );
  XNOR2_X1 U443 ( .A(n466), .B(n355), .ZN(n467) );
  XNOR2_X1 U444 ( .A(n373), .B(n372), .ZN(n735) );
  INV_X1 U445 ( .A(KEYINPUT42), .ZN(n372) );
  OR2_X1 U446 ( .A1(n626), .A2(n514), .ZN(n373) );
  AND2_X1 U447 ( .A1(n358), .A2(n357), .ZN(n570) );
  INV_X1 U448 ( .A(n569), .ZN(n357) );
  XNOR2_X1 U449 ( .A(n360), .B(n359), .ZN(n358) );
  OR2_X1 U450 ( .A1(n572), .A2(n563), .ZN(n666) );
  XNOR2_X1 U451 ( .A(n684), .B(n683), .ZN(n685) );
  INV_X1 U452 ( .A(n600), .ZN(n395) );
  AND2_X1 U453 ( .A1(n550), .A2(n395), .ZN(n565) );
  XOR2_X1 U454 ( .A(n380), .B(KEYINPUT22), .Z(n347) );
  XOR2_X1 U455 ( .A(n418), .B(n417), .Z(n348) );
  XNOR2_X1 U456 ( .A(n480), .B(KEYINPUT39), .ZN(n546) );
  OR2_X1 U457 ( .A1(n586), .A2(n585), .ZN(n349) );
  NOR2_X1 U458 ( .A1(n512), .A2(n569), .ZN(n350) );
  AND2_X1 U459 ( .A1(n365), .A2(n639), .ZN(n351) );
  BUF_X1 U460 ( .A(n562), .Z(n604) );
  INV_X1 U461 ( .A(n510), .ZN(n394) );
  XOR2_X1 U462 ( .A(KEYINPUT86), .B(KEYINPUT45), .Z(n352) );
  XNOR2_X1 U463 ( .A(n371), .B(n370), .ZN(n704) );
  XNOR2_X2 U464 ( .A(n640), .B(KEYINPUT2), .ZN(n642) );
  NAND2_X1 U465 ( .A1(n568), .A2(n580), .ZN(n360) );
  NAND2_X2 U466 ( .A1(n363), .A2(n361), .ZN(n723) );
  NAND2_X1 U467 ( .A1(n369), .A2(n368), .ZN(n364) );
  AND2_X1 U468 ( .A1(n731), .A2(KEYINPUT87), .ZN(n368) );
  NAND2_X1 U469 ( .A1(n613), .A2(n616), .ZN(n375) );
  OR2_X2 U470 ( .A1(n524), .A2(n515), .ZN(n547) );
  NAND2_X1 U471 ( .A1(n377), .A2(n587), .ZN(n376) );
  NAND2_X1 U472 ( .A1(n571), .A2(n729), .ZN(n379) );
  NAND2_X1 U473 ( .A1(n583), .A2(n381), .ZN(n380) );
  NAND2_X1 U474 ( .A1(n385), .A2(n383), .ZN(n382) );
  XNOR2_X1 U475 ( .A(n386), .B(KEYINPUT67), .ZN(n385) );
  NAND2_X1 U476 ( .A1(n540), .A2(n539), .ZN(n386) );
  AND2_X1 U477 ( .A1(n509), .A2(n510), .ZN(n387) );
  INV_X1 U478 ( .A(n534), .ZN(n388) );
  NAND2_X1 U479 ( .A1(n390), .A2(n389), .ZN(n514) );
  NAND2_X1 U480 ( .A1(n393), .A2(n531), .ZN(n391) );
  NAND2_X1 U481 ( .A1(n604), .A2(n394), .ZN(n393) );
  XNOR2_X2 U482 ( .A(n396), .B(n348), .ZN(n550) );
  INV_X1 U483 ( .A(n615), .ZN(n397) );
  AND2_X1 U484 ( .A1(n398), .A2(n350), .ZN(n637) );
  INV_X1 U485 ( .A(n735), .ZN(n400) );
  XNOR2_X1 U486 ( .A(n401), .B(G131), .ZN(G33) );
  NOR2_X1 U487 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U488 ( .A1(n657), .A2(n701), .ZN(n659) );
  NOR2_X1 U489 ( .A1(n648), .A2(n701), .ZN(n650) );
  NOR2_X1 U490 ( .A1(n691), .A2(n701), .ZN(n692) );
  XNOR2_X1 U491 ( .A(n415), .B(n719), .ZN(n698) );
  XNOR2_X1 U492 ( .A(n413), .B(n412), .ZN(n415) );
  XNOR2_X1 U493 ( .A(n409), .B(n408), .ZN(n413) );
  AND2_X1 U494 ( .A1(G227), .A2(n725), .ZN(n402) );
  XOR2_X1 U495 ( .A(KEYINPUT76), .B(KEYINPUT95), .Z(n403) );
  INV_X1 U496 ( .A(n679), .ZN(n539) );
  XNOR2_X1 U497 ( .A(n407), .B(n406), .ZN(n408) );
  BUF_X1 U498 ( .A(n640), .Z(n590) );
  INV_X1 U499 ( .A(n562), .ZN(n509) );
  BUF_X1 U500 ( .A(n716), .Z(n717) );
  XNOR2_X1 U501 ( .A(n425), .B(n424), .ZN(n430) );
  XNOR2_X1 U502 ( .A(n688), .B(n687), .ZN(n689) );
  INV_X1 U503 ( .A(KEYINPUT119), .ZN(n634) );
  XNOR2_X1 U504 ( .A(n636), .B(n635), .ZN(G75) );
  XOR2_X1 U505 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n405) );
  XNOR2_X1 U506 ( .A(G128), .B(KEYINPUT68), .ZN(n404) );
  XNOR2_X1 U507 ( .A(n405), .B(n404), .ZN(n409) );
  XNOR2_X1 U508 ( .A(G119), .B(G110), .ZN(n407) );
  NAND2_X1 U509 ( .A1(n725), .A2(G234), .ZN(n411) );
  XNOR2_X1 U510 ( .A(n411), .B(n410), .ZN(n499) );
  NAND2_X1 U511 ( .A1(n499), .A2(G221), .ZN(n412) );
  XOR2_X2 U512 ( .A(G137), .B(G140), .Z(n426) );
  XNOR2_X1 U513 ( .A(n482), .B(n426), .ZN(n719) );
  XOR2_X1 U514 ( .A(KEYINPUT97), .B(KEYINPUT25), .Z(n418) );
  NAND2_X1 U515 ( .A1(G234), .A2(n641), .ZN(n416) );
  XNOR2_X1 U516 ( .A(KEYINPUT20), .B(n416), .ZN(n419) );
  NAND2_X1 U517 ( .A1(n419), .A2(G217), .ZN(n417) );
  XOR2_X1 U518 ( .A(KEYINPUT99), .B(KEYINPUT21), .Z(n421) );
  NAND2_X1 U519 ( .A1(n419), .A2(G221), .ZN(n420) );
  XNOR2_X1 U520 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U521 ( .A(KEYINPUT98), .B(n422), .ZN(n600) );
  XNOR2_X1 U522 ( .A(G107), .B(KEYINPUT75), .ZN(n423) );
  XNOR2_X1 U523 ( .A(n403), .B(n423), .ZN(n425) );
  XOR2_X1 U524 ( .A(n426), .B(G104), .Z(n427) );
  XNOR2_X1 U525 ( .A(n427), .B(G101), .ZN(n428) );
  INV_X1 U526 ( .A(n428), .ZN(n429) );
  XNOR2_X2 U527 ( .A(G143), .B(G128), .ZN(n496) );
  XNOR2_X2 U528 ( .A(n496), .B(KEYINPUT4), .ZN(n468) );
  INV_X1 U529 ( .A(G134), .ZN(n431) );
  XNOR2_X1 U530 ( .A(n431), .B(G131), .ZN(n432) );
  XNOR2_X2 U531 ( .A(n468), .B(n432), .ZN(n716) );
  XNOR2_X1 U532 ( .A(n433), .B(n448), .ZN(n682) );
  NAND2_X1 U533 ( .A1(n565), .A2(n531), .ZN(n437) );
  INV_X1 U534 ( .A(KEYINPUT100), .ZN(n436) );
  INV_X1 U535 ( .A(KEYINPUT73), .ZN(n438) );
  XNOR2_X1 U536 ( .A(n439), .B(n438), .ZN(n481) );
  NAND2_X1 U537 ( .A1(n481), .A2(G210), .ZN(n441) );
  XNOR2_X1 U538 ( .A(n440), .B(G119), .ZN(n465) );
  XNOR2_X1 U539 ( .A(n441), .B(n465), .ZN(n446) );
  XNOR2_X1 U540 ( .A(n442), .B(KEYINPUT71), .ZN(n444) );
  XNOR2_X1 U541 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U542 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U543 ( .A(n448), .B(n447), .ZN(n644) );
  OR2_X2 U544 ( .A1(n644), .A2(G902), .ZN(n450) );
  INV_X1 U545 ( .A(G472), .ZN(n449) );
  XNOR2_X2 U546 ( .A(n450), .B(n449), .ZN(n562) );
  NAND2_X1 U547 ( .A1(n476), .A2(G214), .ZN(n452) );
  INV_X1 U548 ( .A(KEYINPUT92), .ZN(n451) );
  XNOR2_X1 U549 ( .A(n452), .B(n451), .ZN(n614) );
  INV_X1 U550 ( .A(KEYINPUT30), .ZN(n453) );
  XNOR2_X1 U551 ( .A(n454), .B(n453), .ZN(n461) );
  XNOR2_X1 U552 ( .A(n455), .B(KEYINPUT93), .ZN(n456) );
  XOR2_X1 U553 ( .A(KEYINPUT14), .B(n456), .Z(n457) );
  NAND2_X1 U554 ( .A1(G952), .A2(n457), .ZN(n625) );
  NOR2_X1 U555 ( .A1(G953), .A2(n625), .ZN(n554) );
  AND2_X1 U556 ( .A1(G953), .A2(n457), .ZN(n458) );
  NAND2_X1 U557 ( .A1(G902), .A2(n458), .ZN(n552) );
  NOR2_X1 U558 ( .A1(G900), .A2(n552), .ZN(n459) );
  OR2_X1 U559 ( .A1(n554), .A2(n459), .ZN(n460) );
  XNOR2_X1 U560 ( .A(n460), .B(KEYINPUT80), .ZN(n507) );
  AND2_X1 U561 ( .A1(n461), .A2(n507), .ZN(n462) );
  NAND2_X1 U562 ( .A1(n578), .A2(n462), .ZN(n463) );
  XNOR2_X1 U563 ( .A(n469), .B(n468), .ZN(n474) );
  XOR2_X1 U564 ( .A(KEYINPUT90), .B(KEYINPUT17), .Z(n472) );
  NAND2_X1 U565 ( .A1(G224), .A2(n725), .ZN(n470) );
  XNOR2_X1 U566 ( .A(n470), .B(KEYINPUT18), .ZN(n471) );
  XNOR2_X1 U567 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U568 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U569 ( .A(n704), .B(n475), .ZN(n654) );
  NAND2_X1 U570 ( .A1(n654), .A2(n641), .ZN(n478) );
  NAND2_X1 U571 ( .A1(G210), .A2(n476), .ZN(n477) );
  XNOR2_X2 U572 ( .A(n478), .B(n477), .ZN(n512) );
  INV_X1 U573 ( .A(KEYINPUT38), .ZN(n479) );
  NAND2_X1 U574 ( .A1(G214), .A2(n481), .ZN(n490) );
  XNOR2_X1 U575 ( .A(G131), .B(n483), .ZN(n484) );
  XNOR2_X1 U576 ( .A(n485), .B(n484), .ZN(n489) );
  NOR2_X1 U577 ( .A1(G902), .A2(n686), .ZN(n492) );
  XNOR2_X1 U578 ( .A(KEYINPUT13), .B(G475), .ZN(n491) );
  XOR2_X1 U579 ( .A(KEYINPUT9), .B(KEYINPUT102), .Z(n494) );
  XNOR2_X1 U580 ( .A(G134), .B(G122), .ZN(n493) );
  XNOR2_X1 U581 ( .A(n494), .B(n493), .ZN(n503) );
  XOR2_X1 U582 ( .A(KEYINPUT7), .B(KEYINPUT103), .Z(n495) );
  XOR2_X1 U583 ( .A(n496), .B(n495), .Z(n498) );
  XNOR2_X1 U584 ( .A(n498), .B(n497), .ZN(n501) );
  NAND2_X1 U585 ( .A1(n499), .A2(G217), .ZN(n500) );
  XOR2_X1 U586 ( .A(n501), .B(n500), .Z(n502) );
  XNOR2_X1 U587 ( .A(n503), .B(n502), .ZN(n695) );
  NOR2_X1 U588 ( .A1(G902), .A2(n695), .ZN(n504) );
  INV_X1 U589 ( .A(n504), .ZN(n505) );
  XNOR2_X2 U590 ( .A(G478), .B(n505), .ZN(n523) );
  INV_X1 U591 ( .A(n523), .ZN(n515) );
  NAND2_X1 U592 ( .A1(n524), .A2(n515), .ZN(n533) );
  INV_X1 U593 ( .A(n533), .ZN(n673) );
  NAND2_X1 U594 ( .A1(n546), .A2(n673), .ZN(n506) );
  NOR2_X1 U595 ( .A1(n524), .A2(n523), .ZN(n616) );
  NOR2_X1 U596 ( .A1(n550), .A2(n600), .ZN(n508) );
  NAND2_X1 U597 ( .A1(n508), .A2(n507), .ZN(n534) );
  XOR2_X1 U598 ( .A(KEYINPUT106), .B(KEYINPUT28), .Z(n510) );
  XNOR2_X1 U599 ( .A(KEYINPUT89), .B(KEYINPUT46), .ZN(n511) );
  INV_X1 U600 ( .A(KEYINPUT84), .ZN(n518) );
  NOR2_X2 U601 ( .A1(n514), .A2(n556), .ZN(n670) );
  INV_X1 U602 ( .A(n670), .ZN(n516) );
  XNOR2_X1 U603 ( .A(n612), .B(KEYINPUT85), .ZN(n586) );
  NOR2_X1 U604 ( .A1(n516), .A2(n586), .ZN(n517) );
  NOR2_X1 U605 ( .A1(n518), .A2(n517), .ZN(n519) );
  NOR2_X1 U606 ( .A1(KEYINPUT47), .A2(n519), .ZN(n528) );
  INV_X1 U607 ( .A(n612), .ZN(n520) );
  NAND2_X1 U608 ( .A1(n521), .A2(n670), .ZN(n522) );
  NAND2_X1 U609 ( .A1(n522), .A2(KEYINPUT47), .ZN(n526) );
  NAND2_X1 U610 ( .A1(n524), .A2(n523), .ZN(n569) );
  INV_X1 U611 ( .A(n637), .ZN(n525) );
  NAND2_X1 U612 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U613 ( .A(n529), .B(KEYINPUT70), .ZN(n540) );
  XNOR2_X1 U614 ( .A(KEYINPUT1), .B(KEYINPUT64), .ZN(n530) );
  INV_X1 U615 ( .A(KEYINPUT6), .ZN(n532) );
  XNOR2_X1 U616 ( .A(n562), .B(n532), .ZN(n573) );
  NOR2_X1 U617 ( .A1(n533), .A2(n573), .ZN(n536) );
  NOR2_X1 U618 ( .A1(n614), .A2(n534), .ZN(n535) );
  NAND2_X1 U619 ( .A1(n536), .A2(n535), .ZN(n542) );
  NOR2_X1 U620 ( .A1(n512), .A2(n542), .ZN(n537) );
  XOR2_X1 U621 ( .A(KEYINPUT36), .B(n537), .Z(n538) );
  NOR2_X1 U622 ( .A1(n561), .A2(n538), .ZN(n679) );
  INV_X1 U623 ( .A(KEYINPUT48), .ZN(n541) );
  OR2_X1 U624 ( .A1(n542), .A2(n596), .ZN(n543) );
  XNOR2_X1 U625 ( .A(n543), .B(KEYINPUT43), .ZN(n544) );
  AND2_X1 U626 ( .A1(n544), .A2(n512), .ZN(n545) );
  XNOR2_X1 U627 ( .A(n545), .B(KEYINPUT105), .ZN(n731) );
  INV_X1 U628 ( .A(n547), .ZN(n676) );
  NAND2_X1 U629 ( .A1(n546), .A2(n676), .ZN(n639) );
  XNOR2_X1 U630 ( .A(KEYINPUT32), .B(KEYINPUT77), .ZN(n560) );
  XOR2_X1 U631 ( .A(KEYINPUT79), .B(n573), .Z(n548) );
  NAND2_X1 U632 ( .A1(n548), .A2(n596), .ZN(n549) );
  NOR2_X1 U633 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U634 ( .A(n551), .B(KEYINPUT78), .ZN(n558) );
  NOR2_X1 U635 ( .A1(G898), .A2(n552), .ZN(n553) );
  NOR2_X1 U636 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U637 ( .A1(n558), .A2(n347), .ZN(n559) );
  XNOR2_X1 U638 ( .A(n560), .B(n559), .ZN(n733) );
  NAND2_X1 U639 ( .A1(n561), .A2(n347), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n601), .A2(n604), .ZN(n563) );
  INV_X1 U641 ( .A(n666), .ZN(n564) );
  NOR2_X1 U642 ( .A1(n733), .A2(n564), .ZN(n571) );
  NAND2_X1 U643 ( .A1(n565), .A2(n596), .ZN(n582) );
  XOR2_X1 U644 ( .A(KEYINPUT33), .B(KEYINPUT69), .Z(n566) );
  XNOR2_X1 U645 ( .A(n567), .B(n566), .ZN(n627) );
  INV_X1 U646 ( .A(n627), .ZN(n568) );
  XNOR2_X1 U647 ( .A(n570), .B(KEYINPUT35), .ZN(n729) );
  INV_X1 U648 ( .A(n572), .ZN(n576) );
  INV_X1 U649 ( .A(n573), .ZN(n574) );
  NOR2_X1 U650 ( .A1(n574), .A2(n601), .ZN(n575) );
  NAND2_X1 U651 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U652 ( .A(KEYINPUT104), .B(n577), .ZN(n730) );
  AND2_X1 U653 ( .A1(n578), .A2(n604), .ZN(n579) );
  NAND2_X1 U654 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U655 ( .A(KEYINPUT101), .B(n581), .ZN(n661) );
  NOR2_X1 U656 ( .A1(n582), .A2(n604), .ZN(n608) );
  NAND2_X1 U657 ( .A1(n583), .A2(n608), .ZN(n584) );
  XNOR2_X1 U658 ( .A(n584), .B(KEYINPUT31), .ZN(n677) );
  NOR2_X1 U659 ( .A1(n661), .A2(n677), .ZN(n585) );
  AND2_X1 U660 ( .A1(n730), .A2(n349), .ZN(n587) );
  NOR2_X2 U661 ( .A1(n723), .A2(n710), .ZN(n640) );
  XOR2_X1 U662 ( .A(KEYINPUT2), .B(KEYINPUT83), .Z(n593) );
  NOR2_X1 U663 ( .A1(n593), .A2(KEYINPUT81), .ZN(n588) );
  OR2_X1 U664 ( .A1(n590), .A2(n588), .ZN(n592) );
  NOR2_X1 U665 ( .A1(KEYINPUT2), .A2(KEYINPUT81), .ZN(n589) );
  NAND2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U668 ( .A1(n593), .A2(KEYINPUT81), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n632) );
  XNOR2_X1 U670 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n598) );
  NOR2_X1 U671 ( .A1(n565), .A2(n596), .ZN(n597) );
  XNOR2_X1 U672 ( .A(n598), .B(n597), .ZN(n599) );
  XNOR2_X1 U673 ( .A(n599), .B(KEYINPUT116), .ZN(n607) );
  XOR2_X1 U674 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n603) );
  NAND2_X1 U675 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U676 ( .A(n603), .B(n602), .ZN(n605) );
  NOR2_X1 U677 ( .A1(n605), .A2(n509), .ZN(n606) );
  AND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n609) );
  NOR2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U680 ( .A(KEYINPUT51), .B(n610), .Z(n611) );
  NOR2_X1 U681 ( .A1(n626), .A2(n611), .ZN(n622) );
  NAND2_X1 U682 ( .A1(n612), .A2(n613), .ZN(n619) );
  NAND2_X1 U683 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U684 ( .A1(n617), .A2(n616), .ZN(n618) );
  AND2_X1 U685 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U686 ( .A1(n620), .A2(n627), .ZN(n621) );
  NOR2_X1 U687 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U688 ( .A(n623), .B(KEYINPUT52), .ZN(n624) );
  NOR2_X1 U689 ( .A1(n625), .A2(n624), .ZN(n629) );
  NOR2_X1 U690 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U691 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U692 ( .A(n630), .B(KEYINPUT118), .ZN(n631) );
  NAND2_X1 U693 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U694 ( .A1(G953), .A2(n633), .ZN(n636) );
  XNOR2_X1 U695 ( .A(n634), .B(KEYINPUT53), .ZN(n635) );
  XOR2_X1 U696 ( .A(G143), .B(n637), .Z(G45) );
  XOR2_X1 U697 ( .A(G134), .B(KEYINPUT113), .Z(n638) );
  XNOR2_X1 U698 ( .A(n639), .B(n638), .ZN(G36) );
  NOR2_X4 U699 ( .A1(n642), .A2(n641), .ZN(n697) );
  NAND2_X1 U700 ( .A1(n697), .A2(G472), .ZN(n646) );
  XOR2_X1 U701 ( .A(KEYINPUT107), .B(KEYINPUT62), .Z(n643) );
  XNOR2_X1 U702 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U703 ( .A(n646), .B(n645), .ZN(n648) );
  INV_X1 U704 ( .A(G952), .ZN(n647) );
  XOR2_X1 U705 ( .A(KEYINPUT108), .B(KEYINPUT63), .Z(n649) );
  XNOR2_X1 U706 ( .A(n650), .B(n649), .ZN(G57) );
  NAND2_X1 U707 ( .A1(n697), .A2(G210), .ZN(n656) );
  XNOR2_X1 U708 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n652) );
  XNOR2_X1 U709 ( .A(KEYINPUT55), .B(KEYINPUT82), .ZN(n651) );
  XNOR2_X1 U710 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U711 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U712 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U713 ( .A(KEYINPUT88), .B(KEYINPUT56), .ZN(n658) );
  XNOR2_X1 U714 ( .A(n659), .B(n658), .ZN(G51) );
  NAND2_X1 U715 ( .A1(n661), .A2(n673), .ZN(n660) );
  XNOR2_X1 U716 ( .A(n660), .B(G104), .ZN(G6) );
  XOR2_X1 U717 ( .A(KEYINPUT109), .B(KEYINPUT26), .Z(n663) );
  NAND2_X1 U718 ( .A1(n661), .A2(n676), .ZN(n662) );
  XNOR2_X1 U719 ( .A(n663), .B(n662), .ZN(n665) );
  XOR2_X1 U720 ( .A(G107), .B(KEYINPUT27), .Z(n664) );
  XNOR2_X1 U721 ( .A(n665), .B(n664), .ZN(G9) );
  XNOR2_X1 U722 ( .A(G110), .B(KEYINPUT110), .ZN(n667) );
  XNOR2_X1 U723 ( .A(n667), .B(n666), .ZN(G12) );
  XOR2_X1 U724 ( .A(G128), .B(KEYINPUT29), .Z(n669) );
  NAND2_X1 U725 ( .A1(n670), .A2(n676), .ZN(n668) );
  XNOR2_X1 U726 ( .A(n669), .B(n668), .ZN(G30) );
  XOR2_X1 U727 ( .A(G146), .B(KEYINPUT111), .Z(n672) );
  NAND2_X1 U728 ( .A1(n670), .A2(n673), .ZN(n671) );
  XNOR2_X1 U729 ( .A(n672), .B(n671), .ZN(G48) );
  NAND2_X1 U730 ( .A1(n677), .A2(n673), .ZN(n674) );
  XNOR2_X1 U731 ( .A(n674), .B(KEYINPUT112), .ZN(n675) );
  XNOR2_X1 U732 ( .A(G113), .B(n675), .ZN(G15) );
  NAND2_X1 U733 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U734 ( .A(n678), .B(G116), .ZN(G18) );
  XNOR2_X1 U735 ( .A(G125), .B(n679), .ZN(n680) );
  XNOR2_X1 U736 ( .A(n680), .B(KEYINPUT37), .ZN(G27) );
  BUF_X1 U737 ( .A(n697), .Z(n693) );
  NAND2_X1 U738 ( .A1(n693), .A2(G469), .ZN(n684) );
  XOR2_X1 U739 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n681) );
  XNOR2_X1 U740 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U741 ( .A1(n701), .A2(n685), .ZN(G54) );
  NAND2_X1 U742 ( .A1(n697), .A2(G475), .ZN(n690) );
  INV_X1 U743 ( .A(n686), .ZN(n688) );
  XOR2_X1 U744 ( .A(KEYINPUT59), .B(KEYINPUT91), .Z(n687) );
  XNOR2_X1 U745 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U746 ( .A(KEYINPUT60), .B(n692), .ZN(G60) );
  NAND2_X1 U747 ( .A1(n693), .A2(G478), .ZN(n694) );
  XNOR2_X1 U748 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U749 ( .A1(n701), .A2(n696), .ZN(G63) );
  NAND2_X1 U750 ( .A1(n697), .A2(G217), .ZN(n700) );
  XOR2_X1 U751 ( .A(n698), .B(KEYINPUT121), .Z(n699) );
  XNOR2_X1 U752 ( .A(n700), .B(n699), .ZN(n702) );
  XNOR2_X1 U753 ( .A(n703), .B(KEYINPUT122), .ZN(G66) );
  INV_X1 U754 ( .A(G898), .ZN(n709) );
  NAND2_X1 U755 ( .A1(n709), .A2(G953), .ZN(n705) );
  NAND2_X1 U756 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U757 ( .A(n706), .B(KEYINPUT124), .ZN(n715) );
  NAND2_X1 U758 ( .A1(G953), .A2(G224), .ZN(n707) );
  XOR2_X1 U759 ( .A(KEYINPUT61), .B(n707), .Z(n708) );
  NOR2_X1 U760 ( .A1(n709), .A2(n708), .ZN(n712) );
  NOR2_X1 U761 ( .A1(G953), .A2(n710), .ZN(n711) );
  NOR2_X1 U762 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U763 ( .A(n713), .B(KEYINPUT123), .Z(n714) );
  XNOR2_X1 U764 ( .A(n715), .B(n714), .ZN(G69) );
  XOR2_X1 U765 ( .A(KEYINPUT125), .B(n717), .Z(n718) );
  XNOR2_X1 U766 ( .A(n719), .B(n718), .ZN(n724) );
  XNOR2_X1 U767 ( .A(KEYINPUT126), .B(n724), .ZN(n720) );
  XNOR2_X1 U768 ( .A(G227), .B(n720), .ZN(n721) );
  NAND2_X1 U769 ( .A1(n721), .A2(G900), .ZN(n722) );
  NAND2_X1 U770 ( .A1(n722), .A2(G953), .ZN(n728) );
  XNOR2_X1 U771 ( .A(n723), .B(n724), .ZN(n726) );
  NAND2_X1 U772 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U773 ( .A1(n728), .A2(n727), .ZN(G72) );
  XNOR2_X1 U774 ( .A(G122), .B(n729), .ZN(G24) );
  XNOR2_X1 U775 ( .A(G101), .B(n730), .ZN(G3) );
  XNOR2_X1 U776 ( .A(G140), .B(KEYINPUT114), .ZN(n732) );
  XNOR2_X1 U777 ( .A(n732), .B(n731), .ZN(G42) );
  XNOR2_X1 U778 ( .A(G119), .B(KEYINPUT127), .ZN(n734) );
  XNOR2_X1 U779 ( .A(n734), .B(n733), .ZN(G21) );
  XOR2_X1 U780 ( .A(G137), .B(n735), .Z(G39) );
endmodule

