//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT74), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n190), .B2(KEYINPUT16), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G140), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(KEYINPUT74), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n189), .B1(new_n192), .B2(KEYINPUT73), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT73), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(G125), .A3(G140), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n194), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n187), .B1(new_n196), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(new_n199), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT16), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n203), .A2(G146), .A3(new_n191), .A4(new_n195), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  OR3_X1    g020(.A1(new_n206), .A2(KEYINPUT70), .A3(G128), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT70), .B1(new_n206), .B2(G128), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n207), .B(new_n208), .C1(G119), .C2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT24), .B(G110), .ZN(new_n211));
  OR2_X1    g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT23), .B1(new_n209), .B2(G119), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT71), .B1(new_n206), .B2(G128), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n213), .B(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT72), .ZN(new_n216));
  OAI21_X1  g030(.A(G110), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n218), .B1(new_n206), .B2(G128), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n219), .B(new_n214), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(KEYINPUT72), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n205), .B(new_n212), .C1(new_n217), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n210), .A2(new_n211), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n223), .B1(new_n220), .B2(G110), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n189), .A2(G125), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT75), .B1(new_n193), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n192), .A2(G140), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT75), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n190), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(G146), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n224), .A2(new_n204), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT22), .B(G137), .ZN(new_n233));
  INV_X1    g047(.A(G953), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(G221), .A3(G234), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n233), .B(new_n235), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n222), .A2(new_n232), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n236), .B1(new_n222), .B2(new_n232), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G902), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(KEYINPUT25), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n222), .A2(new_n232), .ZN(new_n242));
  INV_X1    g056(.A(new_n236), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n222), .A2(new_n232), .A3(new_n236), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n240), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT25), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n241), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G217), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(G234), .B2(new_n240), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n251), .A2(G902), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n249), .A2(new_n251), .B1(new_n239), .B2(new_n252), .ZN(new_n253));
  XOR2_X1   g067(.A(KEYINPUT26), .B(G101), .Z(new_n254));
  NOR2_X1   g068(.A1(G237), .A2(G953), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G210), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n254), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT11), .ZN(new_n261));
  INV_X1    g075(.A(G134), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n261), .B1(new_n262), .B2(G137), .ZN(new_n263));
  INV_X1    g077(.A(G137), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(KEYINPUT11), .A3(G134), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n262), .A2(G137), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G131), .ZN(new_n268));
  INV_X1    g082(.A(G131), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n263), .A2(new_n265), .A3(new_n269), .A4(new_n266), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n187), .A2(G143), .ZN(new_n272));
  INV_X1    g086(.A(G143), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G146), .ZN(new_n274));
  AND2_X1   g088(.A1(KEYINPUT0), .A2(G128), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(G143), .B(G146), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT0), .B(G128), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n271), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT65), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT1), .B1(new_n273), .B2(G146), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n273), .A2(G146), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n187), .A2(G143), .ZN(new_n285));
  OAI211_X1 g099(.A(G128), .B(new_n283), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n272), .B(new_n274), .C1(KEYINPUT1), .C2(new_n209), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT66), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n262), .A2(G137), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n264), .A2(G134), .ZN(new_n292));
  OAI21_X1  g106(.A(G131), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n270), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n286), .A2(KEYINPUT66), .A3(new_n287), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n290), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT64), .B1(new_n206), .B2(G116), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT64), .ZN(new_n299));
  INV_X1    g113(.A(G116), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n300), .A3(G119), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n300), .A2(G119), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G113), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT2), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G113), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n302), .A2(new_n304), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(new_n302), .B2(new_n304), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT65), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n271), .A2(new_n313), .A3(new_n280), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n282), .A2(new_n297), .A3(new_n312), .A4(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n312), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n279), .B1(new_n270), .B2(new_n268), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n288), .A2(new_n294), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT28), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n290), .A2(new_n295), .A3(new_n296), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n281), .A2(new_n312), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n320), .A2(KEYINPUT28), .B1(KEYINPUT68), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT68), .ZN(new_n326));
  AOI211_X1 g140(.A(new_n326), .B(new_n321), .C1(new_n315), .C2(new_n319), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n260), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n297), .A2(new_n314), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n317), .A2(new_n313), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT30), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT30), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n312), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n315), .A2(new_n259), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT31), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n335), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT31), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n282), .A2(new_n314), .A3(new_n297), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n332), .B1(new_n339), .B2(KEYINPUT30), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n337), .B(new_n338), .C1(new_n340), .C2(new_n312), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n328), .A2(new_n336), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT32), .ZN(new_n343));
  NOR2_X1   g157(.A1(G472), .A2(G902), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n343), .B1(new_n342), .B2(new_n344), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G472), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n339), .A2(new_n316), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n315), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT28), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n259), .A2(KEYINPUT29), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n324), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT69), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n324), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n350), .B2(KEYINPUT28), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(KEYINPUT69), .A3(new_n353), .ZN(new_n359));
  AOI21_X1  g173(.A(G902), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n334), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n315), .A3(new_n260), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n259), .B1(new_n325), .B2(new_n327), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n348), .B1(new_n360), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n253), .B1(new_n347), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(G214), .B1(G237), .B2(G902), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(G210), .B1(G237), .B2(G902), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n302), .A2(KEYINPUT5), .A3(new_n304), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT5), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n305), .B1(new_n303), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT3), .B1(new_n377), .B2(G107), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n379));
  INV_X1    g193(.A(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G104), .ZN(new_n381));
  INV_X1    g195(.A(G101), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n377), .A2(G107), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n378), .A2(new_n381), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n380), .A2(G104), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n377), .A2(G107), .ZN(new_n386));
  OAI21_X1  g200(.A(G101), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n303), .B1(new_n298), .B2(new_n301), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n309), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n376), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n378), .A2(new_n381), .A3(new_n383), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(G101), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n394), .B1(new_n310), .B2(new_n311), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(G101), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n396), .A2(KEYINPUT4), .A3(new_n384), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n391), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G110), .B(G122), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n391), .B(new_n399), .C1(new_n395), .C2(new_n397), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(KEYINPUT6), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n398), .A2(new_n404), .A3(new_n400), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n286), .A2(new_n192), .A3(new_n287), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n276), .B(G125), .C1(new_n277), .C2(new_n278), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G224), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(G953), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT81), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n408), .B(new_n411), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n403), .A2(new_n405), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT82), .B(KEYINPUT8), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n399), .B(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n373), .A2(new_n375), .B1(new_n389), .B2(new_n309), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT83), .B1(new_n417), .B2(new_n388), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n388), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n417), .A2(KEYINPUT83), .A3(new_n388), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n416), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n411), .A2(KEYINPUT84), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n411), .A2(KEYINPUT7), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n406), .A4(new_n407), .ZN(new_n425));
  OAI211_X1 g239(.A(KEYINPUT7), .B(new_n411), .C1(new_n408), .C2(KEYINPUT84), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n402), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n240), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n372), .B1(new_n413), .B2(new_n428), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n402), .A2(new_n425), .A3(new_n426), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT83), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n391), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n376), .A2(new_n390), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n384), .A2(new_n387), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n421), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n415), .ZN(new_n437));
  AOI21_X1  g251(.A(G902), .B1(new_n430), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n403), .A2(new_n405), .A3(new_n412), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(new_n371), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n370), .B1(new_n429), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G475), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n273), .A2(KEYINPUT85), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n443), .A2(G214), .A3(new_n255), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT85), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G143), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n446), .A2(new_n443), .B1(new_n255), .B2(G214), .ZN(new_n447));
  OAI211_X1 g261(.A(KEYINPUT17), .B(G131), .C1(new_n444), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT89), .ZN(new_n449));
  INV_X1    g263(.A(G214), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n450), .A2(G237), .A3(G953), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n443), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT85), .B(G143), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n452), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT89), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n454), .A2(new_n455), .A3(KEYINPUT17), .A4(G131), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G131), .B1(new_n444), .B2(new_n447), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n452), .B(new_n269), .C1(new_n451), .C2(new_n453), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT17), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n457), .A2(new_n201), .A3(new_n204), .A4(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n202), .A2(new_n187), .ZN(new_n463));
  NAND2_X1  g277(.A1(KEYINPUT18), .A2(G131), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  OAI22_X1  g279(.A1(new_n230), .A2(new_n463), .B1(new_n454), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT86), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n454), .A2(new_n468), .A3(new_n465), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n468), .B1(new_n454), .B2(new_n465), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(G113), .B(G122), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(new_n377), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(KEYINPUT88), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n462), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n461), .A2(new_n201), .A3(new_n204), .ZN(new_n477));
  INV_X1    g291(.A(new_n471), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n469), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n477), .A2(new_n457), .B1(new_n479), .B2(new_n467), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n476), .B1(new_n480), .B2(new_n474), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n442), .B1(new_n481), .B2(new_n240), .ZN(new_n482));
  NOR2_X1   g296(.A1(G475), .A2(G902), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT19), .B1(new_n226), .B2(new_n229), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n197), .A2(KEYINPUT19), .A3(new_n199), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n484), .A2(G146), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n204), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT87), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n458), .A2(new_n459), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT19), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n190), .A2(new_n227), .A3(new_n228), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n228), .B1(new_n190), .B2(new_n227), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(new_n187), .A3(new_n485), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT87), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n496), .A3(new_n204), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n489), .A2(new_n490), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n474), .B1(new_n498), .B2(new_n472), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n462), .A2(new_n472), .A3(new_n475), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n483), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT20), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT20), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n503), .B(new_n483), .C1(new_n499), .C2(new_n500), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n482), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT9), .B(G234), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT76), .ZN(new_n508));
  OR2_X1    g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n508), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n511), .A2(new_n250), .A3(G953), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G122), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G116), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n300), .A2(G122), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n516), .A3(new_n380), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT90), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT90), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n515), .A2(new_n516), .A3(new_n519), .A4(new_n380), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n273), .A2(G128), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n209), .A2(G143), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n522), .A3(new_n262), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n262), .B1(new_n521), .B2(new_n522), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n518), .B(new_n520), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT91), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT14), .B1(new_n514), .B2(G116), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n514), .A2(G116), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT14), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n531), .B1(new_n300), .B2(G122), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(KEYINPUT91), .A3(new_n516), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n534), .B1(new_n516), .B2(KEYINPUT14), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n529), .A2(KEYINPUT92), .A3(new_n531), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n530), .A2(new_n533), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n526), .B1(G107), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT13), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n521), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n273), .A2(KEYINPUT13), .A3(G128), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n541), .A3(new_n522), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n542), .A2(G134), .ZN(new_n543));
  INV_X1    g357(.A(new_n517), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n380), .B1(new_n515), .B2(new_n516), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n523), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n513), .B1(new_n538), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n537), .A2(G107), .ZN(new_n549));
  INV_X1    g363(.A(new_n525), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n550), .A2(new_n523), .B1(KEYINPUT90), .B2(new_n517), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n520), .A3(new_n551), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n543), .A2(new_n546), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n512), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G478), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(KEYINPUT15), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n240), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n558), .B1(new_n555), .B2(new_n240), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n506), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n552), .A2(new_n553), .A3(new_n512), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n512), .B1(new_n552), .B2(new_n553), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n240), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n557), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(KEYINPUT93), .A3(new_n559), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n234), .A2(G952), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(G234), .B2(G237), .ZN(new_n570));
  AOI211_X1 g384(.A(new_n240), .B(new_n234), .C1(G234), .C2(G237), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT21), .B(G898), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n441), .A2(new_n505), .A3(new_n568), .A4(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT80), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n288), .A2(new_n434), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n286), .A2(new_n384), .A3(new_n387), .A4(new_n287), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n580), .A2(KEYINPUT12), .A3(new_n271), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT12), .B1(new_n580), .B2(new_n271), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n384), .A2(new_n387), .A3(KEYINPUT10), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n290), .A2(new_n296), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n396), .A2(KEYINPUT4), .A3(new_n384), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(new_n280), .A3(new_n394), .ZN(new_n587));
  INV_X1    g401(.A(new_n271), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT10), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n579), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n585), .A2(new_n587), .A3(new_n588), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n234), .A2(G227), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(KEYINPUT77), .ZN(new_n593));
  XNOR2_X1  g407(.A(G110), .B(G140), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n577), .B1(new_n583), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n579), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n287), .A2(new_n286), .B1(new_n384), .B2(new_n387), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n271), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT12), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n580), .A2(KEYINPUT12), .A3(new_n271), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n604), .A2(KEYINPUT80), .A3(new_n591), .A4(new_n595), .ZN(new_n605));
  INV_X1    g419(.A(new_n595), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n392), .A2(G101), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n279), .B1(new_n607), .B2(new_n393), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n608), .A2(new_n586), .B1(new_n589), .B2(new_n579), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n588), .B1(new_n609), .B2(new_n585), .ZN(new_n610));
  INV_X1    g424(.A(new_n591), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n606), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n597), .A2(new_n605), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(G469), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n613), .A2(new_n614), .A3(new_n240), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n591), .B1(new_n581), .B2(new_n582), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT78), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n604), .A2(KEYINPUT78), .A3(new_n591), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(new_n606), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT79), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n596), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n610), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n591), .A2(KEYINPUT79), .A3(new_n595), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n620), .A2(G469), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(G469), .A2(G902), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n615), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(G221), .B1(new_n511), .B2(G902), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n576), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n368), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(new_n382), .ZN(G3));
  NAND2_X1  g448(.A1(new_n342), .A2(new_n240), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(G472), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n336), .A2(new_n341), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n320), .A2(KEYINPUT28), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n324), .A2(KEYINPUT68), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n320), .A2(KEYINPUT68), .A3(KEYINPUT28), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n259), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n344), .B1(new_n637), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n636), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n253), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n644), .A2(new_n645), .A3(new_n630), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n429), .A2(KEYINPUT94), .A3(new_n440), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n371), .B1(new_n438), .B2(new_n439), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT94), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n370), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT96), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n565), .B2(new_n556), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT95), .B1(new_n552), .B2(new_n553), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT33), .ZN(new_n655));
  OAI22_X1  g469(.A1(new_n563), .A2(new_n564), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT95), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n657), .B1(new_n538), .B2(new_n547), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n548), .A2(new_n658), .A3(KEYINPUT33), .A4(new_n554), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n556), .A2(G902), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n656), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n656), .A2(new_n659), .A3(new_n652), .A4(new_n660), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n505), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n646), .A2(new_n574), .A3(new_n651), .A4(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n666), .B(KEYINPUT97), .Z(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT34), .B(G104), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  AND3_X1   g483(.A1(new_n566), .A2(KEYINPUT93), .A3(new_n559), .ZN(new_n670));
  AOI21_X1  g484(.A(KEYINPUT93), .B1(new_n566), .B2(new_n559), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n505), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n647), .A2(new_n650), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n673), .A2(new_n674), .A3(new_n573), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n646), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT35), .B(G107), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  NAND2_X1  g492(.A1(new_n249), .A2(new_n251), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n243), .A2(KEYINPUT36), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n242), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n252), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n629), .A3(new_n628), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n644), .A2(new_n684), .A3(new_n575), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT37), .B(G110), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT98), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n685), .B(new_n687), .ZN(G12));
  AOI21_X1  g502(.A(KEYINPUT69), .B1(new_n358), .B2(new_n353), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n321), .B1(new_n349), .B2(new_n315), .ZN(new_n690));
  NOR4_X1   g504(.A1(new_n690), .A2(new_n355), .A3(new_n357), .A4(new_n352), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n240), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT29), .B1(new_n362), .B2(new_n363), .ZN(new_n693));
  OAI21_X1  g507(.A(G472), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n694), .B1(new_n346), .B2(new_n345), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n481), .A2(new_n240), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G475), .ZN(new_n697));
  INV_X1    g511(.A(new_n504), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n466), .B1(new_n478), .B2(new_n469), .ZN(new_n699));
  INV_X1    g513(.A(new_n490), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n495), .A2(new_n204), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n700), .B1(new_n701), .B2(KEYINPUT87), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n699), .B1(new_n702), .B2(new_n497), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n476), .B1(new_n703), .B2(new_n474), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n503), .B1(new_n704), .B2(new_n483), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n697), .B1(new_n698), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n568), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT99), .ZN(new_n708));
  INV_X1    g522(.A(G900), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n571), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n570), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n651), .A2(new_n707), .A3(new_n708), .A4(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n684), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n505), .A2(new_n672), .A3(new_n712), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT99), .B1(new_n715), .B2(new_n674), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n695), .A2(new_n713), .A3(new_n714), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G128), .ZN(G30));
  NAND2_X1  g532(.A1(new_n429), .A2(new_n440), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n719), .B(KEYINPUT38), .Z(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n505), .A2(new_n568), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n369), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n643), .A2(KEYINPUT32), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n260), .B1(new_n361), .B2(new_n315), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n240), .B1(new_n350), .B2(new_n259), .ZN(new_n728));
  OAI21_X1  g542(.A(G472), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n683), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n712), .B(KEYINPUT39), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n631), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n730), .B1(KEYINPUT40), .B2(new_n732), .ZN(new_n733));
  AOI211_X1 g547(.A(new_n723), .B(new_n733), .C1(KEYINPUT40), .C2(new_n732), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n273), .ZN(G45));
  INV_X1    g549(.A(new_n664), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n706), .A2(new_n736), .A3(new_n712), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n674), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n695), .A2(new_n714), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT100), .B(G146), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G48));
  NOR3_X1   g555(.A1(new_n505), .A2(new_n664), .A3(new_n573), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n253), .B(new_n742), .C1(new_n347), .C2(new_n367), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n613), .A2(new_n240), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(G469), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n629), .A3(new_n615), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT101), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT101), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n745), .A2(new_n748), .A3(new_n629), .A4(new_n615), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n747), .A2(new_n651), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT102), .B1(new_n743), .B2(new_n750), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n747), .A2(new_n651), .A3(new_n749), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n645), .B1(new_n726), .B2(new_n694), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT102), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n752), .A2(new_n753), .A3(new_n754), .A4(new_n742), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(KEYINPUT41), .B(G113), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G15));
  AND3_X1   g572(.A1(new_n695), .A2(new_n675), .A3(new_n253), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n747), .A2(new_n749), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(KEYINPUT103), .B(G116), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G18));
  NAND4_X1  g578(.A1(new_n683), .A2(new_n568), .A3(new_n574), .A4(new_n505), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n694), .B2(new_n726), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n752), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G119), .ZN(G21));
  NAND3_X1  g582(.A1(new_n651), .A2(new_n722), .A3(new_n574), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n348), .B1(new_n342), .B2(new_n240), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n260), .B1(new_n690), .B2(new_n357), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n336), .A3(new_n341), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(new_n344), .ZN(new_n774));
  NOR4_X1   g588(.A1(new_n645), .A2(new_n771), .A3(new_n774), .A4(KEYINPUT104), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT104), .ZN(new_n776));
  AOI22_X1  g590(.A1(new_n635), .A2(G472), .B1(new_n344), .B2(new_n773), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n776), .B1(new_n777), .B2(new_n253), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n761), .B(new_n770), .C1(new_n775), .C2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G122), .ZN(G24));
  AOI22_X1  g594(.A1(new_n249), .A2(new_n251), .B1(new_n252), .B2(new_n681), .ZN(new_n781));
  NOR4_X1   g595(.A1(new_n737), .A2(new_n771), .A3(new_n774), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n752), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G125), .ZN(G27));
  XOR2_X1   g598(.A(new_n627), .B(KEYINPUT105), .Z(new_n785));
  NAND3_X1  g599(.A1(new_n615), .A2(new_n626), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT106), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(new_n787), .A3(new_n629), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n429), .A2(new_n369), .A3(new_n440), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT107), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n429), .A2(KEYINPUT107), .A3(new_n369), .A4(new_n440), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n787), .B1(new_n786), .B2(new_n629), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n789), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n737), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n753), .A3(new_n797), .ZN(new_n798));
  XOR2_X1   g612(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT108), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(KEYINPUT42), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n796), .A2(new_n753), .A3(new_n797), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G131), .ZN(G33));
  INV_X1    g620(.A(new_n715), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n794), .A2(new_n795), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n753), .A2(new_n807), .A3(new_n788), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(new_n262), .ZN(G36));
  NOR2_X1   g624(.A1(new_n706), .A2(new_n664), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(KEYINPUT43), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(new_n644), .A3(new_n683), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT44), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n794), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(new_n814), .B2(new_n813), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n816), .A2(KEYINPUT109), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(KEYINPUT109), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT46), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n620), .A2(new_n625), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(KEYINPUT45), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n614), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(KEYINPUT45), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n785), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n819), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n822), .A2(new_n823), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(KEYINPUT46), .A3(new_n785), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n826), .A2(new_n615), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n629), .ZN(new_n830));
  INV_X1    g644(.A(new_n731), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n817), .A2(new_n818), .A3(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(G137), .ZN(G39));
  NOR4_X1   g648(.A1(new_n695), .A2(new_n253), .A3(new_n737), .A4(new_n794), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n835), .B(KEYINPUT110), .Z(new_n836));
  NAND3_X1  g650(.A1(new_n829), .A2(KEYINPUT47), .A3(new_n629), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT47), .B1(new_n829), .B2(new_n629), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  XOR2_X1   g654(.A(KEYINPUT111), .B(G140), .Z(new_n841));
  XNOR2_X1  g655(.A(new_n840), .B(new_n841), .ZN(G42));
  AND2_X1   g656(.A1(new_n812), .A2(new_n570), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n773), .A2(new_n344), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n636), .A2(new_n253), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT104), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n777), .A2(new_n776), .A3(new_n253), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n752), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n569), .B(KEYINPUT118), .Z(new_n851));
  INV_X1    g665(.A(new_n665), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n729), .B1(new_n345), .B2(new_n346), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n853), .A2(new_n645), .A3(new_n711), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n760), .A2(new_n794), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n850), .B(new_n851), .C1(new_n852), .C2(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n843), .A2(new_n855), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n753), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n859), .A2(KEYINPUT48), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(KEYINPUT48), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n857), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n856), .A2(new_n706), .A3(new_n736), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n771), .A2(new_n774), .A3(new_n781), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n863), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n721), .A2(new_n760), .A3(new_n369), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n849), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n867), .B1(new_n849), .B2(new_n868), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n865), .B(KEYINPUT51), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n849), .A2(new_n792), .A3(new_n793), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n838), .A2(new_n839), .ZN(new_n873));
  INV_X1    g687(.A(new_n629), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n745), .A2(new_n874), .A3(new_n615), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n872), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n862), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n869), .A2(new_n870), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT116), .B1(new_n838), .B2(new_n839), .ZN(new_n879));
  INV_X1    g693(.A(new_n839), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT116), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(new_n837), .A3(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n879), .A2(new_n882), .A3(new_n875), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n878), .B(new_n865), .C1(new_n883), .C2(new_n872), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT51), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n877), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n783), .A2(new_n717), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n706), .A2(new_n647), .A3(new_n672), .A4(new_n650), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n786), .A2(new_n629), .ZN(new_n889));
  INV_X1    g703(.A(new_n712), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(new_n781), .A3(new_n853), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n739), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT52), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n684), .B1(new_n726), .B2(new_n694), .ZN(new_n895));
  AOI22_X1  g709(.A1(new_n895), .A2(new_n738), .B1(new_n730), .B2(new_n891), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT52), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n896), .A2(new_n897), .A3(new_n717), .A4(new_n783), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT115), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT115), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n894), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n566), .A2(new_n559), .A3(new_n712), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n904), .B(new_n482), .C1(new_n502), .C2(new_n504), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(new_n792), .A3(new_n793), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT113), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT113), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n905), .A2(new_n792), .A3(new_n908), .A4(new_n793), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n907), .A2(new_n695), .A3(new_n714), .A4(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n808), .A2(new_n797), .A3(new_n864), .A4(new_n788), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI211_X1 g726(.A(new_n809), .B(new_n912), .C1(new_n800), .C2(new_n804), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n685), .B1(new_n759), .B2(new_n761), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n560), .A2(new_n561), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n706), .A2(new_n915), .A3(new_n573), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n646), .A2(new_n441), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n760), .A2(new_n769), .ZN(new_n918));
  AOI22_X1  g732(.A1(new_n848), .A2(new_n918), .B1(new_n766), .B2(new_n752), .ZN(new_n919));
  AND4_X1   g733(.A1(new_n756), .A2(new_n914), .A3(new_n917), .A4(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n630), .A2(new_n645), .ZN(new_n921));
  AOI22_X1  g735(.A1(new_n635), .A2(G472), .B1(new_n344), .B2(new_n342), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n921), .A2(new_n441), .A3(new_n922), .A4(new_n742), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n923), .B1(new_n368), .B2(new_n632), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT112), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n923), .B(KEYINPUT112), .C1(new_n368), .C2(new_n632), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n913), .A2(new_n920), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(KEYINPUT53), .B1(new_n903), .B2(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n779), .A2(new_n767), .A3(new_n917), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n928), .A2(new_n931), .A3(new_n756), .A4(new_n914), .ZN(new_n932));
  INV_X1    g746(.A(new_n809), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n805), .A2(new_n933), .A3(new_n911), .A4(new_n910), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT114), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT114), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n913), .A2(new_n920), .A3(new_n936), .A4(new_n928), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n899), .A2(KEYINPUT53), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n930), .A2(new_n939), .A3(KEYINPUT54), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT53), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n903), .B2(new_n929), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT54), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n894), .A2(new_n898), .A3(KEYINPUT53), .ZN(new_n944));
  OR3_X1    g758(.A1(new_n932), .A2(new_n934), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n886), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(G952), .A2(G953), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n745), .A2(new_n615), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT49), .Z(new_n951));
  NOR3_X1   g765(.A1(new_n645), .A2(new_n370), .A3(new_n874), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n951), .A2(new_n720), .A3(new_n811), .A4(new_n952), .ZN(new_n953));
  OAI22_X1  g767(.A1(new_n948), .A2(new_n949), .B1(new_n853), .B2(new_n953), .ZN(G75));
  NOR2_X1   g768(.A1(new_n234), .A2(G952), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT119), .Z(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n240), .B1(new_n942), .B2(new_n945), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT56), .B1(new_n958), .B2(G210), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n403), .A2(new_n405), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(new_n412), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT55), .Z(new_n962));
  OR2_X1    g776(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n959), .A2(new_n962), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n957), .B1(new_n963), .B2(new_n964), .ZN(G51));
  XOR2_X1   g779(.A(new_n785), .B(KEYINPUT57), .Z(new_n966));
  AND3_X1   g780(.A1(new_n894), .A2(new_n898), .A3(new_n901), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n901), .B1(new_n894), .B2(new_n898), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n932), .A2(new_n934), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT53), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n929), .A2(new_n944), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n971), .A2(KEYINPUT54), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n943), .B1(new_n942), .B2(new_n945), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n966), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n613), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n824), .B(KEYINPUT120), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n958), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n955), .B1(new_n976), .B2(new_n978), .ZN(G54));
  NAND3_X1  g793(.A1(new_n958), .A2(KEYINPUT58), .A3(G475), .ZN(new_n980));
  INV_X1    g794(.A(new_n704), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n982), .A2(new_n983), .A3(new_n955), .ZN(G60));
  NAND2_X1  g798(.A1(new_n656), .A2(new_n659), .ZN(new_n985));
  NAND2_X1  g799(.A1(G478), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT59), .Z(new_n987));
  NOR2_X1   g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT54), .B1(new_n971), .B2(new_n972), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(new_n946), .ZN(new_n991));
  OAI21_X1  g805(.A(KEYINPUT121), .B1(new_n991), .B2(new_n957), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n988), .B1(new_n973), .B2(new_n974), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT121), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n993), .A2(new_n994), .A3(new_n956), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n985), .B1(new_n947), .B2(new_n987), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n992), .A2(new_n995), .A3(new_n996), .ZN(G63));
  INV_X1    g811(.A(KEYINPUT122), .ZN(new_n998));
  NAND2_X1  g812(.A1(G217), .A2(G902), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT60), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(new_n942), .B2(new_n945), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n998), .B1(new_n1001), .B2(new_n681), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n1002), .A2(KEYINPUT61), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n957), .B1(new_n1001), .B2(new_n681), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n971), .A2(new_n972), .ZN(new_n1005));
  OAI22_X1  g819(.A1(new_n1005), .A2(new_n1000), .B1(new_n237), .B2(new_n238), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n1006), .B(new_n1004), .C1(new_n1002), .C2(KEYINPUT61), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(G66));
  OAI21_X1  g824(.A(G953), .B1(new_n572), .B2(new_n409), .ZN(new_n1011));
  INV_X1    g825(.A(new_n932), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1011), .B1(new_n1012), .B2(G953), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n960), .B1(G898), .B2(new_n234), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1013), .B(new_n1014), .ZN(G69));
  NAND2_X1  g829(.A1(new_n494), .A2(new_n485), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n340), .B(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n234), .B1(G227), .B2(G900), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n783), .A2(new_n717), .A3(new_n739), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n734), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT62), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n706), .A2(new_n915), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1022), .A2(new_n665), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT123), .Z(new_n1024));
  OR4_X1    g838(.A1(new_n368), .A2(new_n1024), .A3(new_n732), .A4(new_n794), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n1021), .A2(new_n833), .A3(new_n840), .A4(new_n1025), .ZN(new_n1026));
  AOI211_X1 g840(.A(new_n1017), .B(new_n1018), .C1(new_n1026), .C2(new_n234), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n709), .A2(G227), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n805), .A2(new_n933), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT124), .Z(new_n1030));
  NOR2_X1   g844(.A1(new_n368), .A2(new_n888), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1019), .B1(new_n832), .B2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g846(.A1(new_n1030), .A2(new_n833), .A3(new_n840), .A4(new_n1032), .ZN(new_n1033));
  MUX2_X1   g847(.A(new_n1028), .B(new_n1033), .S(new_n234), .Z(new_n1034));
  AOI21_X1  g848(.A(new_n1027), .B1(new_n1034), .B2(new_n1017), .ZN(G72));
  XNOR2_X1  g849(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n348), .A2(new_n240), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1038), .B1(new_n1026), .B2(new_n932), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n955), .B1(new_n1039), .B2(new_n727), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1038), .B1(new_n1033), .B2(new_n932), .ZN(new_n1041));
  XOR2_X1   g855(.A(new_n362), .B(KEYINPUT126), .Z(new_n1042));
  NAND2_X1  g856(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g857(.A(new_n727), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1044), .A2(new_n362), .A3(new_n1038), .ZN(new_n1045));
  XOR2_X1   g859(.A(new_n1045), .B(KEYINPUT127), .Z(new_n1046));
  NAND3_X1  g860(.A1(new_n930), .A2(new_n939), .A3(new_n1046), .ZN(new_n1047));
  AND3_X1   g861(.A1(new_n1040), .A2(new_n1043), .A3(new_n1047), .ZN(G57));
endmodule


