

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781;

  INV_X1 U375 ( .A(n689), .ZN(n354) );
  INV_X1 U376 ( .A(n689), .ZN(n358) );
  INV_X1 U377 ( .A(n689), .ZN(n362) );
  INV_X1 U378 ( .A(n660), .ZN(n356) );
  INV_X1 U379 ( .A(n672), .ZN(n360) );
  INV_X1 U380 ( .A(n687), .ZN(n364) );
  AND2_X1 U381 ( .A1(n431), .A2(n430), .ZN(n429) );
  AND2_X1 U382 ( .A1(n397), .A2(n396), .ZN(n395) );
  XNOR2_X1 U383 ( .A(n487), .B(n420), .ZN(n755) );
  XNOR2_X1 U384 ( .A(n425), .B(n478), .ZN(n767) );
  XNOR2_X1 U385 ( .A(n522), .B(n463), .ZN(n478) );
  INV_X1 U386 ( .A(n353), .ZN(n665) );
  NAND2_X1 U387 ( .A1(n355), .A2(n354), .ZN(n353) );
  XNOR2_X1 U388 ( .A(n661), .B(n356), .ZN(n355) );
  INV_X1 U389 ( .A(n357), .ZN(n676) );
  NAND2_X1 U390 ( .A1(n359), .A2(n358), .ZN(n357) );
  XNOR2_X1 U391 ( .A(n673), .B(n360), .ZN(n359) );
  INV_X1 U392 ( .A(n361), .ZN(n692) );
  NAND2_X1 U393 ( .A1(n363), .A2(n362), .ZN(n361) );
  XNOR2_X1 U394 ( .A(n688), .B(n364), .ZN(n363) );
  NOR2_X1 U395 ( .A1(n576), .A2(KEYINPUT44), .ZN(n419) );
  XOR2_X1 U396 ( .A(G125), .B(G146), .Z(n476) );
  OR2_X2 U397 ( .A1(n667), .A2(G902), .ZN(n410) );
  OR2_X2 U398 ( .A1(n659), .A2(G902), .ZN(n404) );
  NAND2_X2 U399 ( .A1(n378), .A2(n376), .ZN(n577) );
  XNOR2_X2 U400 ( .A(n499), .B(n435), .ZN(n677) );
  BUF_X1 U401 ( .A(n651), .Z(n693) );
  NAND2_X1 U402 ( .A1(n377), .A2(n370), .ZN(n376) );
  NAND2_X1 U403 ( .A1(n428), .A2(n427), .ZN(n426) );
  XNOR2_X1 U404 ( .A(n410), .B(n367), .ZN(n545) );
  XNOR2_X1 U405 ( .A(n516), .B(G134), .ZN(n425) );
  INV_X2 U406 ( .A(G953), .ZN(n464) );
  NOR2_X1 U407 ( .A1(n415), .A2(n413), .ZN(n412) );
  XOR2_X1 U408 ( .A(G119), .B(G110), .Z(n486) );
  XNOR2_X1 U409 ( .A(n409), .B(n407), .ZN(n521) );
  XNOR2_X1 U410 ( .A(KEYINPUT82), .B(KEYINPUT8), .ZN(n409) );
  NOR2_X1 U411 ( .A1(n408), .A2(G953), .ZN(n407) );
  INV_X1 U412 ( .A(G234), .ZN(n408) );
  AND2_X1 U413 ( .A1(n401), .A2(n559), .ZN(n400) );
  OR2_X1 U414 ( .A1(n677), .A2(n394), .ZN(n393) );
  NAND2_X1 U415 ( .A1(G469), .A2(n531), .ZN(n394) );
  XNOR2_X1 U416 ( .A(n446), .B(KEYINPUT25), .ZN(n447) );
  NAND2_X1 U417 ( .A1(n412), .A2(n411), .ZN(n424) );
  NAND2_X1 U418 ( .A1(n419), .A2(n418), .ZN(n411) );
  XNOR2_X1 U419 ( .A(n387), .B(n513), .ZN(n671) );
  XNOR2_X1 U420 ( .A(n518), .B(n514), .ZN(n387) );
  XNOR2_X1 U421 ( .A(n423), .B(n422), .ZN(n683) );
  XNOR2_X1 U422 ( .A(n477), .B(n481), .ZN(n422) );
  XNOR2_X1 U423 ( .A(n480), .B(n478), .ZN(n423) );
  XNOR2_X1 U424 ( .A(n549), .B(n548), .ZN(n728) );
  XNOR2_X1 U425 ( .A(n392), .B(n372), .ZN(n571) );
  AND2_X1 U426 ( .A1(n504), .A2(n622), .ZN(n392) );
  AND2_X1 U427 ( .A1(n591), .A2(n365), .ZN(n631) );
  NAND2_X1 U428 ( .A1(n375), .A2(n366), .ZN(n380) );
  AND2_X1 U429 ( .A1(n399), .A2(n400), .ZN(n374) );
  NOR2_X1 U430 ( .A1(G953), .A2(G237), .ZN(n506) );
  INV_X1 U431 ( .A(KEYINPUT15), .ZN(n442) );
  NAND2_X1 U432 ( .A1(n472), .A2(G902), .ZN(n396) );
  XNOR2_X1 U433 ( .A(G143), .B(G113), .ZN(n509) );
  XNOR2_X1 U434 ( .A(n383), .B(n382), .ZN(n717) );
  INV_X1 U435 ( .A(KEYINPUT115), .ZN(n382) );
  OR2_X1 U436 ( .A1(n696), .A2(n556), .ZN(n564) );
  XNOR2_X1 U437 ( .A(n540), .B(KEYINPUT0), .ZN(n583) );
  NOR2_X1 U438 ( .A1(n605), .A2(n539), .ZN(n540) );
  XNOR2_X1 U439 ( .A(n482), .B(KEYINPUT3), .ZN(n484) );
  INV_X1 U440 ( .A(KEYINPUT72), .ZN(n482) );
  XNOR2_X1 U441 ( .A(G101), .B(G104), .ZN(n469) );
  XNOR2_X1 U442 ( .A(n406), .B(n405), .ZN(n632) );
  INV_X1 U443 ( .A(KEYINPUT108), .ZN(n405) );
  NAND2_X1 U444 ( .A1(n631), .A2(n630), .ZN(n406) );
  NOR2_X1 U445 ( .A1(n579), .A2(n712), .ZN(n388) );
  NOR2_X1 U446 ( .A1(n474), .A2(n473), .ZN(n475) );
  OR2_X1 U447 ( .A1(n570), .A2(n569), .ZN(n599) );
  AND2_X2 U448 ( .A1(n545), .A2(n695), .ZN(n699) );
  INV_X1 U449 ( .A(n578), .ZN(n402) );
  XNOR2_X1 U450 ( .A(n579), .B(n557), .ZN(n591) );
  XNOR2_X1 U451 ( .A(n441), .B(n768), .ZN(n667) );
  XNOR2_X1 U452 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U453 ( .A(n686), .B(n685), .ZN(n687) );
  NOR2_X1 U454 ( .A1(n464), .A2(G952), .ZN(n689) );
  XNOR2_X1 U455 ( .A(n555), .B(KEYINPUT42), .ZN(n596) );
  NAND2_X1 U456 ( .A1(n379), .A2(n561), .ZN(n378) );
  NAND2_X1 U457 ( .A1(n380), .A2(n374), .ZN(n379) );
  BUF_X1 U458 ( .A(n556), .Z(n389) );
  AND2_X1 U459 ( .A1(n600), .A2(n747), .ZN(n365) );
  AND2_X1 U460 ( .A1(n402), .A2(n403), .ZN(n366) );
  XOR2_X1 U461 ( .A(n448), .B(n447), .Z(n367) );
  AND2_X1 U462 ( .A1(n562), .A2(n579), .ZN(n368) );
  NAND2_X1 U463 ( .A1(n502), .A2(G210), .ZN(n369) );
  AND2_X1 U464 ( .A1(n400), .A2(n398), .ZN(n370) );
  XNOR2_X1 U465 ( .A(KEYINPUT91), .B(KEYINPUT33), .ZN(n371) );
  XOR2_X1 U466 ( .A(n505), .B(KEYINPUT73), .Z(n372) );
  XOR2_X1 U467 ( .A(n503), .B(KEYINPUT30), .Z(n373) );
  INV_X1 U468 ( .A(KEYINPUT75), .ZN(n432) );
  INV_X1 U469 ( .A(KEYINPUT34), .ZN(n403) );
  XNOR2_X1 U470 ( .A(n442), .B(G902), .ZN(n646) );
  INV_X1 U471 ( .A(n711), .ZN(n375) );
  AND2_X1 U472 ( .A1(n380), .A2(n399), .ZN(n377) );
  AND2_X1 U473 ( .A1(n757), .A2(n646), .ZN(n645) );
  XNOR2_X2 U474 ( .A(n424), .B(n594), .ZN(n757) );
  NAND2_X1 U475 ( .A1(n381), .A2(n650), .ZN(n384) );
  NOR2_X1 U476 ( .A1(n649), .A2(n648), .ZN(n381) );
  XNOR2_X1 U477 ( .A(n388), .B(n373), .ZN(n620) );
  NOR2_X1 U478 ( .A1(n713), .A2(n712), .ZN(n383) );
  INV_X1 U479 ( .A(G104), .ZN(n485) );
  NAND2_X1 U480 ( .A1(n384), .A2(n653), .ZN(n654) );
  XNOR2_X1 U481 ( .A(n385), .B(n629), .ZN(n639) );
  NAND2_X1 U482 ( .A1(n626), .A2(n627), .ZN(n385) );
  NAND2_X1 U483 ( .A1(n386), .A2(n428), .ZN(n752) );
  XNOR2_X1 U484 ( .A(n604), .B(KEYINPUT36), .ZN(n386) );
  NAND2_X2 U485 ( .A1(n395), .A2(n393), .ZN(n546) );
  OR2_X2 U486 ( .A1(n571), .A2(n599), .ZN(n573) );
  XNOR2_X1 U487 ( .A(n755), .B(n683), .ZN(n488) );
  XNOR2_X1 U488 ( .A(n515), .B(n433), .ZN(n421) );
  XNOR2_X1 U489 ( .A(n497), .B(n421), .ZN(n420) );
  XNOR2_X2 U490 ( .A(n390), .B(n371), .ZN(n711) );
  NAND2_X1 U491 ( .A1(n704), .A2(n591), .ZN(n390) );
  NAND2_X1 U492 ( .A1(n391), .A2(n590), .ZN(n568) );
  XNOR2_X1 U493 ( .A(n566), .B(KEYINPUT79), .ZN(n391) );
  XNOR2_X2 U494 ( .A(n573), .B(n572), .ZN(n595) );
  XNOR2_X2 U495 ( .A(n546), .B(KEYINPUT1), .ZN(n556) );
  NAND2_X1 U496 ( .A1(n677), .A2(n472), .ZN(n397) );
  INV_X1 U497 ( .A(n561), .ZN(n398) );
  NAND2_X1 U498 ( .A1(n711), .A2(KEYINPUT34), .ZN(n399) );
  NAND2_X1 U499 ( .A1(n578), .A2(KEYINPUT34), .ZN(n401) );
  XNOR2_X2 U500 ( .A(n404), .B(n501), .ZN(n579) );
  XNOR2_X1 U501 ( .A(n499), .B(n498), .ZN(n659) );
  XNOR2_X2 U502 ( .A(n767), .B(G146), .ZN(n499) );
  INV_X1 U503 ( .A(n591), .ZN(n601) );
  NAND2_X1 U504 ( .A1(n414), .A2(n737), .ZN(n413) );
  NAND2_X1 U505 ( .A1(n576), .A2(KEYINPUT44), .ZN(n414) );
  NAND2_X1 U506 ( .A1(n417), .A2(n416), .ZN(n415) );
  NAND2_X1 U507 ( .A1(n577), .A2(KEYINPUT44), .ZN(n416) );
  NAND2_X1 U508 ( .A1(n589), .A2(n609), .ZN(n417) );
  INV_X1 U509 ( .A(n577), .ZN(n418) );
  OR2_X1 U510 ( .A1(n699), .A2(n432), .ZN(n430) );
  NAND2_X2 U511 ( .A1(n429), .A2(n426), .ZN(n704) );
  AND2_X1 U512 ( .A1(n699), .A2(n432), .ZN(n427) );
  INV_X1 U513 ( .A(n556), .ZN(n428) );
  NAND2_X1 U514 ( .A1(n556), .A2(KEYINPUT75), .ZN(n431) );
  AND2_X2 U515 ( .A1(n658), .A2(n657), .ZN(n434) );
  XNOR2_X2 U516 ( .A(n462), .B(G131), .ZN(n516) );
  XNOR2_X2 U517 ( .A(n654), .B(KEYINPUT65), .ZN(n682) );
  XNOR2_X1 U518 ( .A(G116), .B(G107), .ZN(n433) );
  XOR2_X1 U519 ( .A(n471), .B(n470), .Z(n435) );
  INV_X1 U520 ( .A(n476), .ZN(n477) );
  NAND2_X1 U521 ( .A1(n538), .A2(n459), .ZN(n539) );
  BUF_X1 U522 ( .A(n767), .Z(n769) );
  XNOR2_X1 U523 ( .A(n603), .B(n535), .ZN(n605) );
  NAND2_X1 U524 ( .A1(G221), .A2(n521), .ZN(n437) );
  XOR2_X1 U525 ( .A(KEYINPUT94), .B(KEYINPUT23), .Z(n436) );
  XNOR2_X1 U526 ( .A(n437), .B(n436), .ZN(n440) );
  XNOR2_X1 U527 ( .A(G128), .B(KEYINPUT24), .ZN(n438) );
  XNOR2_X1 U528 ( .A(n438), .B(n486), .ZN(n439) );
  XNOR2_X1 U529 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U530 ( .A(KEYINPUT10), .B(n476), .Z(n514) );
  XNOR2_X1 U531 ( .A(G137), .B(G140), .ZN(n466) );
  XNOR2_X1 U532 ( .A(n514), .B(n466), .ZN(n768) );
  INV_X1 U533 ( .A(n646), .ZN(n443) );
  NAND2_X1 U534 ( .A1(n443), .A2(G234), .ZN(n444) );
  XNOR2_X1 U535 ( .A(n444), .B(KEYINPUT96), .ZN(n445) );
  XNOR2_X1 U536 ( .A(KEYINPUT20), .B(n445), .ZN(n449) );
  NAND2_X1 U537 ( .A1(G217), .A2(n449), .ZN(n448) );
  XNOR2_X1 U538 ( .A(KEYINPUT95), .B(KEYINPUT97), .ZN(n446) );
  NAND2_X1 U539 ( .A1(n449), .A2(G221), .ZN(n450) );
  XNOR2_X1 U540 ( .A(n450), .B(KEYINPUT21), .ZN(n452) );
  INV_X1 U541 ( .A(KEYINPUT98), .ZN(n451) );
  XNOR2_X1 U542 ( .A(n452), .B(n451), .ZN(n695) );
  NAND2_X1 U543 ( .A1(G237), .A2(G234), .ZN(n453) );
  XOR2_X1 U544 ( .A(KEYINPUT14), .B(n453), .Z(n725) );
  NAND2_X1 U545 ( .A1(G953), .A2(G902), .ZN(n454) );
  NOR2_X1 U546 ( .A1(n725), .A2(n454), .ZN(n455) );
  XOR2_X1 U547 ( .A(n455), .B(KEYINPUT107), .Z(n457) );
  INV_X1 U548 ( .A(G900), .ZN(n456) );
  NAND2_X1 U549 ( .A1(n457), .A2(n456), .ZN(n461) );
  INV_X1 U550 ( .A(n725), .ZN(n459) );
  NAND2_X1 U551 ( .A1(G952), .A2(n464), .ZN(n537) );
  INV_X1 U552 ( .A(n537), .ZN(n458) );
  NAND2_X1 U553 ( .A1(n459), .A2(n458), .ZN(n460) );
  NAND2_X1 U554 ( .A1(n461), .A2(n460), .ZN(n550) );
  NAND2_X1 U555 ( .A1(n699), .A2(n550), .ZN(n474) );
  XNOR2_X2 U556 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n462) );
  XNOR2_X2 U557 ( .A(G143), .B(G128), .ZN(n522) );
  XNOR2_X1 U558 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n463) );
  NAND2_X1 U559 ( .A1(n464), .A2(G227), .ZN(n465) );
  XNOR2_X1 U560 ( .A(n465), .B(KEYINPUT77), .ZN(n467) );
  XNOR2_X1 U561 ( .A(n467), .B(n466), .ZN(n471) );
  XNOR2_X1 U562 ( .A(G110), .B(G107), .ZN(n468) );
  XNOR2_X1 U563 ( .A(n469), .B(n468), .ZN(n470) );
  INV_X1 U564 ( .A(G469), .ZN(n472) );
  BUF_X1 U565 ( .A(n546), .Z(n473) );
  XNOR2_X1 U566 ( .A(n475), .B(KEYINPUT76), .ZN(n622) );
  NAND2_X1 U567 ( .A1(G224), .A2(n464), .ZN(n479) );
  XNOR2_X1 U568 ( .A(n479), .B(KEYINPUT18), .ZN(n480) );
  XNOR2_X1 U569 ( .A(KEYINPUT17), .B(KEYINPUT93), .ZN(n481) );
  XNOR2_X1 U570 ( .A(G113), .B(G101), .ZN(n483) );
  XNOR2_X1 U571 ( .A(n484), .B(n483), .ZN(n497) );
  XNOR2_X1 U572 ( .A(n485), .B(G122), .ZN(n515) );
  XOR2_X1 U573 ( .A(n486), .B(KEYINPUT16), .Z(n487) );
  NAND2_X1 U574 ( .A1(n488), .A2(n443), .ZN(n490) );
  INV_X1 U575 ( .A(G902), .ZN(n531) );
  INV_X1 U576 ( .A(G237), .ZN(n489) );
  NAND2_X1 U577 ( .A1(n531), .A2(n489), .ZN(n502) );
  XNOR2_X2 U578 ( .A(n490), .B(n369), .ZN(n616) );
  INV_X1 U579 ( .A(KEYINPUT38), .ZN(n491) );
  XNOR2_X1 U580 ( .A(n616), .B(n491), .ZN(n713) );
  NAND2_X1 U581 ( .A1(n506), .A2(G210), .ZN(n493) );
  XNOR2_X1 U582 ( .A(G119), .B(G116), .ZN(n492) );
  XNOR2_X1 U583 ( .A(n493), .B(n492), .ZN(n495) );
  XNOR2_X1 U584 ( .A(KEYINPUT5), .B(G137), .ZN(n494) );
  XNOR2_X1 U585 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U586 ( .A(n497), .B(n496), .ZN(n498) );
  INV_X1 U587 ( .A(KEYINPUT74), .ZN(n500) );
  XNOR2_X1 U588 ( .A(n500), .B(G472), .ZN(n501) );
  NAND2_X1 U589 ( .A1(n502), .A2(G214), .ZN(n630) );
  INV_X1 U590 ( .A(n630), .ZN(n712) );
  INV_X1 U591 ( .A(KEYINPUT111), .ZN(n503) );
  NOR2_X1 U592 ( .A1(n713), .A2(n620), .ZN(n504) );
  XNOR2_X1 U593 ( .A(KEYINPUT88), .B(KEYINPUT39), .ZN(n505) );
  XOR2_X1 U594 ( .A(KEYINPUT11), .B(KEYINPUT100), .Z(n508) );
  NAND2_X1 U595 ( .A1(n506), .A2(G214), .ZN(n507) );
  XNOR2_X1 U596 ( .A(n508), .B(n507), .ZN(n512) );
  XOR2_X1 U597 ( .A(KEYINPUT101), .B(KEYINPUT12), .Z(n510) );
  XNOR2_X1 U598 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U599 ( .A(n512), .B(n511), .Z(n513) );
  XNOR2_X1 U600 ( .A(n515), .B(G140), .ZN(n517) );
  XNOR2_X1 U601 ( .A(n516), .B(n517), .ZN(n518) );
  NAND2_X1 U602 ( .A1(n671), .A2(n531), .ZN(n520) );
  XNOR2_X1 U603 ( .A(KEYINPUT13), .B(G475), .ZN(n519) );
  XNOR2_X1 U604 ( .A(n520), .B(n519), .ZN(n570) );
  NAND2_X1 U605 ( .A1(G217), .A2(n521), .ZN(n524) );
  XNOR2_X1 U606 ( .A(n522), .B(n433), .ZN(n523) );
  XNOR2_X1 U607 ( .A(n524), .B(n523), .ZN(n530) );
  XOR2_X1 U608 ( .A(KEYINPUT7), .B(KEYINPUT103), .Z(n526) );
  XNOR2_X1 U609 ( .A(G122), .B(KEYINPUT102), .ZN(n525) );
  XNOR2_X1 U610 ( .A(n526), .B(n525), .ZN(n528) );
  XOR2_X1 U611 ( .A(G134), .B(KEYINPUT9), .Z(n527) );
  XNOR2_X1 U612 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U613 ( .A(n530), .B(n529), .ZN(n655) );
  NAND2_X1 U614 ( .A1(n655), .A2(n531), .ZN(n533) );
  INV_X1 U615 ( .A(G478), .ZN(n532) );
  XNOR2_X1 U616 ( .A(n533), .B(n532), .ZN(n541) );
  INV_X1 U617 ( .A(n541), .ZN(n569) );
  AND2_X1 U618 ( .A1(n570), .A2(n569), .ZN(n749) );
  INV_X1 U619 ( .A(n749), .ZN(n587) );
  OR2_X1 U620 ( .A1(n571), .A2(n587), .ZN(n637) );
  XNOR2_X1 U621 ( .A(n637), .B(G134), .ZN(G36) );
  INV_X1 U622 ( .A(n616), .ZN(n534) );
  NAND2_X1 U623 ( .A1(n534), .A2(n630), .ZN(n603) );
  XNOR2_X1 U624 ( .A(KEYINPUT19), .B(KEYINPUT67), .ZN(n535) );
  NOR2_X1 U625 ( .A1(G898), .A2(n464), .ZN(n756) );
  NAND2_X1 U626 ( .A1(G902), .A2(n756), .ZN(n536) );
  NAND2_X1 U627 ( .A1(n537), .A2(n536), .ZN(n538) );
  AND2_X1 U628 ( .A1(n570), .A2(n541), .ZN(n714) );
  AND2_X1 U629 ( .A1(n695), .A2(n714), .ZN(n542) );
  NAND2_X1 U630 ( .A1(n583), .A2(n542), .ZN(n544) );
  INV_X1 U631 ( .A(KEYINPUT22), .ZN(n543) );
  XNOR2_X2 U632 ( .A(n544), .B(n543), .ZN(n590) );
  INV_X1 U633 ( .A(n545), .ZN(n562) );
  AND2_X1 U634 ( .A1(n590), .A2(n368), .ZN(n547) );
  NAND2_X1 U635 ( .A1(n547), .A2(n389), .ZN(n574) );
  XNOR2_X1 U636 ( .A(n574), .B(G110), .ZN(G12) );
  AND2_X1 U637 ( .A1(n717), .A2(n714), .ZN(n549) );
  INV_X1 U638 ( .A(KEYINPUT41), .ZN(n548) );
  AND2_X1 U639 ( .A1(n695), .A2(n550), .ZN(n551) );
  AND2_X1 U640 ( .A1(n562), .A2(n551), .ZN(n600) );
  INV_X1 U641 ( .A(n579), .ZN(n703) );
  NAND2_X1 U642 ( .A1(n600), .A2(n703), .ZN(n553) );
  XNOR2_X1 U643 ( .A(KEYINPUT113), .B(KEYINPUT28), .ZN(n552) );
  XNOR2_X1 U644 ( .A(n553), .B(n552), .ZN(n606) );
  INV_X1 U645 ( .A(n473), .ZN(n585) );
  AND2_X1 U646 ( .A1(n606), .A2(n585), .ZN(n554) );
  NAND2_X1 U647 ( .A1(n728), .A2(n554), .ZN(n555) );
  XNOR2_X1 U648 ( .A(n596), .B(G137), .ZN(G39) );
  XNOR2_X1 U649 ( .A(KEYINPUT104), .B(KEYINPUT6), .ZN(n557) );
  INV_X1 U650 ( .A(n583), .ZN(n578) );
  INV_X1 U651 ( .A(n570), .ZN(n558) );
  NAND2_X1 U652 ( .A1(n558), .A2(n569), .ZN(n618) );
  INV_X1 U653 ( .A(n618), .ZN(n559) );
  INV_X1 U654 ( .A(KEYINPUT85), .ZN(n560) );
  XNOR2_X1 U655 ( .A(n560), .B(KEYINPUT35), .ZN(n561) );
  XOR2_X1 U656 ( .A(n577), .B(G122), .Z(G24) );
  XNOR2_X1 U657 ( .A(n562), .B(KEYINPUT105), .ZN(n696) );
  INV_X1 U658 ( .A(KEYINPUT106), .ZN(n563) );
  XNOR2_X1 U659 ( .A(n564), .B(n563), .ZN(n565) );
  NAND2_X1 U660 ( .A1(n565), .A2(n601), .ZN(n566) );
  XNOR2_X1 U661 ( .A(KEYINPUT78), .B(KEYINPUT32), .ZN(n567) );
  XNOR2_X2 U662 ( .A(n568), .B(n567), .ZN(n575) );
  XNOR2_X1 U663 ( .A(n575), .B(G119), .ZN(G21) );
  XNOR2_X1 U664 ( .A(KEYINPUT114), .B(KEYINPUT40), .ZN(n572) );
  XNOR2_X1 U665 ( .A(n595), .B(G131), .ZN(G33) );
  NAND2_X1 U666 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U667 ( .A1(n578), .A2(n579), .ZN(n580) );
  NAND2_X1 U668 ( .A1(n704), .A2(n580), .ZN(n582) );
  XOR2_X1 U669 ( .A(KEYINPUT31), .B(KEYINPUT99), .Z(n581) );
  XNOR2_X1 U670 ( .A(n582), .B(n581), .ZN(n750) );
  NAND2_X1 U671 ( .A1(n699), .A2(n402), .ZN(n584) );
  NOR2_X1 U672 ( .A1(n584), .A2(n703), .ZN(n586) );
  AND2_X1 U673 ( .A1(n586), .A2(n585), .ZN(n739) );
  OR2_X1 U674 ( .A1(n750), .A2(n739), .ZN(n589) );
  NAND2_X1 U675 ( .A1(n587), .A2(n599), .ZN(n716) );
  INV_X1 U676 ( .A(KEYINPUT81), .ZN(n588) );
  XNOR2_X1 U677 ( .A(n716), .B(n588), .ZN(n609) );
  NAND2_X1 U678 ( .A1(n696), .A2(n590), .ZN(n592) );
  NOR2_X1 U679 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U680 ( .A1(n593), .A2(n389), .ZN(n737) );
  XNOR2_X1 U681 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n594) );
  NAND2_X1 U682 ( .A1(n596), .A2(n595), .ZN(n598) );
  XNOR2_X1 U683 ( .A(KEYINPUT87), .B(KEYINPUT46), .ZN(n597) );
  XNOR2_X1 U684 ( .A(n598), .B(n597), .ZN(n627) );
  INV_X1 U685 ( .A(n599), .ZN(n747) );
  XOR2_X1 U686 ( .A(KEYINPUT116), .B(n631), .Z(n602) );
  NOR2_X1 U687 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U688 ( .A1(n605), .A2(n473), .ZN(n607) );
  AND2_X1 U689 ( .A1(n607), .A2(n606), .ZN(n745) );
  NAND2_X1 U690 ( .A1(n745), .A2(n716), .ZN(n608) );
  NAND2_X1 U691 ( .A1(n608), .A2(KEYINPUT47), .ZN(n614) );
  INV_X1 U692 ( .A(n609), .ZN(n611) );
  XOR2_X1 U693 ( .A(KEYINPUT47), .B(KEYINPUT69), .Z(n610) );
  NOR2_X1 U694 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U695 ( .A1(n745), .A2(n612), .ZN(n613) );
  AND2_X1 U696 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U697 ( .A1(n752), .A2(n615), .ZN(n625) );
  BUF_X1 U698 ( .A(n616), .Z(n617) );
  OR2_X1 U699 ( .A1(n617), .A2(n618), .ZN(n619) );
  NOR2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n624) );
  INV_X1 U702 ( .A(KEYINPUT112), .ZN(n623) );
  XNOR2_X1 U703 ( .A(n624), .B(n623), .ZN(n780) );
  NOR2_X1 U704 ( .A1(n625), .A2(n780), .ZN(n626) );
  INV_X1 U705 ( .A(KEYINPUT86), .ZN(n628) );
  XNOR2_X1 U706 ( .A(n628), .B(KEYINPUT48), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n632), .A2(n389), .ZN(n634) );
  XOR2_X1 U708 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n633) );
  XNOR2_X1 U709 ( .A(n634), .B(n633), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n635), .A2(n617), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n636), .B(KEYINPUT110), .ZN(n778) );
  AND2_X1 U712 ( .A1(n778), .A2(n637), .ZN(n638) );
  AND2_X2 U713 ( .A1(n639), .A2(n638), .ZN(n770) );
  NAND2_X1 U714 ( .A1(n757), .A2(n770), .ZN(n651) );
  OR2_X1 U715 ( .A1(KEYINPUT83), .A2(n443), .ZN(n640) );
  NOR2_X1 U716 ( .A1(n651), .A2(n640), .ZN(n643) );
  AND2_X1 U717 ( .A1(KEYINPUT2), .A2(KEYINPUT66), .ZN(n641) );
  AND2_X1 U718 ( .A1(n646), .A2(n641), .ZN(n642) );
  NOR2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n650) );
  NAND2_X1 U720 ( .A1(n770), .A2(KEYINPUT83), .ZN(n644) );
  NOR2_X1 U721 ( .A1(n645), .A2(n644), .ZN(n649) );
  AND2_X1 U722 ( .A1(n646), .A2(KEYINPUT2), .ZN(n647) );
  NOR2_X1 U723 ( .A1(n647), .A2(KEYINPUT66), .ZN(n648) );
  INV_X1 U724 ( .A(n693), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n652), .A2(KEYINPUT2), .ZN(n653) );
  NAND2_X1 U726 ( .A1(n682), .A2(G478), .ZN(n656) );
  XNOR2_X1 U727 ( .A(n656), .B(n655), .ZN(n658) );
  INV_X1 U728 ( .A(n689), .ZN(n657) );
  XNOR2_X1 U729 ( .A(n434), .B(KEYINPUT124), .ZN(G63) );
  NAND2_X1 U730 ( .A1(n682), .A2(G472), .ZN(n661) );
  XNOR2_X1 U731 ( .A(n659), .B(KEYINPUT62), .ZN(n660) );
  XNOR2_X1 U732 ( .A(KEYINPUT92), .B(KEYINPUT63), .ZN(n663) );
  XNOR2_X1 U733 ( .A(n663), .B(KEYINPUT89), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n665), .B(n664), .ZN(G57) );
  BUF_X1 U735 ( .A(n682), .Z(n666) );
  NAND2_X1 U736 ( .A1(n666), .A2(G217), .ZN(n668) );
  XNOR2_X1 U737 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X1 U738 ( .A1(n669), .A2(n689), .ZN(G66) );
  NAND2_X1 U739 ( .A1(n682), .A2(G475), .ZN(n673) );
  XOR2_X1 U740 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n670) );
  XNOR2_X1 U741 ( .A(KEYINPUT68), .B(KEYINPUT60), .ZN(n675) );
  XNOR2_X1 U742 ( .A(n676), .B(n675), .ZN(G60) );
  NAND2_X1 U743 ( .A1(n666), .A2(G469), .ZN(n680) );
  XOR2_X1 U744 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n678) );
  XNOR2_X1 U745 ( .A(n677), .B(n678), .ZN(n679) );
  XNOR2_X1 U746 ( .A(n680), .B(n679), .ZN(n681) );
  NOR2_X1 U747 ( .A1(n681), .A2(n689), .ZN(G54) );
  NAND2_X1 U748 ( .A1(n682), .A2(G210), .ZN(n688) );
  XOR2_X1 U749 ( .A(n683), .B(n755), .Z(n686) );
  XNOR2_X1 U750 ( .A(KEYINPUT90), .B(KEYINPUT54), .ZN(n684) );
  XOR2_X1 U751 ( .A(n684), .B(KEYINPUT55), .Z(n685) );
  XNOR2_X1 U752 ( .A(KEYINPUT122), .B(KEYINPUT56), .ZN(n691) );
  XNOR2_X1 U753 ( .A(n692), .B(n691), .ZN(G51) );
  NAND2_X1 U754 ( .A1(n693), .A2(KEYINPUT80), .ZN(n694) );
  XNOR2_X1 U755 ( .A(n694), .B(KEYINPUT2), .ZN(n735) );
  NOR2_X1 U756 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U757 ( .A(KEYINPUT49), .B(n697), .Z(n698) );
  NOR2_X1 U758 ( .A1(n698), .A2(n703), .ZN(n702) );
  NOR2_X1 U759 ( .A1(n699), .A2(n428), .ZN(n700) );
  XOR2_X1 U760 ( .A(KEYINPUT50), .B(n700), .Z(n701) );
  NAND2_X1 U761 ( .A1(n702), .A2(n701), .ZN(n706) );
  NAND2_X1 U762 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U763 ( .A1(n706), .A2(n705), .ZN(n708) );
  XOR2_X1 U764 ( .A(KEYINPUT51), .B(KEYINPUT120), .Z(n707) );
  XNOR2_X1 U765 ( .A(n708), .B(n707), .ZN(n709) );
  NAND2_X1 U766 ( .A1(n728), .A2(n709), .ZN(n710) );
  XOR2_X1 U767 ( .A(KEYINPUT121), .B(n710), .Z(n722) );
  INV_X1 U768 ( .A(n711), .ZN(n729) );
  NAND2_X1 U769 ( .A1(n713), .A2(n712), .ZN(n715) );
  NAND2_X1 U770 ( .A1(n715), .A2(n714), .ZN(n719) );
  NAND2_X1 U771 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U772 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U773 ( .A1(n729), .A2(n720), .ZN(n721) );
  NAND2_X1 U774 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U775 ( .A(KEYINPUT52), .B(n723), .Z(n724) );
  NOR2_X1 U776 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U777 ( .A1(n726), .A2(G952), .ZN(n727) );
  NAND2_X1 U778 ( .A1(n727), .A2(n464), .ZN(n733) );
  INV_X1 U779 ( .A(n728), .ZN(n731) );
  INV_X1 U780 ( .A(n729), .ZN(n730) );
  NOR2_X1 U781 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U782 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U783 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U784 ( .A(KEYINPUT53), .B(n736), .Z(G75) );
  XNOR2_X1 U785 ( .A(G101), .B(n737), .ZN(G3) );
  NAND2_X1 U786 ( .A1(n739), .A2(n747), .ZN(n738) );
  XNOR2_X1 U787 ( .A(n738), .B(G104), .ZN(G6) );
  XOR2_X1 U788 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n741) );
  NAND2_X1 U789 ( .A1(n739), .A2(n749), .ZN(n740) );
  XNOR2_X1 U790 ( .A(n741), .B(n740), .ZN(n742) );
  XNOR2_X1 U791 ( .A(G107), .B(n742), .ZN(G9) );
  XOR2_X1 U792 ( .A(G128), .B(KEYINPUT29), .Z(n744) );
  NAND2_X1 U793 ( .A1(n745), .A2(n749), .ZN(n743) );
  XNOR2_X1 U794 ( .A(n744), .B(n743), .ZN(G30) );
  NAND2_X1 U795 ( .A1(n745), .A2(n747), .ZN(n746) );
  XNOR2_X1 U796 ( .A(n746), .B(G146), .ZN(G48) );
  NAND2_X1 U797 ( .A1(n750), .A2(n747), .ZN(n748) );
  XNOR2_X1 U798 ( .A(n748), .B(G113), .ZN(G15) );
  NAND2_X1 U799 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U800 ( .A(n751), .B(G116), .ZN(G18) );
  XOR2_X1 U801 ( .A(n752), .B(KEYINPUT118), .Z(n753) );
  XNOR2_X1 U802 ( .A(n753), .B(KEYINPUT37), .ZN(n754) );
  XNOR2_X1 U803 ( .A(G125), .B(n754), .ZN(G27) );
  NOR2_X1 U804 ( .A1(n756), .A2(n755), .ZN(n766) );
  BUF_X1 U805 ( .A(n757), .Z(n758) );
  NAND2_X1 U806 ( .A1(n758), .A2(n464), .ZN(n764) );
  XOR2_X1 U807 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n760) );
  NAND2_X1 U808 ( .A1(G224), .A2(G953), .ZN(n759) );
  XNOR2_X1 U809 ( .A(n760), .B(n759), .ZN(n761) );
  NAND2_X1 U810 ( .A1(G898), .A2(n761), .ZN(n762) );
  XNOR2_X1 U811 ( .A(n762), .B(KEYINPUT126), .ZN(n763) );
  NAND2_X1 U812 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U813 ( .A(n766), .B(n765), .ZN(G69) );
  XOR2_X1 U814 ( .A(n769), .B(n768), .Z(n772) );
  XNOR2_X1 U815 ( .A(n770), .B(n772), .ZN(n771) );
  NAND2_X1 U816 ( .A1(n771), .A2(n464), .ZN(n776) );
  XOR2_X1 U817 ( .A(n772), .B(G227), .Z(n773) );
  NAND2_X1 U818 ( .A1(n773), .A2(G900), .ZN(n774) );
  NAND2_X1 U819 ( .A1(n774), .A2(G953), .ZN(n775) );
  NAND2_X1 U820 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U821 ( .A(KEYINPUT127), .B(n777), .Z(G72) );
  XOR2_X1 U822 ( .A(G140), .B(n778), .Z(n779) );
  XNOR2_X1 U823 ( .A(KEYINPUT119), .B(n779), .ZN(G42) );
  XNOR2_X1 U824 ( .A(G143), .B(KEYINPUT117), .ZN(n781) );
  XNOR2_X1 U825 ( .A(n781), .B(n780), .ZN(G45) );
endmodule

