

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591;

  BUF_X1 U323 ( .A(n567), .Z(n563) );
  NOR2_X1 U324 ( .A1(n530), .A2(n480), .ZN(n410) );
  XNOR2_X1 U325 ( .A(n386), .B(KEYINPUT45), .ZN(n387) );
  XNOR2_X1 U326 ( .A(n410), .B(KEYINPUT54), .ZN(n412) );
  XNOR2_X1 U327 ( .A(n388), .B(n387), .ZN(n390) );
  XNOR2_X1 U328 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U329 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U330 ( .A(n360), .B(n359), .ZN(n361) );
  NOR2_X1 U331 ( .A1(n482), .A2(n456), .ZN(n567) );
  XNOR2_X1 U332 ( .A(n362), .B(n361), .ZN(n580) );
  XNOR2_X1 U333 ( .A(n382), .B(n403), .ZN(n544) );
  XNOR2_X1 U334 ( .A(n342), .B(n341), .ZN(n562) );
  XNOR2_X1 U335 ( .A(n459), .B(G190GAT), .ZN(n460) );
  XNOR2_X1 U336 ( .A(n461), .B(n460), .ZN(G1351GAT) );
  XNOR2_X1 U337 ( .A(G127GAT), .B(G134GAT), .ZN(n291) );
  XNOR2_X1 U338 ( .A(n291), .B(KEYINPUT0), .ZN(n292) );
  XOR2_X1 U339 ( .A(n292), .B(KEYINPUT80), .Z(n294) );
  XNOR2_X1 U340 ( .A(G113GAT), .B(G120GAT), .ZN(n293) );
  XNOR2_X1 U341 ( .A(n294), .B(n293), .ZN(n432) );
  XOR2_X1 U342 ( .A(KEYINPUT20), .B(G71GAT), .Z(n296) );
  XNOR2_X1 U343 ( .A(G15GAT), .B(G176GAT), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n432), .B(n297), .ZN(n309) );
  XOR2_X1 U346 ( .A(G190GAT), .B(KEYINPUT83), .Z(n301) );
  XOR2_X1 U347 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n299) );
  XNOR2_X1 U348 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n298) );
  XNOR2_X1 U349 ( .A(n299), .B(n298), .ZN(n407) );
  XNOR2_X1 U350 ( .A(G43GAT), .B(n407), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U352 ( .A(n302), .B(G99GAT), .Z(n307) );
  XOR2_X1 U353 ( .A(KEYINPUT82), .B(G183GAT), .Z(n304) );
  NAND2_X1 U354 ( .A1(G227GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U355 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U356 ( .A(KEYINPUT81), .B(n305), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U358 ( .A(n309), .B(n308), .ZN(n482) );
  XOR2_X1 U359 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n311) );
  XNOR2_X1 U360 ( .A(G127GAT), .B(G211GAT), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U362 ( .A(G8GAT), .B(G183GAT), .Z(n400) );
  XOR2_X1 U363 ( .A(n312), .B(n400), .Z(n315) );
  XOR2_X1 U364 ( .A(G15GAT), .B(G1GAT), .Z(n329) );
  XNOR2_X1 U365 ( .A(G22GAT), .B(G155GAT), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n313), .B(G78GAT), .ZN(n440) );
  XNOR2_X1 U367 ( .A(n329), .B(n440), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U369 ( .A(KEYINPUT14), .B(KEYINPUT78), .Z(n317) );
  NAND2_X1 U370 ( .A1(G231GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U372 ( .A(n319), .B(n318), .Z(n324) );
  XOR2_X1 U373 ( .A(G57GAT), .B(KEYINPUT13), .Z(n321) );
  XNOR2_X1 U374 ( .A(G71GAT), .B(G64GAT), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U376 ( .A(KEYINPUT70), .B(n322), .Z(n359) );
  XNOR2_X1 U377 ( .A(n359), .B(KEYINPUT79), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n490) );
  XOR2_X1 U379 ( .A(KEYINPUT107), .B(n490), .Z(n540) );
  XOR2_X1 U380 ( .A(G197GAT), .B(G22GAT), .Z(n326) );
  XNOR2_X1 U381 ( .A(G169GAT), .B(G141GAT), .ZN(n325) );
  XNOR2_X1 U382 ( .A(n326), .B(n325), .ZN(n342) );
  XOR2_X1 U383 ( .A(G29GAT), .B(G43GAT), .Z(n328) );
  XNOR2_X1 U384 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n380) );
  XOR2_X1 U386 ( .A(n329), .B(n380), .Z(n331) );
  XNOR2_X1 U387 ( .A(G36GAT), .B(G50GAT), .ZN(n330) );
  XNOR2_X1 U388 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U389 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n333) );
  NAND2_X1 U390 ( .A1(G229GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U392 ( .A(n335), .B(n334), .Z(n340) );
  XOR2_X1 U393 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n337) );
  XNOR2_X1 U394 ( .A(G113GAT), .B(G8GAT), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n338), .B(KEYINPUT68), .ZN(n339) );
  XNOR2_X1 U397 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U398 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n344) );
  XNOR2_X1 U399 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n344), .B(n343), .ZN(n351) );
  XOR2_X1 U401 ( .A(G176GAT), .B(G204GAT), .Z(n399) );
  XOR2_X1 U402 ( .A(KEYINPUT75), .B(KEYINPUT33), .Z(n346) );
  XNOR2_X1 U403 ( .A(G120GAT), .B(G78GAT), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U405 ( .A(n399), .B(n347), .ZN(n349) );
  AND2_X1 U406 ( .A1(G230GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n351), .B(n350), .ZN(n362) );
  XNOR2_X1 U409 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n352) );
  XNOR2_X1 U410 ( .A(n352), .B(G148GAT), .ZN(n452) );
  XNOR2_X1 U411 ( .A(G99GAT), .B(G92GAT), .ZN(n358) );
  INV_X1 U412 ( .A(KEYINPUT74), .ZN(n353) );
  NAND2_X1 U413 ( .A1(G85GAT), .A2(n353), .ZN(n356) );
  INV_X1 U414 ( .A(G85GAT), .ZN(n354) );
  NAND2_X1 U415 ( .A1(n354), .A2(KEYINPUT74), .ZN(n355) );
  NAND2_X1 U416 ( .A1(n356), .A2(n355), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n358), .B(n357), .ZN(n367) );
  XOR2_X1 U418 ( .A(n452), .B(n367), .Z(n360) );
  XNOR2_X1 U419 ( .A(KEYINPUT41), .B(n580), .ZN(n566) );
  AND2_X1 U420 ( .A1(n562), .A2(n566), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n363), .B(KEYINPUT46), .ZN(n364) );
  NOR2_X1 U422 ( .A1(n540), .A2(n364), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n365), .B(KEYINPUT108), .ZN(n383) );
  INV_X1 U424 ( .A(KEYINPUT11), .ZN(n366) );
  XNOR2_X1 U425 ( .A(n367), .B(n366), .ZN(n369) );
  XOR2_X1 U426 ( .A(G50GAT), .B(G162GAT), .Z(n446) );
  XNOR2_X1 U427 ( .A(n446), .B(KEYINPUT9), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n378) );
  XOR2_X1 U429 ( .A(KEYINPUT10), .B(KEYINPUT77), .Z(n371) );
  XNOR2_X1 U430 ( .A(KEYINPUT64), .B(KEYINPUT76), .ZN(n370) );
  XNOR2_X1 U431 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U432 ( .A(G134GAT), .B(n372), .ZN(n376) );
  XOR2_X1 U433 ( .A(G106GAT), .B(KEYINPUT65), .Z(n374) );
  NAND2_X1 U434 ( .A1(G232GAT), .A2(G233GAT), .ZN(n373) );
  XOR2_X1 U435 ( .A(n374), .B(n373), .Z(n375) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n382) );
  XNOR2_X1 U437 ( .A(G36GAT), .B(G190GAT), .ZN(n381) );
  XOR2_X1 U438 ( .A(n381), .B(G218GAT), .Z(n403) );
  INV_X1 U439 ( .A(n544), .ZN(n559) );
  NAND2_X1 U440 ( .A1(n383), .A2(n559), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n384), .B(KEYINPUT47), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n385), .B(KEYINPUT109), .ZN(n393) );
  XNOR2_X1 U443 ( .A(KEYINPUT36), .B(n544), .ZN(n588) );
  NAND2_X1 U444 ( .A1(n588), .A2(n490), .ZN(n388) );
  INV_X1 U445 ( .A(KEYINPUT66), .ZN(n386) );
  INV_X1 U446 ( .A(n562), .ZN(n575) );
  AND2_X1 U447 ( .A1(n580), .A2(n575), .ZN(n389) );
  AND2_X1 U448 ( .A1(n390), .A2(n389), .ZN(n391) );
  XOR2_X1 U449 ( .A(KEYINPUT110), .B(n391), .Z(n392) );
  NAND2_X1 U450 ( .A1(n393), .A2(n392), .ZN(n395) );
  XNOR2_X1 U451 ( .A(KEYINPUT111), .B(KEYINPUT48), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n395), .B(n394), .ZN(n530) );
  XOR2_X1 U453 ( .A(G64GAT), .B(KEYINPUT93), .Z(n397) );
  NAND2_X1 U454 ( .A1(G226GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U456 ( .A(n398), .B(G92GAT), .Z(n402) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n402), .B(n401), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n404), .B(n403), .ZN(n409) );
  XOR2_X1 U460 ( .A(G211GAT), .B(KEYINPUT85), .Z(n406) );
  XNOR2_X1 U461 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n439) );
  XNOR2_X1 U463 ( .A(n407), .B(n439), .ZN(n408) );
  XNOR2_X1 U464 ( .A(n409), .B(n408), .ZN(n480) );
  INV_X1 U465 ( .A(n412), .ZN(n411) );
  NAND2_X1 U466 ( .A1(n411), .A2(KEYINPUT119), .ZN(n415) );
  INV_X1 U467 ( .A(KEYINPUT119), .ZN(n413) );
  NAND2_X1 U468 ( .A1(n413), .A2(n412), .ZN(n414) );
  NAND2_X1 U469 ( .A1(n415), .A2(n414), .ZN(n435) );
  XOR2_X1 U470 ( .A(KEYINPUT6), .B(G57GAT), .Z(n417) );
  XNOR2_X1 U471 ( .A(G1GAT), .B(G155GAT), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U473 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n419) );
  XNOR2_X1 U474 ( .A(KEYINPUT89), .B(KEYINPUT1), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U476 ( .A(n421), .B(n420), .Z(n426) );
  XOR2_X1 U477 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n423) );
  NAND2_X1 U478 ( .A1(G225GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U480 ( .A(KEYINPUT92), .B(n424), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n431) );
  XOR2_X1 U482 ( .A(G85GAT), .B(G162GAT), .Z(n429) );
  XNOR2_X1 U483 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n427), .B(KEYINPUT2), .ZN(n451) );
  XNOR2_X1 U485 ( .A(G29GAT), .B(n451), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U487 ( .A(n431), .B(n430), .Z(n434) );
  XNOR2_X1 U488 ( .A(n432), .B(G148GAT), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n469) );
  NAND2_X1 U490 ( .A1(n435), .A2(n469), .ZN(n572) );
  XOR2_X1 U491 ( .A(KEYINPUT22), .B(G204GAT), .Z(n437) );
  NAND2_X1 U492 ( .A1(G228GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U494 ( .A(n438), .B(KEYINPUT88), .Z(n442) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n450) );
  XOR2_X1 U497 ( .A(KEYINPUT86), .B(KEYINPUT24), .Z(n444) );
  XNOR2_X1 U498 ( .A(KEYINPUT84), .B(KEYINPUT87), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U500 ( .A(n445), .B(KEYINPUT23), .Z(n448) );
  XNOR2_X1 U501 ( .A(n446), .B(G218GAT), .ZN(n447) );
  XNOR2_X1 U502 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U503 ( .A(n450), .B(n449), .Z(n454) );
  XNOR2_X1 U504 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U505 ( .A(n454), .B(n453), .ZN(n471) );
  NOR2_X1 U506 ( .A1(n572), .A2(n471), .ZN(n455) );
  XNOR2_X1 U507 ( .A(n455), .B(KEYINPUT55), .ZN(n456) );
  NAND2_X1 U508 ( .A1(n563), .A2(n540), .ZN(n458) );
  XNOR2_X1 U509 ( .A(G183GAT), .B(KEYINPUT122), .ZN(n457) );
  XNOR2_X1 U510 ( .A(n458), .B(n457), .ZN(G1350GAT) );
  NAND2_X1 U511 ( .A1(n563), .A2(n544), .ZN(n461) );
  XOR2_X1 U512 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n459) );
  INV_X1 U513 ( .A(n469), .ZN(n519) );
  NAND2_X1 U514 ( .A1(n562), .A2(n580), .ZN(n493) );
  INV_X1 U515 ( .A(n490), .ZN(n585) );
  NOR2_X1 U516 ( .A1(n544), .A2(n585), .ZN(n462) );
  XNOR2_X1 U517 ( .A(n462), .B(KEYINPUT16), .ZN(n477) );
  NOR2_X1 U518 ( .A1(n482), .A2(n480), .ZN(n463) );
  NOR2_X1 U519 ( .A1(n471), .A2(n463), .ZN(n464) );
  XNOR2_X1 U520 ( .A(n464), .B(KEYINPUT25), .ZN(n467) );
  XOR2_X1 U521 ( .A(n480), .B(KEYINPUT27), .Z(n472) );
  NAND2_X1 U522 ( .A1(n471), .A2(n482), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n465), .B(KEYINPUT26), .ZN(n573) );
  INV_X1 U524 ( .A(n573), .ZN(n549) );
  NAND2_X1 U525 ( .A1(n472), .A2(n549), .ZN(n466) );
  NAND2_X1 U526 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U527 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n470), .B(KEYINPUT94), .ZN(n475) );
  XNOR2_X1 U529 ( .A(n471), .B(KEYINPUT28), .ZN(n534) );
  NAND2_X1 U530 ( .A1(n472), .A2(n519), .ZN(n529) );
  NOR2_X1 U531 ( .A1(n534), .A2(n529), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n473), .A2(n482), .ZN(n474) );
  NAND2_X1 U533 ( .A1(n475), .A2(n474), .ZN(n476) );
  XOR2_X1 U534 ( .A(KEYINPUT95), .B(n476), .Z(n488) );
  NAND2_X1 U535 ( .A1(n477), .A2(n488), .ZN(n508) );
  NOR2_X1 U536 ( .A1(n493), .A2(n508), .ZN(n486) );
  NAND2_X1 U537 ( .A1(n519), .A2(n486), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n478), .B(KEYINPUT34), .ZN(n479) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(n479), .ZN(G1324GAT) );
  INV_X1 U540 ( .A(n480), .ZN(n522) );
  NAND2_X1 U541 ( .A1(n522), .A2(n486), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT96), .B(KEYINPUT35), .Z(n484) );
  INV_X1 U544 ( .A(n482), .ZN(n531) );
  NAND2_X1 U545 ( .A1(n486), .A2(n531), .ZN(n483) );
  XNOR2_X1 U546 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U547 ( .A(G15GAT), .B(n485), .ZN(G1326GAT) );
  NAND2_X1 U548 ( .A1(n534), .A2(n486), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n487), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U550 ( .A1(n588), .A2(n488), .ZN(n489) );
  NOR2_X1 U551 ( .A1(n490), .A2(n489), .ZN(n492) );
  XNOR2_X1 U552 ( .A(KEYINPUT37), .B(KEYINPUT98), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(n518) );
  NOR2_X1 U554 ( .A1(n493), .A2(n518), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n494), .B(KEYINPUT38), .ZN(n504) );
  NAND2_X1 U556 ( .A1(n504), .A2(n519), .ZN(n498) );
  XOR2_X1 U557 ( .A(KEYINPUT99), .B(KEYINPUT39), .Z(n496) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT97), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NAND2_X1 U561 ( .A1(n504), .A2(n522), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n499), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(KEYINPUT101), .ZN(n503) );
  XOR2_X1 U564 ( .A(KEYINPUT40), .B(KEYINPUT100), .Z(n501) );
  NAND2_X1 U565 ( .A1(n504), .A2(n531), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(G1330GAT) );
  NAND2_X1 U568 ( .A1(n504), .A2(n534), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(KEYINPUT102), .ZN(n506) );
  XNOR2_X1 U570 ( .A(G50GAT), .B(n506), .ZN(G1331GAT) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n510) );
  INV_X1 U572 ( .A(n566), .ZN(n552) );
  NOR2_X1 U573 ( .A1(n552), .A2(n562), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n507), .B(KEYINPUT103), .ZN(n517) );
  NOR2_X1 U575 ( .A1(n517), .A2(n508), .ZN(n514) );
  NAND2_X1 U576 ( .A1(n514), .A2(n519), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n510), .B(n509), .ZN(G1332GAT) );
  NAND2_X1 U578 ( .A1(n522), .A2(n514), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n511), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U580 ( .A1(n531), .A2(n514), .ZN(n512) );
  XNOR2_X1 U581 ( .A(n512), .B(KEYINPUT104), .ZN(n513) );
  XNOR2_X1 U582 ( .A(G71GAT), .B(n513), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U584 ( .A1(n514), .A2(n534), .ZN(n515) );
  XNOR2_X1 U585 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  XOR2_X1 U586 ( .A(G85GAT), .B(KEYINPUT105), .Z(n521) );
  NOR2_X1 U587 ( .A1(n518), .A2(n517), .ZN(n526) );
  NAND2_X1 U588 ( .A1(n526), .A2(n519), .ZN(n520) );
  XNOR2_X1 U589 ( .A(n521), .B(n520), .ZN(G1336GAT) );
  NAND2_X1 U590 ( .A1(n522), .A2(n526), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n523), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U592 ( .A1(n531), .A2(n526), .ZN(n524) );
  XNOR2_X1 U593 ( .A(n524), .B(KEYINPUT106), .ZN(n525) );
  XNOR2_X1 U594 ( .A(G99GAT), .B(n525), .ZN(G1338GAT) );
  NAND2_X1 U595 ( .A1(n534), .A2(n526), .ZN(n527) );
  XNOR2_X1 U596 ( .A(n527), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NOR2_X1 U598 ( .A1(n530), .A2(n529), .ZN(n550) );
  NAND2_X1 U599 ( .A1(n550), .A2(n531), .ZN(n532) );
  XNOR2_X1 U600 ( .A(KEYINPUT112), .B(n532), .ZN(n533) );
  NOR2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n562), .A2(n545), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n535), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n537) );
  NAND2_X1 U605 ( .A1(n545), .A2(n566), .ZN(n536) );
  XNOR2_X1 U606 ( .A(n537), .B(n536), .ZN(n539) );
  XOR2_X1 U607 ( .A(G120GAT), .B(KEYINPUT113), .Z(n538) );
  XNOR2_X1 U608 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n542) );
  NAND2_X1 U610 ( .A1(n545), .A2(n540), .ZN(n541) );
  XNOR2_X1 U611 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U614 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(G134GAT), .B(n548), .ZN(G1343GAT) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n558) );
  NOR2_X1 U618 ( .A1(n575), .A2(n558), .ZN(n551) );
  XOR2_X1 U619 ( .A(G141GAT), .B(n551), .Z(G1344GAT) );
  NOR2_X1 U620 ( .A1(n558), .A2(n552), .ZN(n556) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n553) );
  XNOR2_X1 U623 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  NOR2_X1 U625 ( .A1(n585), .A2(n558), .ZN(n557) );
  XOR2_X1 U626 ( .A(G155GAT), .B(n557), .Z(G1346GAT) );
  NOR2_X1 U627 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U628 ( .A(KEYINPUT118), .B(n560), .Z(n561) );
  XNOR2_X1 U629 ( .A(G162GAT), .B(n561), .ZN(G1347GAT) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1348GAT) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n569) );
  XOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT57), .Z(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n571) );
  XOR2_X1 U636 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(KEYINPUT124), .B(n574), .ZN(n589) );
  INV_X1 U640 ( .A(n589), .ZN(n586) );
  NOR2_X1 U641 ( .A1(n586), .A2(n575), .ZN(n579) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n577) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  NOR2_X1 U646 ( .A1(n580), .A2(n586), .ZN(n584) );
  XOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n582) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n581) );
  XNOR2_X1 U649 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U652 ( .A(G211GAT), .B(n587), .Z(G1354GAT) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(n590), .B(KEYINPUT62), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

