//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT64), .A2(G128), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT64), .A2(G128), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n195), .B1(G143), .B2(new_n187), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n191), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT11), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G137), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT11), .A3(G134), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(G137), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n205), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n204), .A2(G137), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n206), .A2(G134), .ZN(new_n212));
  OAI21_X1  g026(.A(G131), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n210), .A2(new_n213), .A3(KEYINPUT67), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT67), .B1(new_n210), .B2(new_n213), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n202), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  OR2_X1    g031(.A1(KEYINPUT0), .A2(G128), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n191), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n198), .A2(KEYINPUT0), .A3(G128), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n205), .A2(new_n207), .A3(new_n209), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G131), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(new_n210), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n221), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n222), .B1(new_n221), .B2(new_n225), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n216), .B(KEYINPUT30), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n199), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT64), .A2(G128), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n198), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n200), .A2(new_n188), .A3(new_n190), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n210), .B(new_n213), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n224), .A2(new_n210), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n219), .A2(new_n220), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT30), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n229), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n228), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT66), .B1(new_n238), .B2(new_n239), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n221), .A2(new_n225), .A3(new_n222), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n246), .A2(new_n229), .A3(KEYINPUT30), .A4(new_n216), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G119), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT65), .B1(new_n249), .B2(G116), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT65), .ZN(new_n251));
  INV_X1    g065(.A(G116), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n252), .A3(G119), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n250), .A2(new_n253), .B1(G116), .B2(new_n249), .ZN(new_n254));
  XOR2_X1   g068(.A(KEYINPUT2), .B(G113), .Z(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n248), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n256), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n216), .B(new_n258), .C1(new_n226), .C2(new_n227), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT69), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n246), .A2(new_n261), .A3(new_n258), .A4(new_n216), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(G237), .A2(G953), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G210), .ZN(new_n265));
  XOR2_X1   g079(.A(new_n265), .B(KEYINPUT27), .Z(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT26), .B(G101), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n257), .A2(new_n263), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT31), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n240), .A2(new_n256), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n272), .B1(new_n263), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n256), .B1(new_n225), .B2(new_n221), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT28), .B1(new_n275), .B2(new_n216), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n268), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT31), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n257), .A2(new_n278), .A3(new_n263), .A4(new_n269), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n271), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(G472), .A2(G902), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT70), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT32), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n280), .A2(new_n285), .A3(new_n281), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n283), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n269), .B1(new_n274), .B2(new_n276), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n257), .A2(new_n263), .A3(new_n268), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT29), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n246), .A2(new_n216), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n256), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n263), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT28), .ZN(new_n294));
  INV_X1    g108(.A(new_n276), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n269), .A2(KEYINPUT29), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G472), .B1(new_n290), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n280), .A2(KEYINPUT32), .A3(new_n281), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n287), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G221), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT9), .B(G234), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n304), .B1(new_n306), .B2(new_n298), .ZN(new_n307));
  XNOR2_X1  g121(.A(G110), .B(G140), .ZN(new_n308));
  INV_X1    g122(.A(G953), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n309), .A2(G227), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n308), .B(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G104), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT3), .B1(new_n313), .B2(G107), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n315));
  INV_X1    g129(.A(G107), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(G104), .ZN(new_n317));
  INV_X1    g131(.A(G101), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n313), .A2(G107), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n314), .A2(new_n317), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n313), .A2(G107), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n316), .A2(G104), .ZN(new_n322));
  OAI21_X1  g136(.A(G101), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n234), .A2(G128), .B1(new_n188), .B2(new_n190), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n320), .B(new_n323), .C1(new_n324), .C2(new_n236), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n320), .A2(new_n323), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n325), .B1(new_n202), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n225), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT12), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(KEYINPUT12), .A3(new_n225), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n314), .A2(new_n317), .A3(new_n319), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(G101), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT73), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT73), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n333), .A2(new_n337), .A3(new_n334), .A4(G101), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n333), .A2(G101), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(KEYINPUT4), .A3(new_n320), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n221), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT10), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n343), .B1(new_n197), .B2(new_n201), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n326), .A2(new_n344), .B1(new_n325), .B2(new_n343), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n238), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n312), .B1(new_n332), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n312), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n238), .B1(new_n342), .B2(new_n345), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(G469), .B1(new_n351), .B2(G902), .ZN(new_n352));
  INV_X1    g166(.A(G469), .ZN(new_n353));
  INV_X1    g167(.A(new_n349), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n312), .B1(new_n354), .B2(new_n346), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n327), .A2(KEYINPUT12), .A3(new_n225), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT12), .B1(new_n327), .B2(new_n225), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n348), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n353), .B(new_n298), .C1(new_n355), .C2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n307), .B1(new_n352), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G217), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(G234), .B2(new_n298), .ZN(new_n364));
  INV_X1    g178(.A(G140), .ZN(new_n365));
  INV_X1    g179(.A(G125), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n365), .B1(new_n366), .B2(KEYINPUT71), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT71), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(G125), .A3(G140), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(KEYINPUT16), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n365), .A2(G125), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT16), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n370), .A2(new_n187), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT72), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n370), .A2(new_n373), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G146), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n370), .A2(KEYINPUT72), .A3(new_n187), .A4(new_n373), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT23), .B1(new_n199), .B2(G119), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n199), .A2(G119), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n383), .B1(new_n194), .B2(G119), .ZN(new_n386));
  XOR2_X1   g200(.A(KEYINPUT24), .B(G110), .Z(new_n387));
  AOI22_X1  g201(.A1(new_n385), .A2(G110), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n380), .A2(new_n388), .ZN(new_n389));
  OAI22_X1  g203(.A1(new_n385), .A2(G110), .B1(new_n386), .B2(new_n387), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n366), .A2(G140), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n371), .A2(new_n391), .A3(new_n187), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n378), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT22), .B(G137), .ZN(new_n395));
  INV_X1    g209(.A(G234), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n304), .A2(new_n396), .A3(G953), .ZN(new_n397));
  XOR2_X1   g211(.A(new_n395), .B(new_n397), .Z(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n394), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n389), .A2(new_n393), .A3(new_n398), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n402), .A2(KEYINPUT25), .A3(new_n298), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT25), .B1(new_n402), .B2(new_n298), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n364), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n364), .A2(G902), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n362), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G214), .B1(G237), .B2(G902), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT74), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n339), .A2(new_n256), .A3(new_n341), .ZN(new_n413));
  XNOR2_X1  g227(.A(G110), .B(G122), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT5), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(new_n249), .A3(G116), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G113), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n417), .B1(new_n254), .B2(KEYINPUT5), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n254), .A2(new_n255), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(new_n420), .A3(new_n326), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n413), .A2(new_n414), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n239), .A2(G125), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n197), .A2(new_n366), .A3(new_n201), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G224), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT7), .B1(new_n427), .B2(G953), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n428), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n424), .A2(new_n425), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  XOR2_X1   g246(.A(new_n414), .B(KEYINPUT8), .Z(new_n433));
  NAND2_X1  g247(.A1(new_n320), .A2(new_n323), .ZN(new_n434));
  INV_X1    g248(.A(new_n420), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n434), .B1(new_n435), .B2(new_n418), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n433), .B1(new_n421), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n423), .B1(new_n438), .B2(KEYINPUT75), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT75), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n440), .B1(new_n432), .B2(new_n437), .ZN(new_n441));
  AOI21_X1  g255(.A(G902), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(G210), .B1(G237), .B2(G902), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n413), .A2(new_n421), .ZN(new_n444));
  INV_X1    g258(.A(new_n414), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT6), .A3(new_n422), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT6), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(new_n448), .A3(new_n445), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n427), .A2(G953), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n426), .B(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n442), .A2(new_n443), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n443), .B(KEYINPUT76), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n456), .B1(new_n442), .B2(new_n452), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n412), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT87), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n231), .A2(G143), .A3(new_n232), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n189), .A2(G128), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n204), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT83), .B1(new_n252), .B2(G122), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT83), .ZN(new_n465));
  INV_X1    g279(.A(G122), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(G116), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n252), .A2(G122), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n468), .B(new_n469), .C1(KEYINPUT14), .C2(new_n316), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n460), .A2(G134), .A3(new_n461), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n463), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n464), .A2(new_n467), .B1(new_n252), .B2(G122), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT14), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(new_n464), .B2(new_n467), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n473), .A2(new_n475), .A3(new_n316), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT13), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n460), .A2(new_n479), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n480), .A2(G134), .B1(new_n460), .B2(new_n461), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n460), .A2(KEYINPUT13), .A3(G134), .A4(new_n461), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n473), .A2(new_n316), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n468), .A2(new_n316), .A3(new_n469), .ZN(new_n485));
  OAI22_X1  g299(.A1(new_n481), .A2(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT84), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT13), .B1(new_n194), .B2(G143), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n462), .B1(new_n489), .B2(new_n204), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n482), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n473), .B(new_n316), .ZN(new_n492));
  AOI21_X1  g306(.A(KEYINPUT84), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n478), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n305), .A2(new_n363), .A3(G953), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n486), .A2(new_n487), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n491), .A2(KEYINPUT84), .A3(new_n492), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(new_n478), .A3(new_n495), .ZN(new_n501));
  AOI21_X1  g315(.A(G902), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT86), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n495), .B1(new_n500), .B2(new_n478), .ZN(new_n505));
  AOI211_X1 g319(.A(new_n477), .B(new_n496), .C1(new_n498), .C2(new_n499), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n298), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT86), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(G478), .B1(KEYINPUT85), .B2(KEYINPUT15), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(KEYINPUT85), .B2(KEYINPUT15), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n512), .B1(new_n502), .B2(new_n503), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G237), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(new_n309), .A3(G214), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n189), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n264), .A2(G143), .A3(G214), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(KEYINPUT18), .A2(G131), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT78), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT78), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n519), .A2(new_n525), .A3(new_n520), .A4(new_n522), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT77), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n368), .A2(G125), .A3(G140), .ZN(new_n529));
  AOI21_X1  g343(.A(G140), .B1(new_n368), .B2(G125), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n367), .A2(KEYINPUT77), .A3(new_n369), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(G146), .A3(new_n532), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n533), .A2(new_n392), .B1(new_n521), .B2(new_n523), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(KEYINPUT19), .A3(new_n532), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT19), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n371), .A2(new_n391), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n187), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n518), .A2(new_n189), .ZN(new_n539));
  AOI21_X1  g353(.A(G143), .B1(new_n264), .B2(G214), .ZN(new_n540));
  OAI21_X1  g354(.A(G131), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n519), .A2(new_n208), .A3(new_n520), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n541), .A2(new_n542), .B1(new_n377), .B2(G146), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n527), .A2(new_n534), .B1(new_n538), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(G113), .B(G122), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(new_n313), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT79), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n521), .A2(new_n523), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n533), .A2(new_n392), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n527), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n538), .A2(new_n543), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT79), .ZN(new_n553));
  INV_X1    g367(.A(new_n546), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n539), .A2(new_n540), .A3(G131), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n208), .B1(new_n519), .B2(new_n520), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n541), .A2(KEYINPUT17), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n556), .A2(new_n562), .B1(new_n527), .B2(new_n534), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n546), .B(KEYINPUT80), .Z(new_n564));
  AOI22_X1  g378(.A1(new_n547), .A2(new_n555), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(G475), .A2(G902), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT81), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT20), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n563), .A2(new_n564), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n553), .B1(new_n552), .B2(new_n554), .ZN(new_n570));
  AOI211_X1 g384(.A(KEYINPUT79), .B(new_n546), .C1(new_n550), .C2(new_n551), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT20), .ZN(new_n573));
  INV_X1    g387(.A(new_n567), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT82), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n554), .B1(new_n563), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT17), .B1(new_n541), .B2(new_n542), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n559), .A2(new_n557), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n550), .B(new_n576), .C1(new_n580), .C2(new_n380), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n569), .B1(new_n577), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n298), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n568), .A2(new_n575), .B1(new_n584), .B2(G475), .ZN(new_n585));
  INV_X1    g399(.A(G952), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(G953), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n587), .B1(new_n396), .B2(new_n517), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AOI211_X1 g403(.A(new_n298), .B(new_n309), .C1(G234), .C2(G237), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT21), .B(G898), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n585), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n459), .B1(new_n516), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n514), .B1(new_n509), .B2(new_n512), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n596), .A2(KEYINPUT87), .A3(new_n593), .A4(new_n585), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n458), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n303), .A2(new_n409), .A3(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT88), .B(G101), .Z(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G3));
  NAND2_X1  g415(.A1(new_n280), .A2(new_n298), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G472), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n283), .A2(new_n603), .A3(new_n286), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n604), .A2(new_n408), .A3(new_n362), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT89), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n453), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n442), .A2(new_n452), .ZN(new_n608));
  INV_X1    g422(.A(new_n443), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n442), .A2(KEYINPUT89), .A3(new_n443), .A4(new_n452), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n593), .A3(new_n410), .ZN(new_n613));
  INV_X1    g427(.A(G478), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n497), .A2(new_n501), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT90), .ZN(new_n617));
  AOI21_X1  g431(.A(KEYINPUT33), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  AOI211_X1 g433(.A(KEYINPUT90), .B(new_n619), .C1(new_n497), .C2(new_n501), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n615), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n502), .A2(G478), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n568), .A2(new_n575), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n550), .B1(new_n580), .B2(new_n380), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n546), .B1(new_n625), .B2(KEYINPUT82), .ZN(new_n626));
  AOI22_X1  g440(.A1(new_n626), .A2(new_n581), .B1(new_n563), .B2(new_n564), .ZN(new_n627));
  OAI21_X1  g441(.A(G475), .B1(new_n627), .B2(G902), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n621), .A2(new_n623), .B1(new_n624), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n613), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n605), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n632), .B(KEYINPUT91), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT92), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NOR3_X1   g450(.A1(new_n565), .A2(KEYINPUT20), .A3(new_n567), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(KEYINPUT93), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n638), .B(new_n628), .C1(new_n624), .C2(KEYINPUT93), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n639), .A2(new_n596), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n613), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n605), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  AND3_X1   g458(.A1(new_n280), .A2(new_n285), .A3(new_n281), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n285), .B1(new_n280), .B2(new_n281), .ZN(new_n646));
  INV_X1    g460(.A(G472), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n280), .B2(new_n298), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n399), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n394), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n406), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n405), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n598), .A2(new_n649), .A3(new_n361), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT37), .B(G110), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT94), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n654), .B(new_n656), .ZN(G12));
  INV_X1    g471(.A(G900), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n590), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n588), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n640), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n612), .A2(new_n410), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n361), .A2(new_n653), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n645), .A2(new_n646), .A3(KEYINPUT32), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n300), .A2(new_n301), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n662), .B(new_n665), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G128), .ZN(G30));
  OAI21_X1  g483(.A(new_n298), .B1(new_n293), .B2(new_n269), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n268), .B1(new_n257), .B2(new_n263), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n301), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n287), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n674), .A2(KEYINPUT96), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(KEYINPUT96), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT97), .B(KEYINPUT39), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n660), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n361), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n573), .B1(new_n572), .B2(new_n574), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n628), .B1(new_n637), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n516), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n410), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n684), .A2(new_n685), .A3(new_n653), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n454), .A2(new_n457), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n690));
  AND4_X1   g504(.A1(new_n681), .A2(new_n686), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n677), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G143), .ZN(G45));
  INV_X1    g507(.A(new_n615), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n617), .B1(new_n505), .B2(new_n506), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n619), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n617), .B(KEYINPUT33), .C1(new_n505), .C2(new_n506), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n683), .B(new_n660), .C1(new_n698), .C2(new_n622), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT98), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n621), .A2(new_n623), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT98), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n701), .A2(new_n702), .A3(new_n683), .A4(new_n660), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n704), .B(new_n665), .C1(new_n666), .C2(new_n667), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  INV_X1    g520(.A(new_n408), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n298), .B1(new_n355), .B2(new_n359), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(G469), .ZN(new_n709));
  INV_X1    g523(.A(new_n307), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n710), .A3(new_n360), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n303), .A2(new_n707), .A3(new_n631), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT99), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n713), .B(new_n715), .ZN(G15));
  AOI21_X1  g530(.A(new_n408), .B1(new_n287), .B2(new_n302), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n641), .A3(new_n712), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  NAND2_X1  g533(.A1(new_n595), .A2(new_n597), .ZN(new_n720));
  AND4_X1   g534(.A1(new_n410), .A2(new_n612), .A3(new_n653), .A4(new_n712), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n303), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT100), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n287), .A2(new_n302), .B1(new_n595), .B2(new_n597), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT100), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n725), .A3(new_n721), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  NOR3_X1   g542(.A1(new_n596), .A2(new_n711), .A3(new_n585), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n729), .A2(new_n593), .A3(new_n410), .A4(new_n612), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n276), .B1(new_n293), .B2(KEYINPUT28), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n271), .B(new_n279), .C1(new_n269), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n281), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n603), .A2(new_n707), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(KEYINPUT101), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT101), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n602), .A2(G472), .B1(new_n281), .B2(new_n733), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n737), .B1(new_n738), .B2(new_n707), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n731), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT102), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n735), .A2(KEYINPUT101), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n738), .A2(new_n737), .A3(new_n707), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(KEYINPUT102), .A3(new_n731), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g561(.A(KEYINPUT103), .B(G122), .Z(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G24));
  INV_X1    g563(.A(KEYINPUT104), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n702), .B1(new_n629), .B2(new_n660), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n696), .A2(new_n697), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n622), .B1(new_n752), .B2(new_n615), .ZN(new_n753));
  NOR4_X1   g567(.A1(new_n753), .A2(new_n585), .A3(KEYINPUT98), .A4(new_n661), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n750), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n700), .A2(KEYINPUT104), .A3(new_n703), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n721), .A3(new_n738), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G125), .ZN(G27));
  INV_X1    g572(.A(KEYINPUT42), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n454), .A2(new_n457), .A3(new_n685), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n760), .A2(new_n361), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n707), .B(new_n761), .C1(new_n666), .C2(new_n667), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n755), .A2(new_n756), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n301), .A2(KEYINPUT105), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n282), .A2(new_n284), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT105), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n280), .A2(new_n767), .A3(KEYINPUT32), .A4(new_n281), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n765), .A2(new_n766), .A3(new_n300), .A4(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n769), .A2(new_n707), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n700), .A2(KEYINPUT104), .A3(new_n703), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT104), .B1(new_n700), .B2(new_n703), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n761), .A2(KEYINPUT42), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n770), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n764), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G131), .ZN(G33));
  NAND4_X1  g591(.A1(new_n303), .A2(new_n707), .A3(new_n662), .A4(new_n761), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G134), .ZN(G36));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT43), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n701), .A2(new_n781), .A3(new_n585), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT43), .B1(new_n753), .B2(new_n683), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n783), .A3(new_n653), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n780), .B1(new_n649), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n782), .A2(new_n783), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(new_n604), .A3(KEYINPUT44), .A4(new_n653), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n347), .B2(new_n350), .ZN(new_n790));
  INV_X1    g604(.A(new_n346), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n311), .B1(new_n358), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n354), .A2(new_n346), .A3(new_n312), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(KEYINPUT45), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n790), .A2(new_n794), .A3(G469), .ZN(new_n795));
  NAND2_X1  g609(.A1(G469), .A2(G902), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT46), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n795), .A2(KEYINPUT46), .A3(new_n796), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n360), .A3(new_n800), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n710), .A2(new_n801), .A3(new_n679), .A4(new_n760), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n785), .A2(new_n788), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  INV_X1    g618(.A(KEYINPUT47), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n795), .A2(KEYINPUT46), .A3(new_n796), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT46), .B1(new_n795), .B2(new_n796), .ZN(new_n807));
  INV_X1    g621(.A(new_n360), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n805), .B1(new_n809), .B2(new_n307), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n801), .A2(KEYINPUT47), .A3(new_n710), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n645), .A2(new_n646), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n667), .B1(new_n813), .B2(new_n284), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n408), .A2(new_n700), .A3(new_n703), .A4(new_n760), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  NAND3_X1  g631(.A1(new_n707), .A2(new_n710), .A3(new_n412), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT106), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n709), .A2(new_n360), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n820), .A2(KEYINPUT49), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(KEYINPUT49), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n821), .A2(new_n585), .A3(new_n701), .A4(new_n822), .ZN(new_n823));
  OR4_X1    g637(.A1(new_n677), .A2(new_n689), .A3(new_n819), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n586), .A2(new_n309), .ZN(new_n825));
  INV_X1    g639(.A(new_n677), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n760), .A2(new_n712), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n827), .A2(new_n707), .A3(new_n589), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n826), .A2(new_n585), .A3(new_n753), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n786), .A2(new_n588), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n830), .A2(new_n827), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n653), .A3(new_n738), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n833), .A2(KEYINPUT111), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n745), .A2(new_n830), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n689), .A2(new_n410), .A3(new_n711), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT50), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n810), .B(new_n811), .C1(new_n710), .C2(new_n820), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n842), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n760), .A3(new_n835), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n833), .A2(KEYINPUT111), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n834), .A2(new_n840), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n835), .A2(new_n760), .A3(new_n841), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n829), .A2(new_n832), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n839), .B1(new_n849), .B2(new_n838), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n826), .A2(new_n629), .A3(new_n828), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n835), .A2(new_n410), .A3(new_n612), .A4(new_n712), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n851), .A2(new_n587), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n831), .A2(new_n770), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(KEYINPUT48), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT113), .Z(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(KEYINPUT48), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT114), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n853), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n847), .A2(new_n850), .A3(new_n859), .ZN(new_n860));
  XNOR2_X1  g674(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n742), .A2(new_n746), .B1(new_n723), .B2(new_n726), .ZN(new_n862));
  OR3_X1    g676(.A1(new_n596), .A2(KEYINPUT107), .A3(new_n683), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT107), .B1(new_n596), .B2(new_n683), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n864), .A3(new_n630), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n458), .A2(new_n592), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n865), .A2(new_n649), .A3(new_n409), .A4(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n713), .A2(new_n599), .A3(new_n654), .A4(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n718), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n738), .ZN(new_n871));
  OR3_X1    g685(.A1(new_n516), .A2(new_n639), .A3(new_n661), .ZN(new_n872));
  OAI22_X1  g686(.A1(new_n763), .A2(new_n871), .B1(new_n814), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n761), .A2(new_n653), .ZN(new_n874));
  INV_X1    g688(.A(new_n762), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n873), .A2(new_n874), .B1(new_n875), .B2(new_n662), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n862), .A2(new_n870), .A3(new_n776), .A4(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n303), .B(new_n665), .C1(new_n662), .C2(new_n704), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n663), .A2(new_n684), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n362), .A2(new_n653), .A3(new_n661), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n674), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n878), .A2(new_n757), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT52), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n861), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT102), .B1(new_n745), .B2(new_n731), .ZN(new_n887));
  AOI211_X1 g701(.A(new_n741), .B(new_n730), .C1(new_n743), .C2(new_n744), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n725), .A2(new_n303), .A3(new_n720), .A4(new_n721), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n725), .B1(new_n724), .B2(new_n721), .ZN(new_n890));
  OAI22_X1  g704(.A1(new_n887), .A2(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n458), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n720), .A2(new_n409), .A3(new_n892), .ZN(new_n893));
  AOI211_X1 g707(.A(new_n458), .B(new_n664), .C1(new_n595), .C2(new_n597), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n893), .A2(new_n303), .B1(new_n894), .B2(new_n649), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n895), .A2(new_n713), .A3(new_n718), .A4(new_n867), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n873), .A2(new_n874), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n776), .A2(new_n898), .A3(new_n778), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT108), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n882), .A2(new_n900), .A3(KEYINPUT52), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n882), .A2(new_n900), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT52), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n897), .A2(new_n899), .A3(new_n901), .A4(new_n904), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n884), .B(new_n885), .C1(new_n886), .C2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n861), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n877), .A2(new_n883), .ZN(new_n908));
  AOI22_X1  g722(.A1(new_n907), .A2(new_n908), .B1(new_n905), .B2(new_n886), .ZN(new_n909));
  OAI211_X1 g723(.A(KEYINPUT110), .B(new_n906), .C1(new_n909), .C2(new_n885), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT110), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n905), .A2(new_n886), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n877), .A2(new_n883), .A3(new_n861), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n911), .B(KEYINPUT54), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n860), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT115), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n825), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI211_X1 g731(.A(KEYINPUT115), .B(new_n860), .C1(new_n910), .C2(new_n914), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n824), .B1(new_n917), .B2(new_n918), .ZN(G75));
  INV_X1    g733(.A(new_n877), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n920), .A2(KEYINPUT53), .A3(new_n901), .A4(new_n904), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n884), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(G902), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT117), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n298), .B1(new_n921), .B2(new_n884), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT117), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n925), .A2(new_n455), .A3(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n447), .A2(new_n449), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(new_n451), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT55), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(KEYINPUT56), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT116), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n926), .A2(new_n934), .A3(G210), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT56), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n934), .B1(new_n926), .B2(G210), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n931), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n309), .A2(G952), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n933), .A2(new_n939), .A3(new_n941), .ZN(G51));
  XNOR2_X1  g756(.A(new_n922), .B(new_n885), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n796), .B(KEYINPUT57), .ZN(new_n944));
  OAI22_X1  g758(.A1(new_n943), .A2(new_n944), .B1(new_n355), .B2(new_n359), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n795), .B(KEYINPUT118), .Z(new_n946));
  NAND3_X1  g760(.A1(new_n925), .A2(new_n927), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n940), .B1(new_n945), .B2(new_n947), .ZN(G54));
  AND2_X1   g762(.A1(KEYINPUT58), .A2(G475), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n925), .A2(new_n927), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n565), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n925), .A2(new_n572), .A3(new_n927), .A4(new_n949), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n951), .A2(new_n941), .A3(new_n952), .ZN(G60));
  NAND2_X1  g767(.A1(G478), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT59), .Z(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n752), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n941), .B1(new_n943), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n752), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n910), .A2(new_n914), .A3(new_n956), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(G63));
  NAND2_X1  g775(.A1(G217), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT119), .Z(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT60), .Z(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n921), .B2(new_n884), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n651), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(KEYINPUT120), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT121), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n969), .A2(KEYINPUT61), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n941), .B(new_n970), .C1(new_n966), .C2(new_n402), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT120), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n966), .A2(new_n972), .A3(new_n651), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n968), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n922), .A2(new_n964), .ZN(new_n975));
  INV_X1    g789(.A(new_n402), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n940), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n977), .A2(new_n969), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n977), .A2(new_n967), .A3(new_n970), .ZN(new_n979));
  AOI22_X1  g793(.A1(new_n974), .A2(new_n978), .B1(KEYINPUT61), .B2(new_n979), .ZN(G66));
  INV_X1    g794(.A(new_n591), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n309), .B1(new_n981), .B2(G224), .ZN(new_n982));
  INV_X1    g796(.A(new_n897), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n982), .B1(new_n983), .B2(new_n309), .ZN(new_n984));
  INV_X1    g798(.A(G898), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n929), .B1(new_n985), .B2(G953), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n984), .B(new_n986), .ZN(G69));
  INV_X1    g801(.A(KEYINPUT124), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n535), .A2(new_n537), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n248), .B(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n801), .A2(new_n710), .A3(new_n679), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n992), .A2(new_n769), .A3(new_n707), .A4(new_n879), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n816), .A2(new_n778), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(new_n764), .B2(new_n775), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT122), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n757), .A2(new_n668), .A3(new_n705), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n996), .B1(new_n997), .B2(new_n803), .ZN(new_n998));
  AND4_X1   g812(.A1(new_n996), .A2(new_n803), .A3(new_n757), .A4(new_n878), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n995), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n309), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n309), .A2(G900), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(KEYINPUT123), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n785), .A2(new_n788), .A3(new_n802), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n757), .A2(new_n705), .A3(new_n668), .ZN(new_n1006));
  OAI21_X1  g820(.A(KEYINPUT122), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n803), .A2(new_n996), .A3(new_n757), .A4(new_n878), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(G953), .B1(new_n1009), .B2(new_n995), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT123), .ZN(new_n1011));
  NOR3_X1   g825(.A1(new_n1010), .A2(new_n1011), .A3(new_n1002), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n991), .B1(new_n1004), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n309), .B1(G227), .B2(G900), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n875), .A2(new_n679), .A3(new_n865), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1016), .A2(new_n803), .A3(new_n816), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n692), .A2(new_n997), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1017), .B1(new_n1018), .B2(KEYINPUT62), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT62), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n692), .A2(new_n1020), .A3(new_n997), .ZN(new_n1021));
  AOI21_X1  g835(.A(G953), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1015), .B1(new_n1022), .B2(new_n991), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n988), .B1(new_n1013), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1011), .B1(new_n1010), .B2(new_n1002), .ZN(new_n1026));
  AND3_X1   g840(.A1(new_n816), .A2(new_n778), .A3(new_n993), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1027), .A2(new_n776), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1028), .B1(new_n1008), .B2(new_n1007), .ZN(new_n1029));
  OAI211_X1 g843(.A(KEYINPUT123), .B(new_n1003), .C1(new_n1029), .C2(G953), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n990), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1031));
  NOR3_X1   g845(.A1(new_n1031), .A2(KEYINPUT124), .A3(new_n1023), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT125), .ZN(new_n1033));
  OAI211_X1 g847(.A(new_n1033), .B(new_n991), .C1(new_n1004), .C2(new_n1012), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1034), .A2(new_n1014), .ZN(new_n1035));
  OAI21_X1  g849(.A(KEYINPUT125), .B1(new_n1022), .B2(new_n991), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1037));
  OAI22_X1  g851(.A1(new_n1025), .A2(new_n1032), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT126), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g854(.A(new_n1034), .B(new_n1014), .C1(new_n1031), .C2(new_n1036), .ZN(new_n1041));
  OAI211_X1 g855(.A(new_n1041), .B(KEYINPUT126), .C1(new_n1025), .C2(new_n1032), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1040), .A2(new_n1042), .ZN(G72));
  NAND3_X1  g857(.A1(new_n1019), .A2(new_n897), .A3(new_n1021), .ZN(new_n1044));
  NAND2_X1  g858(.A1(G472), .A2(G902), .ZN(new_n1045));
  XOR2_X1   g859(.A(new_n1045), .B(KEYINPUT63), .Z(new_n1046));
  NAND2_X1  g860(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1047), .A2(new_n671), .ZN(new_n1048));
  XNOR2_X1  g862(.A(new_n1048), .B(KEYINPUT127), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n289), .A2(new_n1046), .ZN(new_n1050));
  NOR3_X1   g864(.A1(new_n909), .A2(new_n671), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g865(.A(new_n1046), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1052), .B1(new_n1029), .B2(new_n897), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n941), .B1(new_n1053), .B2(new_n289), .ZN(new_n1054));
  NOR3_X1   g868(.A1(new_n1049), .A2(new_n1051), .A3(new_n1054), .ZN(G57));
endmodule


