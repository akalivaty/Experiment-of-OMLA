//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1265, new_n1266, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  AND2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n202), .A2(new_n203), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n203), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G107), .ZN(new_n227));
  INV_X1    g0027(.A(G264), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n225), .B1(new_n206), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n212), .B(new_n219), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT65), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n201), .A2(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n203), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n244), .B(new_n249), .ZN(G351));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G1), .A3(G13), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G274), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n252), .A2(new_n255), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n256), .B1(G226), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT3), .B(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G222), .A2(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G223), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n252), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n264), .B(new_n265), .C1(G77), .C2(new_n260), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G200), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(G190), .B2(new_n267), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT68), .ZN(new_n271));
  AOI21_X1  g0071(.A(KEYINPUT10), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n273), .A2(new_n216), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n205), .A2(new_n217), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT66), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G58), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT8), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G150), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n280), .A2(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n275), .B1(new_n276), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n254), .A2(G13), .A3(G20), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n274), .B1(G1), .B2(new_n217), .ZN(new_n290));
  MUX2_X1   g0090(.A(new_n289), .B(new_n290), .S(G50), .Z(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT9), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n270), .ZN(new_n294));
  XOR2_X1   g0094(.A(new_n272), .B(new_n294), .Z(new_n295));
  INV_X1    g0095(.A(G179), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n267), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(new_n292), .C1(G169), .C2(new_n267), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  INV_X1    g0100(.A(G232), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G1698), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n260), .B(new_n302), .C1(G226), .C2(G1698), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G97), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n252), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n255), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(new_n252), .A3(G274), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(new_n221), .B2(new_n257), .ZN(new_n308));
  OR3_X1    g0108(.A1(new_n305), .A2(KEYINPUT13), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT13), .B1(new_n305), .B2(new_n308), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n300), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT14), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT70), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n311), .A2(KEYINPUT70), .A3(new_n312), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n309), .A2(new_n310), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n311), .A2(new_n312), .B1(new_n318), .B2(new_n296), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n285), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n283), .B2(new_n206), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n323), .A2(KEYINPUT11), .A3(new_n275), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT12), .ZN(new_n325));
  INV_X1    g0125(.A(new_n289), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n203), .ZN(new_n327));
  NOR3_X1   g0127(.A1(new_n289), .A2(KEYINPUT12), .A3(G68), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n290), .A2(new_n203), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT11), .B1(new_n323), .B2(new_n275), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n324), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n321), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n318), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n332), .B1(new_n335), .B2(G190), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n318), .A2(G200), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT69), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n260), .A2(G232), .A3(new_n262), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n227), .B2(new_n260), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT3), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G33), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n345), .A2(new_n221), .A3(new_n262), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n265), .B1(new_n341), .B2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n347), .B(new_n307), .C1(new_n226), .C2(new_n257), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n300), .ZN(new_n349));
  XOR2_X1   g0149(.A(KEYINPUT8), .B(G58), .Z(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT67), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n285), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT15), .B(G87), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n354), .A2(new_n282), .B1(G20), .B2(G77), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n274), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n326), .A2(new_n206), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n290), .B2(new_n206), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n349), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n348), .A2(G179), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n356), .A2(new_n358), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n348), .A2(G200), .ZN(new_n363));
  INV_X1    g0163(.A(G190), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n362), .B(new_n363), .C1(new_n364), .C2(new_n348), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NOR4_X1   g0166(.A1(new_n299), .A2(new_n334), .A3(new_n339), .A4(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n278), .B(KEYINPUT8), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n290), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n280), .A2(new_n289), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT74), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT72), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n202), .B2(new_n203), .ZN(new_n375));
  NAND3_X1  g0175(.A1(KEYINPUT72), .A2(G58), .A3(G68), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n375), .A2(new_n213), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G159), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n377), .A2(new_n217), .B1(new_n378), .B2(new_n286), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT71), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n343), .ZN(new_n381));
  NAND2_X1  g0181(.A1(KEYINPUT71), .A2(KEYINPUT3), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(G33), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n342), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n217), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT7), .ZN(new_n386));
  AOI21_X1  g0186(.A(G20), .B1(new_n383), .B2(new_n342), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n203), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n379), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n274), .B1(new_n390), .B2(KEYINPUT16), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT16), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT73), .ZN(new_n393));
  AND2_X1   g0193(.A1(KEYINPUT71), .A2(KEYINPUT3), .ZN(new_n394));
  NOR2_X1   g0194(.A1(KEYINPUT71), .A2(KEYINPUT3), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n393), .B(new_n281), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n388), .A2(G20), .ZN(new_n397));
  AOI21_X1  g0197(.A(G33), .B1(new_n381), .B2(new_n382), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n344), .A2(KEYINPUT73), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n396), .B(new_n397), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n388), .B1(new_n260), .B2(G20), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n203), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n392), .B1(new_n402), .B2(new_n379), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n373), .B1(new_n391), .B2(new_n403), .ZN(new_n404));
  MUX2_X1   g0204(.A(G223), .B(G226), .S(G1698), .Z(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(new_n383), .A3(new_n342), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G33), .A2(G87), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n252), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n307), .B1(new_n301), .B2(new_n257), .ZN(new_n409));
  NOR4_X1   g0209(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT75), .A4(G179), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT75), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n408), .A2(new_n409), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n411), .B1(new_n412), .B2(new_n296), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n300), .B1(new_n408), .B2(new_n409), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n410), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT18), .B1(new_n404), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n386), .A2(new_n389), .ZN(new_n417));
  INV_X1    g0217(.A(new_n379), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(KEYINPUT16), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(new_n275), .A3(new_n403), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n371), .B(KEYINPUT74), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n412), .A2(new_n296), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(KEYINPUT75), .A3(new_n414), .ZN(new_n424));
  INV_X1    g0224(.A(new_n410), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT18), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n422), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n416), .A2(new_n428), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n408), .A2(new_n364), .A3(new_n409), .ZN(new_n430));
  INV_X1    g0230(.A(new_n409), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n406), .A2(new_n407), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n431), .B1(new_n432), .B2(new_n252), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n430), .B1(G200), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n420), .A2(new_n434), .A3(new_n421), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT17), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n420), .A2(new_n434), .A3(KEYINPUT17), .A4(new_n421), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT76), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n437), .A2(KEYINPUT76), .A3(new_n438), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n429), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n367), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n326), .A2(KEYINPUT25), .A3(new_n227), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT25), .B1(new_n326), .B2(new_n227), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n254), .A2(G33), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n289), .A2(new_n447), .A3(new_n216), .A4(new_n273), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n445), .A2(new_n446), .B1(new_n227), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT24), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n222), .A2(G20), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT22), .B1(new_n260), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n217), .A2(G33), .A3(G116), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n227), .A2(KEYINPUT23), .A3(G20), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT23), .B1(new_n227), .B2(G20), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT22), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(new_n222), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n383), .A2(new_n217), .A3(new_n342), .A4(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n450), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n451), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n458), .B1(new_n345), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G116), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(G20), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT23), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(new_n217), .B2(G107), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n227), .A2(KEYINPUT23), .A3(G20), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND4_X1   g0269(.A1(new_n450), .A2(new_n460), .A3(new_n463), .A4(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n275), .B1(new_n461), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT84), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(KEYINPUT84), .B(new_n275), .C1(new_n461), .C2(new_n470), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n449), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g0275(.A1(G257), .A2(G1698), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n383), .A2(KEYINPUT85), .A3(new_n342), .A4(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n383), .A2(G250), .A3(new_n262), .A4(new_n342), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G294), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n342), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n394), .A2(new_n395), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(G33), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT85), .B1(new_n483), .B2(new_n476), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n265), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G45), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(G1), .ZN(new_n487));
  AND2_X1   g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  NOR2_X1   g0288(.A1(KEYINPUT5), .A2(G41), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n490), .A2(new_n252), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G264), .ZN(new_n492));
  XNOR2_X1  g0292(.A(KEYINPUT5), .B(G41), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n493), .A2(G274), .A3(new_n252), .A4(new_n487), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n485), .A2(new_n364), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n485), .A2(new_n492), .A3(new_n494), .ZN(new_n496));
  AOI22_X1  g0296(.A1(KEYINPUT86), .A2(new_n495), .B1(new_n496), .B2(new_n268), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n496), .A2(KEYINPUT86), .A3(new_n268), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n475), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT87), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n475), .B(KEYINPUT87), .C1(new_n497), .C2(new_n498), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(G257), .A2(G1698), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(new_n228), .B2(G1698), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(new_n383), .A3(new_n342), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n345), .A2(G303), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT80), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n506), .A2(KEYINPUT80), .A3(new_n507), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n265), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n490), .A2(G270), .A3(new_n252), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n513), .A2(KEYINPUT79), .A3(new_n494), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT79), .B1(new_n513), .B2(new_n494), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n289), .A2(new_n447), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT81), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n518), .A2(new_n519), .A3(G116), .A4(new_n274), .ZN(new_n520));
  INV_X1    g0320(.A(G116), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT81), .B1(new_n448), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n326), .A2(new_n521), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n273), .A2(new_n216), .B1(G20), .B2(new_n521), .ZN(new_n526));
  NOR2_X1   g0326(.A1(KEYINPUT82), .A2(KEYINPUT20), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G283), .ZN(new_n528));
  INV_X1    g0328(.A(G97), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n528), .B(new_n217), .C1(G33), .C2(new_n529), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n526), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n527), .B1(new_n526), .B2(new_n530), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT82), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT20), .ZN(new_n534));
  OAI22_X1  g0334(.A1(new_n531), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n300), .B1(new_n525), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT21), .B1(new_n517), .B2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n274), .A2(G116), .A3(new_n447), .A4(new_n289), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n538), .A2(KEYINPUT81), .B1(new_n521), .B2(new_n326), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n520), .A3(new_n539), .ZN(new_n540));
  AND4_X1   g0340(.A1(G179), .A2(new_n512), .A3(new_n540), .A4(new_n516), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n533), .A2(new_n534), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n526), .A2(new_n530), .ZN(new_n544));
  INV_X1    g0344(.A(new_n527), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n526), .A2(new_n527), .A3(new_n530), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n543), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(G169), .B1(new_n548), .B2(new_n524), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n512), .B2(new_n516), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT83), .B1(new_n550), .B2(KEYINPUT21), .ZN(new_n551));
  AND4_X1   g0351(.A1(KEYINPUT83), .A2(new_n517), .A3(new_n536), .A4(KEYINPUT21), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n542), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n354), .A2(new_n289), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n448), .A2(new_n222), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT19), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n282), .A2(new_n556), .A3(G97), .ZN(new_n557));
  NOR2_X1   g0357(.A1(G97), .A2(G107), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n558), .A2(new_n222), .B1(new_n304), .B2(new_n217), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n557), .B1(new_n559), .B2(new_n556), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n383), .A2(new_n217), .A3(G68), .A4(new_n342), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI211_X1 g0362(.A(new_n554), .B(new_n555), .C1(new_n562), .C2(new_n275), .ZN(new_n563));
  NOR2_X1   g0363(.A1(G238), .A2(G1698), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n226), .B2(G1698), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n565), .A2(new_n383), .A3(new_n342), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n252), .B1(new_n566), .B2(new_n464), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n487), .A2(new_n223), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n252), .ZN(new_n569));
  INV_X1    g0369(.A(new_n487), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n569), .B1(new_n570), .B2(new_n253), .ZN(new_n571));
  OAI21_X1  g0371(.A(G200), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n253), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(new_n487), .B1(new_n252), .B2(new_n568), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n566), .A2(new_n464), .ZN(new_n575));
  OAI211_X1 g0375(.A(G190), .B(new_n574), .C1(new_n575), .C2(new_n252), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n563), .A2(new_n572), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n562), .A2(new_n275), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n518), .A2(new_n354), .A3(new_n274), .ZN(new_n579));
  INV_X1    g0379(.A(new_n554), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n296), .B(new_n574), .C1(new_n575), .C2(new_n252), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n300), .B1(new_n567), .B2(new_n571), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n506), .A2(KEYINPUT80), .A3(new_n507), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT80), .B1(new_n506), .B2(new_n507), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n586), .A2(new_n587), .A3(new_n252), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n513), .A2(new_n494), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT79), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n513), .A2(KEYINPUT79), .A3(new_n494), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(G200), .B1(new_n588), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n540), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n512), .A2(new_n516), .A3(G190), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n260), .A2(G250), .A3(G1698), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT4), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(new_n226), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n600), .A2(new_n262), .A3(new_n342), .A4(new_n344), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(new_n528), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n383), .A2(G244), .A3(new_n262), .A4(new_n342), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n599), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n252), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n491), .A2(G257), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n494), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n300), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n494), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(G257), .B2(new_n491), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n602), .B1(new_n599), .B2(new_n604), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n296), .B(new_n611), .C1(new_n612), .C2(new_n252), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n227), .B1(new_n400), .B2(new_n401), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT6), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n529), .A2(new_n227), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n616), .B1(new_n617), .B2(new_n558), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n227), .A2(KEYINPUT6), .A3(G97), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G20), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n285), .A2(G77), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n622), .B(KEYINPUT77), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n274), .B1(new_n615), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n448), .A2(G97), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(G97), .B2(new_n326), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n627), .B(KEYINPUT78), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n609), .B(new_n613), .C1(new_n625), .C2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(G200), .B1(new_n606), .B2(new_n608), .ZN(new_n630));
  OAI211_X1 g0430(.A(G190), .B(new_n611), .C1(new_n612), .C2(new_n252), .ZN(new_n631));
  INV_X1    g0431(.A(new_n620), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n623), .B1(new_n632), .B2(new_n217), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n275), .B1(new_n633), .B2(new_n614), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT78), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n627), .B(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n630), .A2(new_n631), .A3(new_n634), .A4(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n585), .A2(new_n597), .A3(new_n629), .A4(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n496), .A2(new_n300), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n485), .A2(new_n296), .A3(new_n492), .A4(new_n494), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n475), .A2(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n553), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n444), .A2(new_n503), .A3(new_n643), .ZN(G372));
  AND2_X1   g0444(.A1(new_n416), .A2(new_n428), .ZN(new_n645));
  INV_X1    g0445(.A(new_n361), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n334), .B1(new_n338), .B2(new_n646), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n437), .A2(KEYINPUT76), .A3(new_n438), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n648), .A2(new_n439), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n645), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n295), .ZN(new_n651));
  INV_X1    g0451(.A(new_n629), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT26), .B1(new_n652), .B2(new_n585), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n577), .A2(new_n584), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n629), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n584), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n585), .A2(new_n629), .A3(new_n637), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n512), .A2(new_n540), .A3(new_n516), .A4(G179), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n550), .B2(KEYINPUT21), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n517), .A2(new_n536), .A3(KEYINPUT21), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT83), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n550), .A2(KEYINPUT83), .A3(KEYINPUT21), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n660), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n475), .A2(new_n641), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n658), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n657), .B1(new_n667), .B2(new_n503), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n298), .B(new_n651), .C1(new_n443), .C2(new_n668), .ZN(G369));
  NAND3_X1  g0469(.A1(new_n254), .A2(new_n217), .A3(G13), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n595), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n553), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n597), .ZN(new_n679));
  INV_X1    g0479(.A(G330), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n666), .A2(new_n675), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n475), .A2(new_n676), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n503), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n682), .B1(new_n684), .B2(new_n666), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n666), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n665), .A2(new_n675), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n682), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n686), .A2(new_n689), .ZN(G399));
  INV_X1    g0490(.A(new_n210), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G41), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n558), .A2(new_n222), .A3(new_n521), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n692), .A2(new_n693), .A3(new_n254), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n215), .B2(new_n692), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT28), .Z(new_n696));
  NAND2_X1  g0496(.A1(new_n667), .A2(new_n503), .ZN(new_n697));
  INV_X1    g0497(.A(new_n657), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n675), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(KEYINPUT91), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT29), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT31), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n643), .B2(new_n503), .ZN(new_n703));
  NOR4_X1   g0503(.A1(new_n517), .A2(new_n296), .A3(new_n606), .A4(new_n608), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT88), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n567), .A2(new_n571), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n485), .A2(new_n705), .A3(new_n706), .A4(new_n492), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n485), .A2(new_n492), .A3(new_n706), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT88), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n704), .A2(KEYINPUT30), .A3(new_n707), .A4(new_n709), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n588), .A2(new_n593), .A3(new_n296), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n606), .A2(new_n608), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n709), .A2(new_n711), .A3(new_n712), .A4(new_n707), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n296), .B1(new_n567), .B2(new_n571), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(new_n496), .A3(new_n517), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n710), .A2(new_n715), .A3(new_n702), .A4(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n719), .A2(new_n675), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n703), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n676), .A2(new_n702), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n717), .A2(new_n496), .A3(new_n517), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n714), .B2(new_n713), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT89), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n710), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n715), .A2(new_n718), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(KEYINPUT89), .ZN(new_n728));
  OAI211_X1 g0528(.A(KEYINPUT90), .B(new_n722), .C1(new_n726), .C2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n722), .B1(new_n726), .B2(new_n728), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT90), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n721), .A2(new_n729), .A3(new_n732), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n733), .A2(G330), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n701), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n696), .B1(new_n735), .B2(G1), .ZN(G364));
  INV_X1    g0536(.A(new_n679), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G13), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n740), .A2(new_n486), .A3(G20), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT92), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n742), .A2(new_n254), .A3(new_n692), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n681), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n217), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT95), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT97), .Z(new_n748));
  OR2_X1    g0548(.A1(new_n737), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n217), .A2(new_n296), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(G190), .A3(new_n268), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G179), .A2(G200), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(G20), .A3(new_n364), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n752), .A2(G322), .B1(G329), .B2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G311), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G190), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n750), .A2(new_n758), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n756), .B(new_n345), .C1(new_n757), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n750), .A2(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G190), .ZN(new_n762));
  INV_X1    g0562(.A(G317), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(KEYINPUT33), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n763), .A2(KEYINPUT33), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n762), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n761), .A2(new_n364), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G326), .ZN(new_n768));
  INV_X1    g0568(.A(G303), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n217), .A2(G179), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n766), .B(new_n768), .C1(new_n769), .C2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n770), .A2(new_n364), .A3(G200), .ZN(new_n773));
  INV_X1    g0573(.A(G283), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n217), .B1(new_n753), .B2(G190), .ZN(new_n775));
  INV_X1    g0575(.A(G294), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n773), .A2(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n760), .A2(new_n772), .A3(new_n777), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n751), .A2(new_n202), .B1(new_n759), .B2(new_n206), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT96), .ZN(new_n780));
  INV_X1    g0580(.A(new_n767), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n260), .B1(new_n781), .B2(new_n201), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n773), .A2(new_n227), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n771), .A2(new_n222), .ZN(new_n784));
  NOR4_X1   g0584(.A1(new_n780), .A2(new_n782), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n755), .A2(G159), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT32), .ZN(new_n787));
  INV_X1    g0587(.A(new_n762), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n788), .A2(new_n203), .B1(new_n775), .B2(new_n529), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n778), .B1(new_n785), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n216), .B1(G20), .B2(new_n300), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n743), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n691), .A2(new_n345), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n795), .A2(G355), .B1(new_n521), .B2(new_n691), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n384), .A2(new_n210), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT93), .Z(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n215), .A2(new_n486), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n249), .B2(new_n486), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n796), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n802), .A2(KEYINPUT94), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n747), .A2(new_n793), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(new_n802), .B2(KEYINPUT94), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n794), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n739), .A2(new_n744), .B1(new_n749), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  NOR2_X1   g0608(.A1(new_n792), .A2(new_n745), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n743), .B1(G77), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n773), .A2(new_n222), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n771), .A2(new_n227), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n812), .B(new_n813), .C1(G303), .C2(new_n767), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n260), .B1(new_n752), .B2(G294), .ZN(new_n815));
  INV_X1    g0615(.A(new_n759), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n816), .A2(G116), .B1(new_n755), .B2(G311), .ZN(new_n817));
  INV_X1    g0617(.A(new_n775), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n762), .A2(G283), .B1(G97), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n814), .A2(new_n815), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n773), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(G68), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n822), .B1(new_n201), .B2(new_n771), .C1(new_n202), .C2(new_n775), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n384), .B(new_n823), .C1(G132), .C2(new_n755), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n752), .A2(G143), .B1(new_n816), .B2(G159), .ZN(new_n825));
  INV_X1    g0625(.A(G137), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n825), .B1(new_n781), .B2(new_n826), .C1(new_n284), .C2(new_n788), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT34), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n827), .A2(new_n828), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n820), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n811), .B1(new_n832), .B2(new_n792), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n361), .A2(new_n675), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n365), .B1(new_n362), .B2(new_n676), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n361), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n745), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n833), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n668), .A2(new_n838), .A3(new_n675), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(KEYINPUT98), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n699), .A2(new_n839), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n843), .B(new_n844), .Z(new_n845));
  AND2_X1   g0645(.A1(new_n845), .A2(new_n734), .ZN(new_n846));
  INV_X1    g0646(.A(new_n743), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n845), .B2(new_n734), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n841), .B1(new_n846), .B2(new_n848), .ZN(G384));
  OR2_X1    g0649(.A1(new_n620), .A2(KEYINPUT35), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n620), .A2(KEYINPUT35), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n850), .A2(G116), .A3(new_n218), .A4(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT36), .Z(new_n853));
  NAND4_X1  g0653(.A1(new_n215), .A2(G77), .A3(new_n375), .A4(new_n376), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n254), .B(G13), .C1(new_n854), .C2(new_n245), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n701), .A2(new_n444), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n651), .A2(new_n298), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n645), .B1(new_n648), .B2(new_n439), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n390), .A2(KEYINPUT16), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n373), .B1(new_n861), .B2(new_n391), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(new_n673), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n435), .B1(new_n862), .B2(new_n673), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n862), .A2(new_n415), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT37), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n422), .A2(new_n426), .ZN(new_n868));
  INV_X1    g0668(.A(new_n673), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n422), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n868), .A2(new_n870), .A3(new_n871), .A4(new_n435), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n864), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT38), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n864), .A2(KEYINPUT38), .A3(new_n873), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n331), .A2(new_n676), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n339), .B2(new_n321), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT99), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n321), .A2(new_n881), .A3(new_n332), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n319), .B1(new_n315), .B2(new_n316), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT99), .B1(new_n883), .B2(new_n331), .ZN(new_n884));
  INV_X1    g0684(.A(new_n879), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n882), .A2(new_n884), .A3(new_n338), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n878), .B(new_n887), .C1(new_n834), .C2(new_n842), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT39), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n416), .A2(new_n437), .A3(new_n428), .A4(new_n438), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n404), .A2(new_n673), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n890), .A2(KEYINPUT101), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT101), .B1(new_n890), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n435), .B1(new_n404), .B2(new_n415), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT37), .B1(new_n895), .B2(new_n891), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT100), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n896), .A2(new_n897), .A3(new_n872), .ZN(new_n898));
  OAI211_X1 g0698(.A(KEYINPUT100), .B(KEYINPUT37), .C1(new_n895), .C2(new_n891), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT38), .B1(new_n894), .B2(new_n900), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n864), .A2(KEYINPUT38), .A3(new_n873), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n889), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n876), .A2(KEYINPUT39), .A3(new_n877), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n882), .A2(new_n884), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n906), .A2(new_n675), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n888), .B1(new_n645), .B2(new_n869), .C1(new_n905), .C2(new_n908), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n859), .B(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n901), .A2(new_n902), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n838), .B1(new_n880), .B2(new_n886), .ZN(new_n912));
  INV_X1    g0712(.A(new_n710), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n722), .B1(new_n727), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n703), .B2(new_n720), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT40), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT40), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n878), .A2(new_n918), .A3(new_n915), .A4(new_n912), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n443), .B1(new_n721), .B2(new_n914), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n922), .A2(new_n923), .A3(new_n680), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n910), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(G1), .B1(new_n740), .B2(G20), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n910), .B2(new_n924), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n856), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT102), .Z(G367));
  INV_X1    g0729(.A(KEYINPUT104), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n675), .B1(new_n625), .B2(new_n628), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n629), .A2(new_n637), .A3(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n666), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n676), .B1(new_n933), .B2(new_n652), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT42), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n685), .A2(new_n688), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n652), .A2(new_n675), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n932), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n936), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n685), .A2(KEYINPUT42), .A3(new_n688), .A4(new_n939), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n935), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n584), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n563), .A2(new_n676), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n654), .B2(new_n945), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n947), .A2(KEYINPUT103), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT43), .B1(new_n947), .B2(KEYINPUT103), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n943), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT105), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT105), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n943), .B2(new_n953), .ZN(new_n957));
  INV_X1    g0757(.A(new_n950), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n943), .A2(new_n958), .ZN(new_n959));
  AND4_X1   g0759(.A1(new_n930), .A2(new_n955), .A3(new_n957), .A4(new_n959), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n954), .A2(KEYINPUT105), .B1(new_n943), .B2(new_n958), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n930), .B1(new_n961), .B2(new_n957), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n960), .A2(new_n962), .B1(new_n686), .B2(new_n940), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n957), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(KEYINPUT104), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n686), .A2(new_n940), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n961), .A2(new_n930), .A3(new_n957), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n692), .B(new_n969), .Z(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n689), .A2(new_n939), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT45), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(KEYINPUT45), .B1(new_n689), .B2(new_n939), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n689), .A2(new_n939), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT44), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n976), .A2(new_n978), .A3(new_n686), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n977), .A2(KEYINPUT44), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT44), .ZN(new_n981));
  NOR3_X1   g0781(.A1(new_n689), .A2(new_n981), .A3(new_n939), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n980), .A2(new_n982), .B1(new_n974), .B2(new_n975), .ZN(new_n983));
  INV_X1    g0783(.A(new_n686), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n737), .A2(G330), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT107), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n986), .A2(new_n987), .A3(new_n937), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n986), .B1(new_n937), .B2(new_n987), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n989), .A2(new_n990), .B1(new_n685), .B2(new_n688), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n937), .A2(new_n987), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n681), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n685), .A2(new_n688), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n993), .A2(new_n994), .A3(new_n988), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n991), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n979), .A2(new_n985), .A3(new_n735), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n971), .B1(new_n997), .B2(new_n735), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n742), .A2(new_n254), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n963), .B(new_n968), .C1(new_n998), .C2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n804), .B1(new_n691), .B2(new_n354), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n799), .B2(new_n236), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n743), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n775), .A2(new_n203), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n751), .A2(new_n284), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(G143), .C2(new_n767), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n1007), .A2(KEYINPUT108), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n260), .B1(new_n754), .B2(new_n826), .C1(new_n759), .C2(new_n201), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n821), .A2(G77), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n202), .B2(new_n771), .C1(new_n788), .C2(new_n378), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(KEYINPUT108), .B2(new_n1007), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n771), .A2(new_n521), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT46), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n776), .A2(new_n788), .B1(new_n781), .B2(new_n757), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G97), .B2(new_n821), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n751), .A2(new_n769), .B1(new_n759), .B2(new_n774), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G317), .B2(new_n755), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n483), .B1(G107), .B2(new_n818), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1017), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1013), .B1(new_n1015), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT47), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1004), .B1(new_n1023), .B2(new_n792), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n947), .A2(new_n748), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1001), .A2(new_n1026), .ZN(G387));
  NAND2_X1  g0827(.A1(new_n996), .A2(new_n1000), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n751), .A2(new_n201), .B1(new_n759), .B2(new_n203), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G150), .B2(new_n755), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n771), .A2(new_n206), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n368), .B2(new_n762), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n767), .A2(G159), .B1(new_n354), .B2(new_n818), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n384), .B1(G97), .B2(new_n821), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1030), .A2(new_n1032), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(G322), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n757), .A2(new_n788), .B1(new_n781), .B2(new_n1036), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1037), .A2(KEYINPUT110), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(KEYINPUT110), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n752), .A2(G317), .B1(new_n816), .B2(G303), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT48), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n771), .A2(new_n776), .B1(new_n775), .B2(new_n774), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1043), .A2(KEYINPUT49), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n483), .B1(G326), .B2(new_n755), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(new_n521), .C2(new_n773), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT49), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1035), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n792), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n795), .A2(new_n693), .B1(new_n227), .B2(new_n691), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n351), .A2(new_n201), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT50), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n486), .B1(new_n203), .B2(new_n206), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1054), .A2(new_n693), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n798), .B1(new_n240), .B2(new_n486), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1052), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1058), .A2(KEYINPUT109), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n804), .B1(new_n1058), .B2(KEYINPUT109), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n847), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1051), .B(new_n1061), .C1(new_n685), .C2(new_n748), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n996), .A2(new_n735), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n692), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n996), .A2(new_n735), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1028), .B(new_n1062), .C1(new_n1064), .C2(new_n1065), .ZN(G393));
  AND2_X1   g0866(.A1(new_n997), .A2(new_n692), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT111), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n979), .A2(new_n985), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n1063), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n692), .A3(new_n997), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT111), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n979), .A2(new_n985), .A3(new_n1000), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n781), .A2(new_n284), .B1(new_n378), .B2(new_n751), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT51), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n788), .A2(new_n201), .B1(new_n203), .B2(new_n771), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n775), .A2(new_n206), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n1078), .A2(new_n812), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n351), .A2(new_n816), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n384), .B1(G143), .B2(new_n755), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1077), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n781), .A2(new_n763), .B1(new_n757), .B2(new_n751), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT52), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n771), .A2(new_n774), .B1(new_n775), .B2(new_n521), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n783), .B(new_n1086), .C1(G303), .C2(new_n762), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n345), .B1(new_n754), .B2(new_n1036), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G294), .B2(new_n816), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n793), .B1(new_n1083), .B2(new_n1090), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n799), .A2(new_n244), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n804), .B1(G97), .B2(new_n691), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n847), .B(new_n1091), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n939), .B2(new_n747), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1075), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1074), .A2(new_n1096), .ZN(G390));
  INV_X1    g0897(.A(KEYINPUT115), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n722), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n913), .B1(new_n727), .B2(KEYINPUT89), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n724), .A2(new_n725), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n1102), .A2(KEYINPUT90), .B1(new_n703), .B2(new_n720), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n729), .ZN(new_n1104));
  OAI211_X1 g0904(.A(G330), .B(new_n912), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(KEYINPUT114), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT114), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n733), .A2(new_n1107), .A3(G330), .A4(new_n912), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n915), .A2(G330), .A3(new_n839), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n887), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(KEYINPUT112), .B1(new_n842), .B2(new_n834), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n834), .B1(new_n699), .B2(new_n839), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT112), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1112), .A2(new_n1113), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1098), .B1(new_n1109), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n733), .A2(G330), .A3(new_n839), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n1111), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n915), .A2(G330), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n912), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1114), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1118), .A2(new_n1124), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1109), .A2(new_n1117), .A3(new_n1098), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n858), .B(new_n857), .C1(new_n444), .C2(new_n1122), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n908), .B1(new_n1114), .B2(new_n1111), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(KEYINPUT113), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT113), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1133), .B(new_n908), .C1(new_n1114), .C2(new_n1111), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(new_n905), .A3(new_n1134), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n842), .A2(KEYINPUT112), .A3(new_n834), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n697), .A2(new_n698), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1137), .A2(new_n676), .A3(new_n839), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1115), .B1(new_n1138), .B2(new_n835), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n887), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n911), .A2(new_n907), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1135), .A2(new_n1142), .A3(new_n1109), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1131), .A2(KEYINPUT113), .B1(new_n903), .B2(new_n904), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1144), .A2(new_n1134), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1143), .B1(new_n1145), .B2(new_n1123), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1130), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1135), .A2(new_n1142), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1148), .A2(new_n912), .A3(new_n1122), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1128), .A2(new_n1129), .A3(new_n1143), .A4(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1147), .A2(new_n1150), .A3(new_n692), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n781), .A2(new_n774), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1079), .B(new_n1152), .C1(G107), .C2(new_n762), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n784), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n751), .A2(new_n521), .B1(new_n776), .B2(new_n754), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n260), .B(new_n1155), .C1(G97), .C2(new_n816), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1153), .A2(new_n1154), .A3(new_n822), .A4(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(G132), .ZN(new_n1158));
  INV_X1    g0958(.A(G125), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n751), .A2(new_n1158), .B1(new_n1159), .B2(new_n754), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT54), .B(G143), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n345), .B(new_n1160), .C1(new_n816), .C2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n771), .A2(new_n284), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT53), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n767), .A2(G128), .B1(new_n821), .B2(G50), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n762), .A2(G137), .B1(G159), .B2(new_n818), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1163), .A2(new_n1165), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT117), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1157), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n792), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1173), .B(new_n743), .C1(new_n368), .C2(new_n810), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n905), .B2(new_n745), .ZN(new_n1175));
  OR3_X1    g0975(.A1(new_n1146), .A2(KEYINPUT116), .A3(new_n999), .ZN(new_n1176));
  OAI21_X1  g0976(.A(KEYINPUT116), .B1(new_n1146), .B2(new_n999), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1151), .A2(new_n1178), .ZN(G378));
  NOR3_X1   g0979(.A1(new_n1126), .A2(new_n1118), .A3(new_n1124), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1129), .B1(new_n1180), .B2(new_n1146), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n299), .A2(new_n292), .A3(new_n869), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n292), .A2(new_n869), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n295), .A2(new_n298), .A3(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1182), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1185), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n920), .B2(G330), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n909), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n920), .A2(G330), .A3(new_n1189), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n680), .B(new_n1188), .C1(new_n917), .C2(new_n919), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n909), .B1(new_n1195), .B2(new_n1190), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1181), .A2(KEYINPUT57), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT57), .B1(new_n1181), .B2(new_n1197), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n692), .B(new_n1198), .C1(new_n1199), .C2(KEYINPUT121), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT121), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1201), .B(KEYINPUT57), .C1(new_n1181), .C2(new_n1197), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1188), .A2(new_n745), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n810), .A2(G50), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n752), .A2(G107), .B1(G283), .B2(new_n755), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1031), .A2(new_n1005), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n353), .C2(new_n759), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n767), .A2(G116), .B1(new_n821), .B2(G58), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n529), .B2(new_n788), .ZN(new_n1210));
  NOR4_X1   g1010(.A1(new_n1208), .A2(new_n1210), .A3(G41), .A4(new_n483), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT120), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1212), .A2(KEYINPUT58), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(KEYINPUT58), .ZN(new_n1214));
  INV_X1    g1014(.A(G41), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n281), .A2(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT118), .ZN(new_n1217));
  AOI211_X1 g1017(.A(G50), .B(new_n1217), .C1(new_n1215), .C2(new_n384), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT119), .Z(new_n1219));
  OAI22_X1  g1019(.A1(new_n1159), .A2(new_n781), .B1(new_n788), .B2(new_n1158), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G150), .B2(new_n818), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n752), .A2(G128), .B1(new_n816), .B2(G137), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1221), .B(new_n1222), .C1(new_n771), .C2(new_n1161), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n755), .A2(G124), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1217), .B(new_n1225), .C1(new_n378), .C2(new_n773), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1223), .B2(KEYINPUT59), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1219), .B1(new_n1224), .B2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1213), .A2(new_n1214), .A3(new_n1228), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n847), .B(new_n1205), .C1(new_n1229), .C2(new_n792), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1204), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1197), .B2(new_n1000), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1203), .A2(new_n1232), .ZN(G375));
  OAI22_X1  g1033(.A1(new_n521), .A2(new_n788), .B1(new_n781), .B2(new_n776), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n771), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1234), .B1(G97), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n818), .A2(new_n354), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n751), .A2(new_n774), .B1(new_n759), .B2(new_n227), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n260), .B(new_n1238), .C1(G303), .C2(new_n755), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1236), .A2(new_n1010), .A3(new_n1237), .A4(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(G128), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n759), .A2(new_n284), .B1(new_n754), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G137), .B2(new_n752), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n767), .A2(G132), .B1(new_n1235), .B2(G159), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n762), .A2(new_n1162), .B1(G50), .B2(new_n818), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n384), .B1(G58), .B2(new_n821), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n793), .B1(new_n1240), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n743), .B1(G68), .B2(new_n810), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1248), .B(new_n1249), .C1(new_n1111), .C2(new_n745), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1128), .B2(new_n1000), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT122), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n859), .B1(new_n443), .B2(new_n1121), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1180), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1130), .A2(new_n1254), .A3(new_n970), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1252), .A2(new_n1255), .ZN(G381));
  OR4_X1    g1056(.A1(G396), .A2(G378), .A3(G384), .A4(G393), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1001), .A2(new_n1026), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1075), .A2(new_n1095), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  OR4_X1    g1061(.A1(G375), .A2(new_n1257), .A3(G381), .A4(new_n1261), .ZN(G407));
  INV_X1    g1062(.A(G378), .ZN(new_n1263));
  INV_X1    g1063(.A(G213), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1264), .A2(G343), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G407), .B(G213), .C1(G375), .C2(new_n1266), .ZN(G409));
  INV_X1    g1067(.A(KEYINPUT124), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G390), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1260), .A2(KEYINPUT124), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(G387), .A3(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(G393), .B(new_n807), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT125), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(new_n1258), .B2(G390), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(G387), .A2(KEYINPUT125), .A3(new_n1260), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1271), .B(new_n1273), .C1(new_n1275), .C2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(G387), .A2(G390), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1261), .A2(new_n1272), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G378), .B(new_n1232), .C1(new_n1200), .C2(new_n1202), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1232), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1181), .A2(new_n970), .A3(new_n1197), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1151), .B(new_n1178), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1265), .B1(new_n1282), .B2(new_n1285), .ZN(new_n1286));
  XOR2_X1   g1086(.A(G384), .B(KEYINPUT123), .Z(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT122), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1251), .B(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1180), .A2(KEYINPUT60), .A3(new_n1253), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n692), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1130), .A2(KEYINPUT60), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1254), .B2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1288), .B1(new_n1290), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(new_n1254), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1292), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  OR2_X1    g1098(.A1(G384), .A2(KEYINPUT123), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n1252), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1295), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(KEYINPUT62), .B1(new_n1286), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT126), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1282), .A2(new_n1285), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1265), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1304), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  AOI211_X1 g1107(.A(KEYINPUT126), .B(new_n1265), .C1(new_n1282), .C2(new_n1285), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1302), .A2(KEYINPUT62), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1303), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1265), .A2(G2897), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1295), .A2(new_n1300), .A3(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1312), .B1(new_n1295), .B2(new_n1300), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1316), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT61), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1281), .B1(new_n1311), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1315), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1313), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1280), .B(new_n1318), .C1(new_n1322), .C2(new_n1286), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT63), .B1(new_n1286), .B2(new_n1302), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1309), .A2(KEYINPUT63), .A3(new_n1302), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1320), .A2(new_n1327), .ZN(G405));
  NAND2_X1  g1128(.A1(new_n1280), .A2(KEYINPUT127), .ZN(new_n1329));
  AOI21_X1  g1129(.A(G378), .B1(new_n1203), .B2(new_n1232), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1282), .ZN(new_n1331));
  OR3_X1    g1131(.A1(new_n1330), .A2(new_n1302), .A3(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1302), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1329), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1280), .A2(KEYINPUT127), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(new_n1334), .B(new_n1335), .ZN(G402));
endmodule


