

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801;

  BUF_X1 U378 ( .A(n700), .Z(n356) );
  AND2_X1 U379 ( .A1(n384), .A2(n385), .ZN(n383) );
  AND2_X1 U380 ( .A1(n381), .A2(n380), .ZN(n432) );
  NAND2_X1 U381 ( .A1(n411), .A2(n454), .ZN(n641) );
  OR2_X1 U382 ( .A1(n647), .A2(n646), .ZN(n749) );
  NAND2_X1 U383 ( .A1(n370), .A2(n688), .ZN(n621) );
  NOR2_X1 U384 ( .A1(n672), .A2(n671), .ZN(n564) );
  AND2_X1 U385 ( .A1(n357), .A2(n469), .ZN(n365) );
  INV_X1 U386 ( .A(KEYINPUT34), .ZN(n353) );
  OR2_X2 U387 ( .A1(n409), .A2(n407), .ZN(n372) );
  NAND2_X1 U388 ( .A1(n408), .A2(n452), .ZN(n407) );
  XOR2_X1 U389 ( .A(n531), .B(n530), .Z(n374) );
  XNOR2_X1 U390 ( .A(n528), .B(n514), .ZN(n732) );
  XNOR2_X1 U391 ( .A(n522), .B(n521), .ZN(n781) );
  INV_X1 U392 ( .A(G953), .ZN(n793) );
  XNOR2_X1 U393 ( .A(n373), .B(n374), .ZN(n371) );
  AND2_X1 U394 ( .A1(n633), .A2(n353), .ZN(n354) );
  NAND2_X2 U395 ( .A1(n633), .A2(n626), .ZN(n627) );
  XNOR2_X2 U396 ( .A(n618), .B(n617), .ZN(n370) );
  NOR2_X2 U397 ( .A1(n739), .A2(n774), .ZN(n740) );
  XNOR2_X2 U398 ( .A(n618), .B(n617), .ZN(n633) );
  AND2_X2 U399 ( .A1(n716), .A2(G953), .ZN(n774) );
  XNOR2_X2 U400 ( .A(n581), .B(KEYINPUT19), .ZN(n615) );
  NAND2_X2 U401 ( .A1(n615), .A2(n614), .ZN(n618) );
  AND2_X2 U402 ( .A1(n423), .A2(n422), .ZN(n376) );
  NAND2_X1 U403 ( .A1(n611), .A2(n610), .ZN(n662) );
  NAND2_X2 U404 ( .A1(n580), .A2(n681), .ZN(n764) );
  NAND2_X1 U405 ( .A1(n354), .A2(n415), .ZN(n413) );
  XNOR2_X2 U406 ( .A(G116), .B(G113), .ZN(n447) );
  NAND2_X1 U407 ( .A1(n355), .A2(n432), .ZN(n430) );
  NOR2_X2 U408 ( .A1(n429), .A2(n428), .ZN(n355) );
  NOR2_X2 U409 ( .A1(n594), .A2(n755), .ZN(n462) );
  NOR2_X2 U410 ( .A1(n488), .A2(n565), .ZN(n518) );
  OR2_X2 U411 ( .A1(n595), .A2(n607), .ZN(n597) );
  XNOR2_X1 U412 ( .A(n449), .B(n466), .ZN(n448) );
  NAND2_X2 U413 ( .A1(n629), .A2(n426), .ZN(n643) );
  XNOR2_X2 U414 ( .A(n528), .B(n404), .ZN(n735) );
  NAND2_X1 U415 ( .A1(n757), .A2(n751), .ZN(n624) );
  XNOR2_X1 U416 ( .A(n465), .B(KEYINPUT82), .ZN(n758) );
  OR2_X1 U417 ( .A1(n599), .A2(n584), .ZN(n757) );
  XNOR2_X2 U418 ( .A(n446), .B(n444), .ZN(n522) );
  XNOR2_X2 U419 ( .A(n570), .B(KEYINPUT111), .ZN(n583) );
  XNOR2_X2 U420 ( .A(n510), .B(n509), .ZN(n528) );
  AND2_X2 U421 ( .A1(n651), .A2(n650), .ZN(n393) );
  AND2_X2 U422 ( .A1(n413), .A2(n412), .ZN(n411) );
  XNOR2_X2 U423 ( .A(n478), .B(n477), .ZN(n713) );
  NAND2_X2 U424 ( .A1(n376), .A2(n419), .ZN(n723) );
  AND2_X1 U425 ( .A1(n455), .A2(n639), .ZN(n454) );
  INV_X1 U426 ( .A(n624), .ZN(n673) );
  INV_X1 U427 ( .A(n757), .ZN(n421) );
  INV_X1 U428 ( .A(n563), .ZN(n669) );
  INV_X1 U429 ( .A(n628), .ZN(n357) );
  AND2_X1 U430 ( .A1(n601), .A2(n600), .ZN(n755) );
  AND2_X1 U431 ( .A1(n418), .A2(n439), .ZN(n377) );
  NOR2_X1 U432 ( .A1(n356), .A2(n699), .ZN(n701) );
  INV_X1 U433 ( .A(n619), .ZN(n358) );
  XNOR2_X1 U434 ( .A(n437), .B(G125), .ZN(n526) );
  XOR2_X1 U435 ( .A(KEYINPUT73), .B(G131), .Z(n550) );
  BUF_X1 U436 ( .A(n662), .Z(n359) );
  BUF_X1 U437 ( .A(n382), .Z(n360) );
  XNOR2_X1 U438 ( .A(n735), .B(n736), .ZN(n737) );
  AND2_X2 U439 ( .A1(n370), .A2(n623), .ZN(n744) );
  NAND2_X2 U440 ( .A1(n371), .A2(n668), .ZN(n581) );
  XNOR2_X1 U441 ( .A(n445), .B(G119), .ZN(n444) );
  XNOR2_X1 U442 ( .A(n447), .B(n472), .ZN(n446) );
  INV_X1 U443 ( .A(KEYINPUT74), .ZN(n445) );
  NOR2_X1 U444 ( .A1(n770), .A2(G902), .ZN(n503) );
  AND2_X1 U445 ( .A1(n624), .A2(n443), .ZN(n442) );
  INV_X1 U446 ( .A(KEYINPUT104), .ZN(n443) );
  AND2_X1 U447 ( .A1(n624), .A2(n369), .ZN(n463) );
  INV_X1 U448 ( .A(KEYINPUT86), .ZN(n467) );
  INV_X1 U449 ( .A(n480), .ZN(n453) );
  NAND2_X1 U450 ( .A1(n480), .A2(G902), .ZN(n452) );
  NOR2_X1 U451 ( .A1(n480), .A2(G902), .ZN(n451) );
  XNOR2_X1 U452 ( .A(KEYINPUT71), .B(KEYINPUT4), .ZN(n470) );
  XNOR2_X1 U453 ( .A(n402), .B(n653), .ZN(n707) );
  NAND2_X1 U454 ( .A1(n387), .A2(n383), .ZN(n402) );
  XNOR2_X1 U455 ( .A(G119), .B(G110), .ZN(n489) );
  XNOR2_X1 U456 ( .A(G128), .B(G137), .ZN(n492) );
  XNOR2_X1 U457 ( .A(n550), .B(n473), .ZN(n792) );
  XNOR2_X1 U458 ( .A(G137), .B(G134), .ZN(n473) );
  XNOR2_X1 U459 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n523) );
  XNOR2_X1 U460 ( .A(n427), .B(n527), .ZN(n406) );
  INV_X1 U461 ( .A(n526), .ZN(n427) );
  XNOR2_X1 U462 ( .A(n520), .B(G122), .ZN(n521) );
  XOR2_X1 U463 ( .A(KEYINPUT16), .B(KEYINPUT78), .Z(n520) );
  XNOR2_X1 U464 ( .A(G122), .B(KEYINPUT102), .ZN(n533) );
  XOR2_X1 U465 ( .A(KEYINPUT101), .B(KEYINPUT9), .Z(n534) );
  XNOR2_X1 U466 ( .A(n536), .B(n535), .ZN(n537) );
  INV_X1 U467 ( .A(KEYINPUT7), .ZN(n535) );
  XNOR2_X1 U468 ( .A(G116), .B(G107), .ZN(n536) );
  XNOR2_X1 U469 ( .A(n547), .B(n546), .ZN(n599) );
  XNOR2_X1 U470 ( .A(G478), .B(KEYINPUT103), .ZN(n546) );
  NOR2_X1 U471 ( .A1(n767), .A2(G902), .ZN(n547) );
  INV_X1 U472 ( .A(KEYINPUT22), .ZN(n401) );
  XNOR2_X1 U473 ( .A(n499), .B(n498), .ZN(n770) );
  INV_X1 U474 ( .A(n790), .ZN(n498) );
  OR2_X1 U475 ( .A1(n587), .A2(n589), .ZN(n588) );
  OR2_X1 U476 ( .A1(n624), .A2(n443), .ZN(n440) );
  INV_X1 U477 ( .A(KEYINPUT79), .ZN(n398) );
  NAND2_X1 U478 ( .A1(n458), .A2(n461), .ZN(n457) );
  INV_X1 U479 ( .A(G237), .ZN(n481) );
  XNOR2_X1 U480 ( .A(G902), .B(KEYINPUT15), .ZN(n709) );
  INV_X1 U481 ( .A(KEYINPUT85), .ZN(n466) );
  XNOR2_X1 U482 ( .A(n435), .B(n434), .ZN(n603) );
  INV_X1 U483 ( .A(KEYINPUT108), .ZN(n434) );
  OR2_X1 U484 ( .A1(n679), .A2(n678), .ZN(n619) );
  XNOR2_X1 U485 ( .A(G110), .B(G107), .ZN(n508) );
  XNOR2_X1 U486 ( .A(n495), .B(n395), .ZN(n540) );
  XNOR2_X1 U487 ( .A(n396), .B(KEYINPUT72), .ZN(n395) );
  INV_X1 U488 ( .A(KEYINPUT8), .ZN(n396) );
  INV_X1 U489 ( .A(KEYINPUT23), .ZN(n491) );
  NOR2_X1 U490 ( .A1(G953), .A2(G237), .ZN(n548) );
  XNOR2_X1 U491 ( .A(G113), .B(G122), .ZN(n552) );
  XOR2_X1 U492 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n553) );
  XNOR2_X1 U493 ( .A(n526), .B(n436), .ZN(n790) );
  XNOR2_X1 U494 ( .A(G140), .B(KEYINPUT10), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n781), .B(n405), .ZN(n404) );
  XNOR2_X1 U496 ( .A(n406), .B(n525), .ZN(n405) );
  NAND2_X1 U497 ( .A1(n421), .A2(n468), .ZN(n420) );
  NAND2_X1 U498 ( .A1(n757), .A2(n424), .ZN(n422) );
  XNOR2_X1 U499 ( .A(n603), .B(n433), .ZN(n576) );
  INV_X1 U500 ( .A(KEYINPUT116), .ZN(n433) );
  NAND2_X1 U501 ( .A1(n568), .A2(n358), .ZN(n622) );
  INV_X1 U502 ( .A(n795), .ZN(n410) );
  XNOR2_X1 U503 ( .A(n543), .B(n397), .ZN(n544) );
  XNOR2_X1 U504 ( .A(n538), .B(n537), .ZN(n539) );
  BUF_X1 U505 ( .A(n760), .Z(n394) );
  BUF_X1 U506 ( .A(n758), .Z(n399) );
  NOR2_X1 U507 ( .A1(n630), .A2(n357), .ZN(n425) );
  XNOR2_X1 U508 ( .A(n770), .B(KEYINPUT124), .ZN(n771) );
  AND2_X1 U509 ( .A1(n703), .A2(n793), .ZN(n400) );
  AND2_X1 U510 ( .A1(n712), .A2(G475), .ZN(n361) );
  INV_X1 U511 ( .A(G902), .ZN(n515) );
  AND2_X1 U512 ( .A1(n378), .A2(G469), .ZN(n362) );
  AND2_X1 U513 ( .A1(n375), .A2(n361), .ZN(n363) );
  AND2_X1 U514 ( .A1(n419), .A2(n461), .ZN(n364) );
  AND2_X1 U515 ( .A1(n681), .A2(n679), .ZN(n366) );
  INV_X1 U516 ( .A(G146), .ZN(n437) );
  XOR2_X1 U517 ( .A(KEYINPUT105), .B(KEYINPUT6), .Z(n367) );
  XOR2_X1 U518 ( .A(KEYINPUT67), .B(KEYINPUT1), .Z(n368) );
  XOR2_X1 U519 ( .A(KEYINPUT70), .B(KEYINPUT47), .Z(n369) );
  XNOR2_X1 U520 ( .A(n560), .B(n559), .ZN(n598) );
  NAND2_X1 U521 ( .A1(n390), .A2(n389), .ZN(n388) );
  XNOR2_X1 U522 ( .A(n373), .B(n374), .ZN(n575) );
  NOR2_X2 U523 ( .A1(n735), .A2(n706), .ZN(n373) );
  OR2_X1 U524 ( .A1(n407), .A2(n409), .ZN(n684) );
  XNOR2_X1 U525 ( .A(n494), .B(n493), .ZN(n497) );
  NAND2_X1 U526 ( .A1(n448), .A2(n711), .ZN(n375) );
  NAND2_X1 U527 ( .A1(n448), .A2(n711), .ZN(n403) );
  XNOR2_X1 U528 ( .A(n386), .B(KEYINPUT107), .ZN(n385) );
  NAND2_X1 U529 ( .A1(n800), .A2(n649), .ZN(n392) );
  NAND2_X1 U530 ( .A1(n713), .A2(n451), .ZN(n408) );
  AND2_X1 U531 ( .A1(n375), .A2(n712), .ZN(n378) );
  AND2_X2 U532 ( .A1(n403), .A2(n712), .ZN(n769) );
  BUF_X1 U533 ( .A(n581), .Z(n379) );
  BUF_X1 U534 ( .A(n707), .Z(n775) );
  NAND2_X1 U535 ( .A1(n725), .A2(n749), .ZN(n651) );
  AND2_X1 U536 ( .A1(n629), .A2(n425), .ZN(n741) );
  NAND2_X1 U537 ( .A1(n364), .A2(n376), .ZN(n380) );
  NAND2_X1 U538 ( .A1(n460), .A2(n723), .ZN(n381) );
  AND2_X1 U539 ( .A1(n382), .A2(n775), .ZN(n654) );
  NOR2_X1 U540 ( .A1(n658), .A2(n360), .ZN(n659) );
  NAND2_X1 U541 ( .A1(n450), .A2(n382), .ZN(n449) );
  XNOR2_X1 U542 ( .A(n360), .B(n410), .ZN(n794) );
  XNOR2_X2 U543 ( .A(n662), .B(KEYINPUT89), .ZN(n382) );
  XNOR2_X2 U544 ( .A(n568), .B(n368), .ZN(n681) );
  XNOR2_X2 U545 ( .A(n516), .B(G469), .ZN(n568) );
  OR2_X2 U546 ( .A1(n800), .A2(n650), .ZN(n384) );
  NAND2_X1 U547 ( .A1(n632), .A2(n631), .ZN(n386) );
  NAND2_X1 U548 ( .A1(n391), .A2(n388), .ZN(n387) );
  NAND2_X1 U549 ( .A1(n800), .A2(n648), .ZN(n389) );
  INV_X1 U550 ( .A(n651), .ZN(n390) );
  NAND2_X1 U551 ( .A1(n393), .A2(n392), .ZN(n391) );
  XNOR2_X2 U552 ( .A(n641), .B(n640), .ZN(n800) );
  NOR2_X1 U553 ( .A1(n713), .A2(n453), .ZN(n409) );
  INV_X1 U554 ( .A(n542), .ZN(n397) );
  XNOR2_X1 U555 ( .A(n585), .B(n398), .ZN(n459) );
  XNOR2_X2 U556 ( .A(n573), .B(n572), .ZN(n801) );
  AND2_X1 U557 ( .A1(n441), .A2(n440), .ZN(n439) );
  NOR2_X1 U558 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U559 ( .A1(n656), .A2(n655), .ZN(n660) );
  NAND2_X1 U560 ( .A1(n667), .A2(n400), .ZN(n705) );
  INV_X1 U561 ( .A(n629), .ZN(n647) );
  XNOR2_X2 U562 ( .A(n627), .B(n401), .ZN(n629) );
  XNOR2_X2 U563 ( .A(n789), .B(n471), .ZN(n510) );
  XNOR2_X2 U564 ( .A(n542), .B(n470), .ZN(n789) );
  NAND2_X1 U565 ( .A1(n700), .A2(KEYINPUT34), .ZN(n412) );
  INV_X1 U566 ( .A(n700), .ZN(n415) );
  NOR2_X1 U567 ( .A1(n628), .A2(n619), .ZN(n634) );
  XNOR2_X2 U568 ( .A(n372), .B(n367), .ZN(n628) );
  NAND2_X1 U569 ( .A1(n377), .A2(n416), .ZN(n632) );
  NAND2_X1 U570 ( .A1(n417), .A2(n438), .ZN(n416) );
  INV_X1 U571 ( .A(n760), .ZN(n417) );
  NAND2_X1 U572 ( .A1(n760), .A2(n442), .ZN(n418) );
  OR2_X1 U573 ( .A1(n609), .A2(n420), .ZN(n419) );
  NAND2_X1 U574 ( .A1(n609), .A2(n424), .ZN(n423) );
  INV_X1 U575 ( .A(n468), .ZN(n424) );
  AND2_X1 U576 ( .A1(n628), .A2(n366), .ZN(n426) );
  INV_X1 U577 ( .A(n758), .ZN(n464) );
  NOR2_X2 U578 ( .A1(n717), .A2(n774), .ZN(n719) );
  NAND2_X1 U579 ( .A1(n462), .A2(n457), .ZN(n428) );
  XNOR2_X1 U580 ( .A(n708), .B(n467), .ZN(n450) );
  NAND2_X1 U581 ( .A1(n459), .A2(n764), .ZN(n429) );
  XNOR2_X1 U582 ( .A(n430), .B(n602), .ZN(n611) );
  NAND2_X1 U583 ( .A1(n365), .A2(n421), .ZN(n435) );
  NOR2_X1 U584 ( .A1(n744), .A2(n443), .ZN(n438) );
  NAND2_X1 U585 ( .A1(n744), .A2(n442), .ZN(n441) );
  XNOR2_X2 U586 ( .A(n621), .B(KEYINPUT31), .ZN(n760) );
  NAND2_X1 U587 ( .A1(n637), .A2(KEYINPUT34), .ZN(n455) );
  XNOR2_X2 U588 ( .A(n636), .B(n635), .ZN(n700) );
  XNOR2_X2 U589 ( .A(n456), .B(G143), .ZN(n542) );
  XNOR2_X2 U590 ( .A(G128), .B(KEYINPUT65), .ZN(n456) );
  INV_X1 U591 ( .A(n801), .ZN(n458) );
  AND2_X1 U592 ( .A1(n801), .A2(n574), .ZN(n460) );
  INV_X1 U593 ( .A(n574), .ZN(n461) );
  NAND2_X1 U594 ( .A1(n464), .A2(n463), .ZN(n585) );
  NAND2_X1 U595 ( .A1(n583), .A2(n582), .ZN(n465) );
  XNOR2_X1 U596 ( .A(n510), .B(n522), .ZN(n478) );
  XOR2_X1 U597 ( .A(n562), .B(n561), .Z(n468) );
  AND2_X1 U598 ( .A1(n679), .A2(n566), .ZN(n469) );
  INV_X1 U599 ( .A(KEYINPUT5), .ZN(n474) );
  AND2_X1 U600 ( .A1(n372), .A2(n469), .ZN(n567) );
  XNOR2_X1 U601 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U602 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U603 ( .A(n513), .B(n476), .ZN(n477) );
  XNOR2_X1 U604 ( .A(n558), .B(n726), .ZN(n559) );
  XNOR2_X1 U605 ( .A(n497), .B(n496), .ZN(n499) );
  INV_X1 U606 ( .A(KEYINPUT63), .ZN(n718) );
  XNOR2_X1 U607 ( .A(n772), .B(n771), .ZN(n773) );
  XNOR2_X1 U608 ( .A(n705), .B(n704), .ZN(G75) );
  XNOR2_X1 U609 ( .A(KEYINPUT69), .B(G101), .ZN(n471) );
  INV_X1 U610 ( .A(KEYINPUT3), .ZN(n472) );
  XNOR2_X1 U611 ( .A(n792), .B(n437), .ZN(n513) );
  NAND2_X1 U612 ( .A1(n548), .A2(G210), .ZN(n475) );
  INV_X1 U613 ( .A(KEYINPUT77), .ZN(n479) );
  XNOR2_X1 U614 ( .A(n479), .B(G472), .ZN(n480) );
  NAND2_X1 U615 ( .A1(n515), .A2(n481), .ZN(n529) );
  NAND2_X1 U616 ( .A1(n529), .A2(G214), .ZN(n668) );
  NAND2_X1 U617 ( .A1(n684), .A2(n668), .ZN(n482) );
  XNOR2_X1 U618 ( .A(n482), .B(KEYINPUT30), .ZN(n488) );
  NAND2_X1 U619 ( .A1(G234), .A2(G237), .ZN(n483) );
  XNOR2_X1 U620 ( .A(n483), .B(KEYINPUT14), .ZN(n696) );
  INV_X1 U621 ( .A(G952), .ZN(n716) );
  NAND2_X1 U622 ( .A1(n793), .A2(n716), .ZN(n485) );
  OR2_X1 U623 ( .A1(n793), .A2(G902), .ZN(n484) );
  AND2_X1 U624 ( .A1(n485), .A2(n484), .ZN(n486) );
  AND2_X1 U625 ( .A1(n696), .A2(n486), .ZN(n613) );
  NAND2_X1 U626 ( .A1(G953), .A2(G900), .ZN(n487) );
  NAND2_X1 U627 ( .A1(n613), .A2(n487), .ZN(n565) );
  XOR2_X1 U628 ( .A(KEYINPUT98), .B(KEYINPUT24), .Z(n490) );
  XNOR2_X1 U629 ( .A(n490), .B(n489), .ZN(n494) );
  NAND2_X1 U630 ( .A1(G234), .A2(n793), .ZN(n495) );
  NAND2_X1 U631 ( .A1(G221), .A2(n540), .ZN(n496) );
  NAND2_X1 U632 ( .A1(G234), .A2(n709), .ZN(n500) );
  XNOR2_X1 U633 ( .A(KEYINPUT20), .B(n500), .ZN(n504) );
  AND2_X1 U634 ( .A1(G217), .A2(n504), .ZN(n501) );
  XNOR2_X1 U635 ( .A(KEYINPUT25), .B(n501), .ZN(n502) );
  XNOR2_X2 U636 ( .A(n503), .B(n502), .ZN(n679) );
  AND2_X1 U637 ( .A1(n504), .A2(G221), .ZN(n506) );
  INV_X1 U638 ( .A(KEYINPUT21), .ZN(n505) );
  XNOR2_X1 U639 ( .A(n506), .B(n505), .ZN(n678) );
  INV_X1 U640 ( .A(G104), .ZN(n507) );
  XNOR2_X1 U641 ( .A(n508), .B(n507), .ZN(n782) );
  XNOR2_X1 U642 ( .A(n782), .B(KEYINPUT75), .ZN(n509) );
  NAND2_X1 U643 ( .A1(n793), .A2(G227), .ZN(n511) );
  XNOR2_X1 U644 ( .A(n511), .B(G140), .ZN(n512) );
  XNOR2_X1 U645 ( .A(n513), .B(n512), .ZN(n514) );
  NAND2_X1 U646 ( .A1(n732), .A2(n515), .ZN(n516) );
  XNOR2_X1 U647 ( .A(n622), .B(KEYINPUT109), .ZN(n517) );
  NAND2_X1 U648 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U649 ( .A(n519), .B(KEYINPUT80), .ZN(n595) );
  XOR2_X1 U650 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n524) );
  XNOR2_X1 U651 ( .A(n524), .B(n523), .ZN(n525) );
  NAND2_X1 U652 ( .A1(G224), .A2(n793), .ZN(n527) );
  INV_X1 U653 ( .A(n709), .ZN(n706) );
  NAND2_X1 U654 ( .A1(n529), .A2(G210), .ZN(n531) );
  XNOR2_X1 U655 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n530) );
  XNOR2_X1 U656 ( .A(n575), .B(KEYINPUT38), .ZN(n563) );
  NOR2_X1 U657 ( .A1(n595), .A2(n563), .ZN(n532) );
  XNOR2_X1 U658 ( .A(n532), .B(KEYINPUT39), .ZN(n609) );
  XNOR2_X1 U659 ( .A(n534), .B(n533), .ZN(n538) );
  XOR2_X1 U660 ( .A(n539), .B(KEYINPUT100), .Z(n545) );
  NAND2_X1 U661 ( .A1(n540), .A2(G217), .ZN(n541) );
  XNOR2_X1 U662 ( .A(n541), .B(G134), .ZN(n543) );
  XNOR2_X1 U663 ( .A(n545), .B(n544), .ZN(n767) );
  NAND2_X1 U664 ( .A1(G214), .A2(n548), .ZN(n549) );
  XNOR2_X1 U665 ( .A(n790), .B(n549), .ZN(n557) );
  XNOR2_X1 U666 ( .A(n550), .B(G143), .ZN(n551) );
  XNOR2_X1 U667 ( .A(n551), .B(G104), .ZN(n555) );
  XNOR2_X1 U668 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U669 ( .A(n555), .B(n554), .Z(n556) );
  XNOR2_X1 U670 ( .A(n557), .B(n556), .ZN(n727) );
  NOR2_X1 U671 ( .A1(G902), .A2(n727), .ZN(n560) );
  XNOR2_X1 U672 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n558) );
  INV_X1 U673 ( .A(G475), .ZN(n726) );
  INV_X1 U674 ( .A(n598), .ZN(n584) );
  XNOR2_X1 U675 ( .A(KEYINPUT113), .B(KEYINPUT40), .ZN(n562) );
  INV_X1 U676 ( .A(KEYINPUT112), .ZN(n561) );
  NAND2_X1 U677 ( .A1(n669), .A2(n668), .ZN(n672) );
  OR2_X1 U678 ( .A1(n599), .A2(n598), .ZN(n671) );
  XOR2_X1 U679 ( .A(KEYINPUT41), .B(n564), .Z(n677) );
  NOR2_X1 U680 ( .A1(n678), .A2(n565), .ZN(n566) );
  XNOR2_X1 U681 ( .A(n567), .B(KEYINPUT28), .ZN(n569) );
  NAND2_X1 U682 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U683 ( .A1(n677), .A2(n583), .ZN(n573) );
  XOR2_X1 U684 ( .A(KEYINPUT115), .B(KEYINPUT42), .Z(n571) );
  XNOR2_X1 U685 ( .A(n571), .B(KEYINPUT114), .ZN(n572) );
  XNOR2_X1 U686 ( .A(KEYINPUT91), .B(KEYINPUT46), .ZN(n574) );
  NOR2_X1 U687 ( .A1(n576), .A2(n379), .ZN(n579) );
  INV_X1 U688 ( .A(KEYINPUT93), .ZN(n577) );
  XNOR2_X1 U689 ( .A(n577), .B(KEYINPUT36), .ZN(n578) );
  XNOR2_X1 U690 ( .A(n579), .B(n578), .ZN(n580) );
  BUF_X1 U691 ( .A(n615), .Z(n582) );
  NAND2_X1 U692 ( .A1(n599), .A2(n584), .ZN(n751) );
  NOR2_X1 U693 ( .A1(KEYINPUT83), .A2(n624), .ZN(n587) );
  NAND2_X1 U694 ( .A1(KEYINPUT47), .A2(n673), .ZN(n586) );
  AND2_X1 U695 ( .A1(n586), .A2(KEYINPUT83), .ZN(n589) );
  NOR2_X1 U696 ( .A1(n758), .A2(n588), .ZN(n593) );
  INV_X1 U697 ( .A(n589), .ZN(n591) );
  INV_X1 U698 ( .A(KEYINPUT47), .ZN(n590) );
  AND2_X1 U699 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U700 ( .A1(n593), .A2(n592), .ZN(n594) );
  INV_X1 U701 ( .A(n575), .ZN(n607) );
  INV_X1 U702 ( .A(KEYINPUT110), .ZN(n596) );
  XNOR2_X1 U703 ( .A(n597), .B(n596), .ZN(n601) );
  NAND2_X1 U704 ( .A1(n599), .A2(n598), .ZN(n638) );
  INV_X1 U705 ( .A(n638), .ZN(n600) );
  INV_X1 U706 ( .A(KEYINPUT48), .ZN(n602) );
  AND2_X1 U707 ( .A1(n603), .A2(n668), .ZN(n605) );
  INV_X1 U708 ( .A(n681), .ZN(n604) );
  NAND2_X1 U709 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U710 ( .A(n606), .B(KEYINPUT43), .ZN(n608) );
  NAND2_X1 U711 ( .A1(n608), .A2(n607), .ZN(n721) );
  OR2_X1 U712 ( .A1(n609), .A2(n751), .ZN(n722) );
  AND2_X1 U713 ( .A1(n721), .A2(n722), .ZN(n610) );
  NAND2_X1 U714 ( .A1(G953), .A2(G898), .ZN(n612) );
  AND2_X1 U715 ( .A1(n613), .A2(n612), .ZN(n614) );
  INV_X1 U716 ( .A(KEYINPUT68), .ZN(n616) );
  XNOR2_X1 U717 ( .A(n616), .B(KEYINPUT0), .ZN(n617) );
  AND2_X1 U718 ( .A1(n372), .A2(n358), .ZN(n620) );
  AND2_X1 U719 ( .A1(n681), .A2(n620), .ZN(n688) );
  NOR2_X1 U720 ( .A1(n372), .A2(n622), .ZN(n623) );
  NOR2_X1 U721 ( .A1(n671), .A2(n678), .ZN(n625) );
  XNOR2_X1 U722 ( .A(n625), .B(KEYINPUT106), .ZN(n626) );
  OR2_X1 U723 ( .A1(n681), .A2(n679), .ZN(n630) );
  INV_X1 U724 ( .A(n741), .ZN(n631) );
  INV_X1 U725 ( .A(n633), .ZN(n637) );
  NAND2_X1 U726 ( .A1(n634), .A2(n681), .ZN(n636) );
  XOR2_X1 U727 ( .A(KEYINPUT33), .B(KEYINPUT76), .Z(n635) );
  XNOR2_X1 U728 ( .A(n638), .B(KEYINPUT81), .ZN(n639) );
  INV_X1 U729 ( .A(KEYINPUT35), .ZN(n640) );
  INV_X1 U730 ( .A(KEYINPUT44), .ZN(n650) );
  XNOR2_X1 U731 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n642) );
  XNOR2_X2 U732 ( .A(n643), .B(n642), .ZN(n725) );
  INV_X1 U733 ( .A(n679), .ZN(n644) );
  OR2_X1 U734 ( .A1(n372), .A2(n644), .ZN(n645) );
  OR2_X1 U735 ( .A1(n645), .A2(n681), .ZN(n646) );
  AND2_X1 U736 ( .A1(n650), .A2(KEYINPUT92), .ZN(n648) );
  INV_X1 U737 ( .A(KEYINPUT92), .ZN(n649) );
  XNOR2_X1 U738 ( .A(KEYINPUT90), .B(KEYINPUT45), .ZN(n652) );
  XNOR2_X1 U739 ( .A(n652), .B(KEYINPUT64), .ZN(n653) );
  NOR2_X1 U740 ( .A1(n654), .A2(KEYINPUT2), .ZN(n656) );
  INV_X1 U741 ( .A(KEYINPUT84), .ZN(n655) );
  NOR2_X1 U742 ( .A1(KEYINPUT2), .A2(KEYINPUT84), .ZN(n657) );
  NAND2_X1 U743 ( .A1(n775), .A2(n657), .ZN(n658) );
  NOR2_X1 U744 ( .A1(n660), .A2(n659), .ZN(n665) );
  INV_X1 U745 ( .A(KEYINPUT2), .ZN(n661) );
  NOR2_X1 U746 ( .A1(n359), .A2(n661), .ZN(n663) );
  NAND2_X1 U747 ( .A1(n775), .A2(n663), .ZN(n712) );
  INV_X1 U748 ( .A(n712), .ZN(n664) );
  XNOR2_X1 U749 ( .A(n666), .B(KEYINPUT87), .ZN(n667) );
  NOR2_X1 U750 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U751 ( .A1(n671), .A2(n670), .ZN(n675) );
  NOR2_X1 U752 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U753 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U754 ( .A1(n356), .A2(n676), .ZN(n694) );
  INV_X1 U755 ( .A(n677), .ZN(n699) );
  NAND2_X1 U756 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U757 ( .A(KEYINPUT49), .B(n680), .Z(n687) );
  NOR2_X1 U758 ( .A1(n681), .A2(n358), .ZN(n683) );
  XNOR2_X1 U759 ( .A(KEYINPUT122), .B(KEYINPUT50), .ZN(n682) );
  XNOR2_X1 U760 ( .A(n683), .B(n682), .ZN(n685) );
  NOR2_X1 U761 ( .A1(n685), .A2(n372), .ZN(n686) );
  NAND2_X1 U762 ( .A1(n687), .A2(n686), .ZN(n690) );
  INV_X1 U763 ( .A(n688), .ZN(n689) );
  NAND2_X1 U764 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U765 ( .A(n691), .B(KEYINPUT51), .ZN(n692) );
  NOR2_X1 U766 ( .A1(n699), .A2(n692), .ZN(n693) );
  NOR2_X1 U767 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U768 ( .A(KEYINPUT52), .B(n695), .ZN(n698) );
  NAND2_X1 U769 ( .A1(n696), .A2(G952), .ZN(n697) );
  NOR2_X1 U770 ( .A1(n698), .A2(n697), .ZN(n702) );
  NOR2_X1 U771 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U772 ( .A(KEYINPUT123), .B(KEYINPUT53), .ZN(n704) );
  NAND2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U774 ( .A(n709), .B(KEYINPUT88), .Z(n710) );
  NAND2_X1 U775 ( .A1(n710), .A2(KEYINPUT2), .ZN(n711) );
  NAND2_X1 U776 ( .A1(n769), .A2(G472), .ZN(n715) );
  XOR2_X1 U777 ( .A(KEYINPUT62), .B(n713), .Z(n714) );
  XNOR2_X1 U778 ( .A(n715), .B(n714), .ZN(n717) );
  XNOR2_X1 U779 ( .A(n719), .B(n718), .ZN(G57) );
  INV_X1 U780 ( .A(n751), .ZN(n743) );
  NAND2_X1 U781 ( .A1(n394), .A2(n743), .ZN(n720) );
  XNOR2_X1 U782 ( .A(n720), .B(G116), .ZN(G18) );
  XNOR2_X1 U783 ( .A(n721), .B(G140), .ZN(G42) );
  XNOR2_X1 U784 ( .A(n722), .B(G134), .ZN(G36) );
  XNOR2_X1 U785 ( .A(n723), .B(G131), .ZN(G33) );
  XOR2_X1 U786 ( .A(G119), .B(KEYINPUT127), .Z(n724) );
  XNOR2_X1 U787 ( .A(n725), .B(n724), .ZN(G21) );
  XNOR2_X1 U788 ( .A(n727), .B(KEYINPUT59), .ZN(n728) );
  XNOR2_X1 U789 ( .A(n363), .B(n728), .ZN(n729) );
  NOR2_X1 U790 ( .A1(n729), .A2(n774), .ZN(n730) );
  XNOR2_X1 U791 ( .A(n730), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U792 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n731) );
  XNOR2_X1 U793 ( .A(n732), .B(n731), .ZN(n733) );
  XNOR2_X1 U794 ( .A(n362), .B(n733), .ZN(n734) );
  NOR2_X1 U795 ( .A1(n734), .A2(n774), .ZN(G54) );
  NAND2_X1 U796 ( .A1(n769), .A2(G210), .ZN(n738) );
  XOR2_X1 U797 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n736) );
  XNOR2_X1 U798 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U799 ( .A(n740), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U800 ( .A(n741), .B(G101), .Z(G3) );
  NAND2_X1 U801 ( .A1(n744), .A2(n421), .ZN(n742) );
  XNOR2_X1 U802 ( .A(n742), .B(G104), .ZN(G6) );
  XOR2_X1 U803 ( .A(KEYINPUT27), .B(KEYINPUT117), .Z(n746) );
  NAND2_X1 U804 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U805 ( .A(n746), .B(n745), .ZN(n748) );
  XOR2_X1 U806 ( .A(G107), .B(KEYINPUT26), .Z(n747) );
  XNOR2_X1 U807 ( .A(n748), .B(n747), .ZN(G9) );
  INV_X1 U808 ( .A(n749), .ZN(n750) );
  XOR2_X1 U809 ( .A(G110), .B(n750), .Z(G12) );
  NOR2_X1 U810 ( .A1(n399), .A2(n751), .ZN(n753) );
  XNOR2_X1 U811 ( .A(KEYINPUT118), .B(KEYINPUT29), .ZN(n752) );
  XNOR2_X1 U812 ( .A(n753), .B(n752), .ZN(n754) );
  XNOR2_X1 U813 ( .A(G128), .B(n754), .ZN(G30) );
  XNOR2_X1 U814 ( .A(G143), .B(n755), .ZN(n756) );
  XNOR2_X1 U815 ( .A(n756), .B(KEYINPUT119), .ZN(G45) );
  NOR2_X1 U816 ( .A1(n399), .A2(n757), .ZN(n759) );
  XOR2_X1 U817 ( .A(G146), .B(n759), .Z(G48) );
  NAND2_X1 U818 ( .A1(n394), .A2(n421), .ZN(n761) );
  XNOR2_X1 U819 ( .A(n761), .B(KEYINPUT120), .ZN(n762) );
  XNOR2_X1 U820 ( .A(G113), .B(n762), .ZN(G15) );
  XNOR2_X1 U821 ( .A(KEYINPUT37), .B(KEYINPUT121), .ZN(n763) );
  XNOR2_X1 U822 ( .A(n764), .B(n763), .ZN(n765) );
  XNOR2_X1 U823 ( .A(G125), .B(n765), .ZN(G27) );
  NAND2_X1 U824 ( .A1(n378), .A2(G478), .ZN(n766) );
  XNOR2_X1 U825 ( .A(n767), .B(n766), .ZN(n768) );
  NOR2_X1 U826 ( .A1(n774), .A2(n768), .ZN(G63) );
  NAND2_X1 U827 ( .A1(n378), .A2(G217), .ZN(n772) );
  NOR2_X1 U828 ( .A1(n774), .A2(n773), .ZN(G66) );
  NAND2_X1 U829 ( .A1(n775), .A2(n793), .ZN(n780) );
  XOR2_X1 U830 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n777) );
  NAND2_X1 U831 ( .A1(G224), .A2(G953), .ZN(n776) );
  XNOR2_X1 U832 ( .A(n777), .B(n776), .ZN(n778) );
  NAND2_X1 U833 ( .A1(n778), .A2(G898), .ZN(n779) );
  NAND2_X1 U834 ( .A1(n780), .A2(n779), .ZN(n788) );
  XNOR2_X1 U835 ( .A(n781), .B(G101), .ZN(n783) );
  XNOR2_X1 U836 ( .A(n783), .B(n782), .ZN(n785) );
  NOR2_X1 U837 ( .A1(G898), .A2(n793), .ZN(n784) );
  NOR2_X1 U838 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U839 ( .A(KEYINPUT126), .B(n786), .ZN(n787) );
  XNOR2_X1 U840 ( .A(n788), .B(n787), .ZN(G69) );
  XNOR2_X1 U841 ( .A(n789), .B(n790), .ZN(n791) );
  XNOR2_X1 U842 ( .A(n792), .B(n791), .ZN(n795) );
  NAND2_X1 U843 ( .A1(n794), .A2(n793), .ZN(n799) );
  XNOR2_X1 U844 ( .A(G227), .B(n795), .ZN(n796) );
  NAND2_X1 U845 ( .A1(n796), .A2(G900), .ZN(n797) );
  NAND2_X1 U846 ( .A1(n797), .A2(G953), .ZN(n798) );
  NAND2_X1 U847 ( .A1(n799), .A2(n798), .ZN(G72) );
  XNOR2_X1 U848 ( .A(n800), .B(G122), .ZN(G24) );
  XNOR2_X1 U849 ( .A(G137), .B(n801), .ZN(G39) );
endmodule

