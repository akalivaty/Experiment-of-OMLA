//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G224), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n190), .B(KEYINPUT93), .Z(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT65), .B1(new_n192), .B2(G146), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n199));
  AND4_X1   g013(.A1(new_n193), .A2(new_n196), .A3(new_n197), .A4(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT70), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n195), .A2(G143), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n198), .B1(new_n202), .B2(KEYINPUT1), .ZN(new_n203));
  XNOR2_X1  g017(.A(G143), .B(G146), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n201), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G128), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n202), .A2(new_n197), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(KEYINPUT70), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n200), .B1(new_n205), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G125), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT94), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n208), .B1(KEYINPUT0), .B2(G128), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT0), .A2(G128), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n215), .B(KEYINPUT64), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n193), .A2(new_n196), .A3(new_n197), .ZN(new_n217));
  OAI22_X1  g031(.A1(new_n214), .A2(new_n216), .B1(new_n217), .B2(new_n215), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G125), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n212), .A2(new_n213), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n213), .B1(new_n212), .B2(new_n219), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n191), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n222), .ZN(new_n224));
  INV_X1    g038(.A(new_n191), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n225), .A3(new_n220), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT92), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT5), .ZN(new_n230));
  INV_X1    g044(.A(G119), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n231), .A3(G116), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(G116), .ZN(new_n233));
  INV_X1    g047(.A(G116), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G119), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(G113), .B(new_n232), .C1(new_n236), .C2(new_n230), .ZN(new_n237));
  INV_X1    g051(.A(G113), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT2), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT2), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G113), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(new_n233), .A3(new_n235), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n237), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G104), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT3), .B1(new_n245), .B2(G107), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT3), .ZN(new_n247));
  INV_X1    g061(.A(G107), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(G104), .ZN(new_n249));
  INV_X1    g063(.A(G101), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n245), .A2(G107), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n246), .A2(new_n249), .A3(new_n250), .A4(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n245), .A2(G107), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n248), .A2(G104), .ZN(new_n254));
  OAI21_X1  g068(.A(G101), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n244), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n246), .A2(new_n249), .A3(new_n251), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G101), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT4), .A3(new_n252), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n258), .A2(new_n261), .A3(G101), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT2), .B(G113), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n236), .B1(new_n264), .B2(KEYINPUT71), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n239), .A2(new_n241), .A3(KEYINPUT71), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT72), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n240), .A2(G113), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n238), .A2(KEYINPUT2), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n272), .A2(new_n273), .A3(new_n266), .A4(new_n236), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n268), .A2(new_n243), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n257), .B1(new_n263), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(G110), .B(G122), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n229), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n274), .A2(new_n243), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n242), .A2(new_n269), .B1(new_n233), .B2(new_n235), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n273), .B1(new_n280), .B2(new_n266), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n262), .B(new_n260), .C1(new_n279), .C2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n256), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(new_n243), .A3(new_n237), .ZN(new_n284));
  AND4_X1   g098(.A1(new_n229), .A2(new_n282), .A3(new_n284), .A4(new_n277), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT6), .B1(new_n278), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT91), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n282), .B2(new_n284), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n276), .A2(new_n287), .ZN(new_n290));
  INV_X1    g104(.A(new_n277), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n289), .A2(new_n290), .A3(KEYINPUT6), .A4(new_n291), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n228), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT7), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n191), .A2(new_n296), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n212), .A2(new_n219), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n297), .B1(new_n212), .B2(new_n219), .ZN(new_n299));
  XOR2_X1   g113(.A(new_n277), .B(KEYINPUT8), .Z(new_n300));
  NAND2_X1  g114(.A1(new_n244), .A2(new_n256), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n300), .B1(new_n284), .B2(new_n301), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n298), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n303), .B1(new_n278), .B2(new_n285), .ZN(new_n304));
  INV_X1    g118(.A(G902), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n188), .B1(new_n295), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT6), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n282), .A2(new_n284), .A3(new_n277), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT92), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n276), .A2(new_n229), .A3(new_n277), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI211_X1 g126(.A(KEYINPUT91), .B(new_n257), .C1(new_n263), .C2(new_n275), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n313), .A2(new_n288), .A3(new_n277), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n294), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n227), .ZN(new_n316));
  INV_X1    g130(.A(new_n306), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(new_n187), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n307), .A2(new_n318), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n189), .A2(G952), .ZN(new_n320));
  INV_X1    g134(.A(G234), .ZN(new_n321));
  INV_X1    g135(.A(G237), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  XOR2_X1   g138(.A(KEYINPUT78), .B(G902), .Z(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  AOI211_X1 g140(.A(new_n189), .B(new_n326), .C1(G234), .C2(G237), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT21), .B(G898), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(G214), .B1(G237), .B2(G902), .ZN(new_n331));
  NOR2_X1   g145(.A1(G475), .A2(G902), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(KEYINPUT97), .ZN(new_n333));
  XNOR2_X1  g147(.A(G113), .B(G122), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(new_n245), .ZN(new_n335));
  XNOR2_X1  g149(.A(G125), .B(G140), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT19), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT85), .B1(KEYINPUT84), .B2(G125), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n340), .A2(G140), .ZN(new_n341));
  AND2_X1   g155(.A1(KEYINPUT85), .A2(G125), .ZN(new_n342));
  OAI21_X1  g156(.A(G140), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n195), .B(new_n339), .C1(new_n344), .C2(new_n337), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT96), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT16), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(new_n341), .B2(new_n343), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n347), .B1(new_n211), .B2(G140), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(G146), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  AND2_X1   g165(.A1(KEYINPUT66), .A2(G131), .ZN(new_n352));
  NOR2_X1   g166(.A1(KEYINPUT66), .A2(G131), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(G237), .A2(G953), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(G143), .A3(G214), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(G143), .B1(new_n356), .B2(G214), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n355), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n322), .A2(new_n189), .A3(G214), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n192), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n354), .A3(new_n357), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n341), .A2(new_n343), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n338), .B1(new_n365), .B2(KEYINPUT19), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT96), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(new_n195), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n346), .A2(new_n351), .A3(new_n364), .A4(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n362), .A2(KEYINPUT95), .A3(new_n357), .ZN(new_n370));
  NAND2_X1  g184(.A1(KEYINPUT18), .A2(G131), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n336), .A2(new_n195), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n344), .B2(new_n195), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n335), .B1(new_n369), .B2(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n195), .B(new_n349), .C1(new_n344), .C2(new_n347), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n351), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n355), .B(KEYINPUT17), .C1(new_n358), .C2(new_n359), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n379), .B1(new_n364), .B2(KEYINPUT17), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n375), .B(new_n335), .C1(new_n378), .C2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n333), .B1(new_n376), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT20), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT20), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n385), .B(new_n333), .C1(new_n376), .C2(new_n382), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G475), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n375), .B1(new_n378), .B2(new_n380), .ZN(new_n389));
  INV_X1    g203(.A(new_n335), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n381), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n388), .B1(new_n392), .B2(new_n305), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n192), .A2(G128), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n198), .A2(G143), .ZN(new_n396));
  INV_X1    g210(.A(G134), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G116), .B(G122), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G107), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n248), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n398), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT13), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n395), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n396), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n395), .A2(new_n404), .ZN(new_n407));
  OAI21_X1  g221(.A(G134), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n234), .A2(KEYINPUT14), .A3(G122), .ZN(new_n410));
  OAI211_X1 g224(.A(G107), .B(new_n410), .C1(new_n400), .C2(KEYINPUT14), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n397), .B1(new_n395), .B2(new_n396), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n411), .B(new_n402), .C1(new_n398), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT9), .B(G234), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(G217), .A3(new_n189), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n417), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n409), .A2(new_n413), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(KEYINPUT98), .A3(new_n326), .ZN(new_n422));
  INV_X1    g236(.A(G478), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(KEYINPUT15), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n424), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n421), .A2(KEYINPUT98), .A3(new_n326), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n387), .A2(new_n394), .A3(new_n429), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n319), .A2(new_n330), .A3(new_n331), .A4(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(G110), .B(G140), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(KEYINPUT87), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n189), .A2(G227), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT0), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n204), .B1(new_n436), .B2(new_n198), .ZN(new_n437));
  INV_X1    g251(.A(new_n216), .ZN(new_n438));
  INV_X1    g252(.A(new_n217), .ZN(new_n439));
  INV_X1    g253(.A(new_n215), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n437), .A2(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT10), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n217), .A2(new_n207), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n193), .A2(new_n196), .A3(new_n197), .A4(new_n199), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n283), .A2(new_n445), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n263), .A2(new_n441), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n203), .A2(new_n204), .A3(new_n201), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT70), .B1(new_n207), .B2(new_n208), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n444), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT88), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n252), .A2(new_n255), .A3(KEYINPUT10), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT88), .B1(new_n210), .B2(new_n452), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT11), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n397), .B2(G137), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n397), .A2(G137), .ZN(new_n459));
  INV_X1    g273(.A(G137), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(KEYINPUT11), .A3(G134), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G131), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n354), .A2(new_n459), .A3(new_n458), .A4(new_n461), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT73), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT73), .B1(new_n463), .B2(new_n464), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n447), .A2(new_n456), .A3(new_n467), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n444), .B(new_n256), .C1(new_n448), .C2(new_n449), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n446), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n463), .A2(new_n464), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n471), .A2(KEYINPUT12), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT73), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT73), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n446), .A2(new_n469), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n473), .B1(new_n477), .B2(KEYINPUT12), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n435), .B1(new_n468), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n454), .A2(new_n455), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n446), .A2(new_n442), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n260), .A2(new_n262), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n482), .B1(new_n218), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n480), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n467), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n447), .A2(new_n456), .A3(KEYINPUT89), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n468), .A2(new_n435), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n479), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G469), .B1(new_n490), .B2(G902), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT90), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(KEYINPUT90), .B(G469), .C1(new_n490), .C2(G902), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n489), .A2(new_n478), .ZN(new_n495));
  INV_X1    g309(.A(new_n468), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n447), .A2(new_n456), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n467), .B1(new_n497), .B2(new_n480), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n496), .B1(new_n498), .B2(new_n487), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n495), .B1(new_n499), .B2(new_n435), .ZN(new_n500));
  INV_X1    g314(.A(G469), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n501), .A3(new_n326), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n493), .A2(new_n494), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G221), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(new_n416), .B2(new_n305), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n431), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT77), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT75), .B1(new_n279), .B2(new_n281), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT75), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n268), .A2(new_n511), .A3(new_n243), .A4(new_n274), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT68), .B1(new_n397), .B2(G137), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT68), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(new_n460), .A3(G134), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(new_n516), .A3(new_n459), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G131), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(KEYINPUT69), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT69), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n520), .B1(new_n517), .B2(G131), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n450), .B(new_n464), .C1(new_n519), .C2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n441), .B1(new_n465), .B2(new_n466), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT74), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(KEYINPUT74), .B(new_n441), .C1(new_n465), .C2(new_n466), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n513), .A2(new_n522), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n522), .A3(new_n526), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n527), .B1(new_n529), .B2(new_n513), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT28), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n522), .A2(new_n523), .A3(new_n510), .A4(new_n512), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT28), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n356), .A2(G210), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(KEYINPUT27), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT26), .B(G101), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT29), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n509), .B1(new_n535), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n534), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n441), .A2(new_n471), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT67), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT67), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n441), .A2(new_n548), .A3(new_n471), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(new_n522), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n275), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n527), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n545), .B1(new_n552), .B2(KEYINPUT28), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n539), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT30), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n525), .A2(KEYINPUT30), .A3(new_n522), .A4(new_n526), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(new_n275), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n527), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n540), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n554), .A2(new_n541), .A3(new_n560), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n531), .A2(KEYINPUT77), .A3(new_n534), .A4(new_n542), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n544), .A2(new_n561), .A3(new_n326), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(G472), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n553), .A2(new_n539), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT76), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n525), .A2(new_n526), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n522), .A2(new_n510), .A3(new_n512), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n566), .B(new_n539), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n566), .B1(new_n527), .B2(new_n539), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n558), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT31), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(KEYINPUT31), .B(new_n558), .C1(new_n570), .C2(new_n571), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n565), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(G472), .A2(G902), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n576), .A2(KEYINPUT32), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT32), .ZN(new_n580));
  OR2_X1    g394(.A1(new_n553), .A2(new_n539), .ZN(new_n581));
  INV_X1    g395(.A(new_n575), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n539), .B1(new_n567), .B2(new_n568), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT76), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n569), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT31), .B1(new_n585), .B2(new_n558), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n581), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n580), .B1(new_n587), .B2(new_n577), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n564), .B1(new_n579), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT25), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT24), .B(G110), .ZN(new_n591));
  OR2_X1    g405(.A1(new_n591), .A2(KEYINPUT80), .ZN(new_n592));
  XNOR2_X1  g406(.A(G119), .B(G128), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(KEYINPUT80), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT81), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT80), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n591), .B(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT81), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n599), .A3(new_n593), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n601));
  XOR2_X1   g415(.A(new_n601), .B(KEYINPUT82), .Z(new_n602));
  NOR2_X1   g416(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(G119), .B2(new_n198), .ZN(new_n604));
  NAND2_X1  g418(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n604), .A2(new_n605), .B1(new_n231), .B2(G128), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n596), .A2(new_n600), .B1(G110), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n378), .ZN(new_n609));
  OAI22_X1  g423(.A1(new_n607), .A2(G110), .B1(new_n598), .B2(new_n593), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(new_n351), .A3(new_n373), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT22), .B(G137), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n504), .A2(new_n321), .A3(G953), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n609), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n615), .B1(new_n609), .B2(new_n611), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n590), .B1(new_n619), .B2(new_n326), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n609), .A2(new_n611), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n614), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n622), .A2(new_n590), .A3(new_n326), .A4(new_n616), .ZN(new_n623));
  OAI21_X1  g437(.A(G217), .B1(new_n325), .B2(new_n321), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT79), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n620), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n625), .A2(new_n305), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n629), .B(KEYINPUT86), .Z(new_n630));
  AND2_X1   g444(.A1(new_n619), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n508), .A2(new_n589), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G101), .ZN(G3));
  OAI21_X1  g448(.A(KEYINPUT99), .B1(new_n576), .B2(new_n325), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT99), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n587), .A2(new_n636), .A3(new_n326), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(new_n637), .A3(G472), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n587), .A2(new_n577), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n503), .A2(new_n632), .A3(new_n506), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  AOI211_X1 g457(.A(new_n188), .B(new_n306), .C1(new_n227), .C2(new_n315), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n187), .B1(new_n316), .B2(new_n317), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n330), .B(new_n331), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n367), .B1(new_n366), .B2(new_n195), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n351), .A2(new_n364), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n649), .A2(new_n368), .B1(new_n374), .B2(new_n372), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n381), .B1(new_n650), .B2(new_n335), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n385), .B1(new_n651), .B2(new_n333), .ZN(new_n652));
  INV_X1    g466(.A(new_n386), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n394), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n421), .B(KEYINPUT33), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n325), .A2(new_n423), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n421), .A2(new_n326), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n423), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n643), .A2(new_n646), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT34), .B(G104), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G6));
  INV_X1    g478(.A(KEYINPUT100), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n387), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n384), .A2(KEYINPUT100), .A3(new_n386), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n429), .A2(new_n393), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n643), .A2(new_n646), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT35), .B(G107), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  NOR2_X1   g487(.A1(new_n614), .A2(KEYINPUT36), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n621), .B(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT101), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n675), .A2(new_n676), .A3(new_n630), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n621), .B1(KEYINPUT36), .B2(new_n614), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n609), .A2(new_n611), .A3(new_n674), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n630), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT101), .ZN(new_n681));
  OAI211_X1 g495(.A(new_n677), .B(new_n681), .C1(new_n620), .C2(new_n627), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n638), .A2(new_n639), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT102), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT102), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n638), .A2(new_n685), .A3(new_n639), .A4(new_n682), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n684), .A2(new_n508), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT37), .B(G110), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G12));
  INV_X1    g503(.A(new_n331), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n690), .B1(new_n307), .B2(new_n318), .ZN(new_n691));
  AND4_X1   g505(.A1(new_n506), .A2(new_n691), .A3(new_n503), .A4(new_n682), .ZN(new_n692));
  INV_X1    g506(.A(G900), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n324), .B1(new_n327), .B2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n669), .A2(new_n666), .A3(new_n667), .A4(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n589), .A2(new_n692), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G128), .ZN(G30));
  XOR2_X1   g513(.A(new_n694), .B(KEYINPUT39), .Z(new_n700));
  NAND3_X1  g514(.A1(new_n503), .A2(new_n506), .A3(new_n700), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n701), .A2(KEYINPUT40), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(KEYINPUT40), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n307), .A2(KEYINPUT38), .A3(new_n318), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT38), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n319), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n393), .B1(new_n384), .B2(new_n386), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n429), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n682), .A2(new_n690), .ZN(new_n709));
  AND4_X1   g523(.A1(new_n704), .A2(new_n706), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  AOI22_X1  g524(.A1(new_n585), .A2(new_n558), .B1(new_n540), .B2(new_n530), .ZN(new_n711));
  OAI21_X1  g525(.A(G472), .B1(new_n711), .B2(G902), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n712), .B1(new_n579), .B2(new_n588), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n702), .A2(new_n703), .A3(new_n710), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G143), .ZN(G45));
  NOR2_X1   g529(.A1(new_n661), .A2(new_n694), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n589), .A2(new_n692), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  INV_X1    g532(.A(new_n632), .ZN(new_n719));
  OAI21_X1  g533(.A(KEYINPUT32), .B1(new_n576), .B2(new_n578), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n587), .A2(new_n580), .A3(new_n577), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n719), .B1(new_n722), .B2(new_n564), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n435), .B1(new_n488), .B2(new_n468), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n489), .A2(new_n478), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n326), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n501), .A2(KEYINPUT103), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n727), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n326), .B(new_n729), .C1(new_n724), .C2(new_n725), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n728), .A2(new_n506), .A3(new_n730), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n646), .A2(new_n731), .A3(new_n661), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n723), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT41), .B(G113), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G15));
  NOR3_X1   g549(.A1(new_n670), .A2(new_n646), .A3(new_n731), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n723), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G116), .ZN(G18));
  AOI22_X1  g552(.A1(new_n720), .A2(new_n721), .B1(G472), .B2(new_n563), .ZN(new_n739));
  INV_X1    g553(.A(new_n731), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n430), .A2(new_n682), .A3(new_n330), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n742), .A3(new_n691), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT104), .B1(new_n739), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n319), .A2(new_n331), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n745), .A2(new_n731), .A3(new_n741), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT104), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n589), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G119), .ZN(G21));
  NAND4_X1  g564(.A1(new_n728), .A2(new_n708), .A3(new_n506), .A4(new_n730), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n646), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n535), .A2(new_n540), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n753), .B1(new_n582), .B2(new_n586), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n577), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n574), .A2(new_n575), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n325), .B1(new_n756), .B2(new_n581), .ZN(new_n757));
  INV_X1    g571(.A(G472), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n755), .B(new_n632), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT105), .B1(new_n752), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n587), .A2(new_n326), .ZN(new_n761));
  AOI22_X1  g575(.A1(new_n761), .A2(G472), .B1(new_n577), .B2(new_n754), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n646), .A2(new_n751), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT105), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n632), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G122), .ZN(G24));
  OAI211_X1 g581(.A(new_n755), .B(new_n682), .C1(new_n757), .C2(new_n758), .ZN(new_n768));
  INV_X1    g582(.A(new_n730), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n729), .B1(new_n500), .B2(new_n326), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n691), .A2(new_n771), .A3(new_n716), .A4(new_n506), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(new_n211), .ZN(G27));
  INV_X1    g588(.A(KEYINPUT106), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(new_n739), .B2(new_n719), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n589), .A2(KEYINPUT106), .A3(new_n632), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n319), .A2(new_n690), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n505), .B1(new_n502), .B2(new_n491), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT42), .ZN(new_n781));
  INV_X1    g595(.A(new_n716), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n776), .A2(new_n777), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT107), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n776), .A2(new_n777), .A3(KEYINPUT107), .A4(new_n783), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n780), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n723), .A2(new_n716), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n781), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G131), .ZN(G33));
  XOR2_X1   g607(.A(new_n696), .B(KEYINPUT108), .Z(new_n794));
  NAND3_X1  g608(.A1(new_n723), .A2(new_n789), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G134), .ZN(G36));
  NAND2_X1  g610(.A1(new_n707), .A2(new_n660), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT43), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n682), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n800), .B1(new_n639), .B2(new_n638), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n778), .B1(new_n801), .B2(KEYINPUT44), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT44), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n640), .A2(new_n803), .A3(new_n800), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT110), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n502), .ZN(new_n806));
  NAND2_X1  g620(.A1(G469), .A2(G902), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n490), .A2(KEYINPUT45), .ZN(new_n808));
  OAI21_X1  g622(.A(G469), .B1(new_n490), .B2(KEYINPUT45), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT46), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n806), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n812), .B1(new_n811), .B2(new_n810), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n506), .A3(new_n700), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT109), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n803), .B1(new_n640), .B2(new_n800), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n801), .A2(KEYINPUT44), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT110), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n778), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n805), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  XOR2_X1   g634(.A(KEYINPUT111), .B(G137), .Z(new_n821));
  XNOR2_X1  g635(.A(new_n820), .B(new_n821), .ZN(G39));
  XNOR2_X1  g636(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n813), .A2(new_n506), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n823), .B1(new_n813), .B2(new_n506), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n782), .A2(new_n632), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n739), .A3(new_n778), .A4(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(KEYINPUT113), .B(G140), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n828), .B(new_n829), .ZN(G42));
  OAI21_X1  g644(.A(KEYINPUT116), .B1(new_n654), .B2(new_n429), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n707), .A2(new_n832), .A3(new_n428), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT115), .B1(new_n654), .B2(new_n660), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n655), .A2(new_n656), .B1(new_n658), .B2(new_n423), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n707), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n646), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(new_n639), .A3(new_n638), .A4(new_n641), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n633), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n687), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n723), .B1(new_n732), .B2(new_n736), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n749), .A2(new_n766), .A3(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n682), .A2(new_n394), .A3(new_n429), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n668), .A2(new_n778), .A3(new_n695), .A4(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(new_n589), .A3(new_n506), .A4(new_n503), .ZN(new_n848));
  INV_X1    g662(.A(new_n768), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n849), .A2(new_n789), .A3(new_n716), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n795), .A3(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n843), .A2(new_n845), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n745), .A2(new_n731), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(new_n762), .A3(new_n682), .A4(new_n716), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n682), .A2(new_n694), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n691), .A2(new_n779), .A3(new_n855), .A4(new_n708), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n713), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n698), .A2(new_n717), .A3(new_n854), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n858), .B(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n852), .A2(new_n792), .A3(new_n860), .A4(KEYINPUT53), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n691), .A2(new_n503), .A3(new_n506), .A4(new_n682), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n739), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n773), .B1(new_n863), .B2(new_n697), .ZN(new_n864));
  AND2_X1   g678(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n865));
  NOR2_X1   g679(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n864), .A2(new_n717), .A3(new_n857), .A4(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n858), .A2(new_n865), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n852), .A2(new_n792), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n861), .B1(new_n871), .B2(KEYINPUT53), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT54), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n852), .A2(new_n792), .A3(new_n860), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n852), .A2(new_n792), .A3(new_n870), .A4(KEYINPUT53), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n759), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n799), .A2(new_n324), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n883), .A2(new_n690), .A3(new_n319), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n826), .A2(KEYINPUT118), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n771), .A2(new_n505), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n826), .A2(KEYINPUT118), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n713), .ZN(new_n890));
  NOR4_X1   g704(.A1(new_n731), .A2(new_n319), .A3(new_n323), .A4(new_n690), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n632), .A3(new_n891), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n892), .A2(new_n654), .A3(new_n660), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n891), .A2(new_n799), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n849), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n896));
  AOI211_X1 g710(.A(new_n331), .B(new_n731), .C1(new_n706), .C2(new_n704), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n881), .A3(new_n882), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT50), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n897), .A2(new_n881), .A3(KEYINPUT119), .A4(new_n882), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n896), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n896), .A3(new_n901), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT50), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n903), .B1(new_n904), .B2(new_n898), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n889), .B(new_n895), .C1(new_n902), .C2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT51), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n886), .B1(new_n824), .B2(new_n825), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n907), .B1(new_n909), .B2(new_n884), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n895), .B(new_n910), .C1(new_n905), .C2(new_n902), .ZN(new_n911));
  INV_X1    g725(.A(new_n853), .ZN(new_n912));
  OAI221_X1 g726(.A(new_n320), .B1(new_n883), .B2(new_n912), .C1(new_n892), .C2(new_n661), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n894), .A2(new_n776), .A3(new_n777), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n914), .A2(KEYINPUT48), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(KEYINPUT48), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n908), .A2(new_n911), .A3(new_n917), .ZN(new_n918));
  OAI22_X1  g732(.A1(new_n880), .A2(new_n918), .B1(G952), .B2(G953), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n632), .A2(new_n506), .A3(new_n331), .ZN(new_n920));
  INV_X1    g734(.A(new_n771), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n797), .B(new_n920), .C1(new_n921), .C2(KEYINPUT49), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n706), .A2(new_n704), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n921), .A2(KEYINPUT49), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n922), .A2(new_n890), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT114), .Z(new_n926));
  NAND2_X1  g740(.A1(new_n919), .A2(new_n926), .ZN(G75));
  AOI21_X1  g741(.A(new_n326), .B1(new_n876), .B2(new_n878), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n188), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n315), .B(new_n228), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT55), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n929), .B2(new_n930), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n189), .A2(G952), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(G51));
  XOR2_X1   g750(.A(new_n807), .B(KEYINPUT57), .Z(new_n937));
  INV_X1    g751(.A(new_n879), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n877), .B1(new_n876), .B2(new_n878), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n500), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n808), .A2(new_n809), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n928), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n935), .B1(new_n941), .B2(new_n943), .ZN(G54));
  AND2_X1   g758(.A1(KEYINPUT58), .A2(G475), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n749), .A2(new_n766), .A3(new_n844), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n633), .A2(new_n841), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n431), .A2(new_n507), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n948), .B1(new_n683), .B2(KEYINPUT102), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n947), .B1(new_n686), .B2(new_n949), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n848), .A2(new_n795), .A3(new_n850), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n946), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI22_X1  g766(.A1(new_n786), .A2(new_n787), .B1(new_n781), .B2(new_n790), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(KEYINPUT53), .B1(new_n954), .B2(new_n860), .ZN(new_n955));
  AND4_X1   g769(.A1(KEYINPUT53), .A2(new_n852), .A3(new_n792), .A4(new_n870), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n325), .B(new_n945), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n651), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n935), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n928), .A2(new_n651), .A3(new_n945), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT121), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n959), .A2(new_n961), .A3(KEYINPUT121), .A4(new_n960), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(G60));
  NAND2_X1  g780(.A1(G478), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT59), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n655), .B(new_n968), .C1(new_n938), .C2(new_n939), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n960), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n655), .B1(new_n880), .B2(new_n968), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(G63));
  INV_X1    g786(.A(KEYINPUT61), .ZN(new_n973));
  NAND2_X1  g787(.A1(G217), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT60), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n876), .B2(new_n878), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n675), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n960), .B1(new_n976), .B2(new_n619), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n973), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n976), .A2(new_n619), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n981), .A2(KEYINPUT61), .A3(new_n960), .A4(new_n977), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(G66));
  INV_X1    g797(.A(G224), .ZN(new_n984));
  OAI21_X1  g798(.A(G953), .B1(new_n328), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n843), .A2(new_n845), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(G953), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n293), .B(new_n294), .C1(G898), .C2(new_n189), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT122), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n987), .B(new_n989), .ZN(G69));
  NAND2_X1  g804(.A1(new_n556), .A2(new_n557), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(new_n366), .Z(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n698), .A2(new_n717), .A3(new_n854), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n714), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT62), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n994), .A2(new_n714), .A3(KEYINPUT62), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n839), .A2(new_n834), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n778), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n1000), .A2(new_n701), .ZN(new_n1001));
  AOI22_X1  g815(.A1(new_n997), .A2(new_n998), .B1(new_n723), .B2(new_n1001), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n1002), .A2(new_n820), .A3(new_n828), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n993), .B1(new_n1003), .B2(G953), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n693), .A2(G953), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT123), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n776), .A2(new_n777), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n815), .A2(new_n691), .A3(new_n1007), .A4(new_n708), .ZN(new_n1008));
  AND4_X1   g822(.A1(new_n820), .A2(new_n828), .A3(new_n994), .A4(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT124), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n792), .A2(new_n1010), .A3(new_n795), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1010), .B1(new_n792), .B2(new_n795), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1006), .B1(new_n1013), .B2(new_n189), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1004), .B1(new_n1014), .B2(new_n993), .ZN(new_n1015));
  INV_X1    g829(.A(G227), .ZN(new_n1016));
  OAI221_X1 g830(.A(G953), .B1(new_n1016), .B2(new_n693), .C1(new_n993), .C2(KEYINPUT125), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g833(.A(new_n1017), .B(new_n1004), .C1(new_n1014), .C2(new_n993), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(G72));
  INV_X1    g835(.A(KEYINPUT127), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1002), .A2(new_n820), .A3(new_n828), .A4(new_n986), .ZN(new_n1023));
  NAND2_X1  g837(.A1(G472), .A2(G902), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1024), .B(KEYINPUT63), .Z(new_n1025));
  NAND2_X1  g839(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1026), .A2(new_n539), .A3(new_n559), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1025), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1028), .B1(new_n572), .B2(new_n560), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT126), .Z(new_n1030));
  AOI21_X1  g844(.A(new_n935), .B1(new_n872), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n559), .A2(new_n539), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1033), .ZN(new_n1034));
  OAI211_X1 g848(.A(new_n1009), .B(new_n986), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1034), .B1(new_n1035), .B2(new_n1025), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1022), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1035), .A2(new_n1025), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1038), .A2(new_n1033), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n1039), .A2(KEYINPUT127), .A3(new_n1027), .A4(new_n1031), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1037), .A2(new_n1040), .ZN(G57));
endmodule


