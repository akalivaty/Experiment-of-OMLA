//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n202));
  XNOR2_X1  g001(.A(G211gat), .B(G218gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT76), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n206));
  OR2_X1    g005(.A1(G197gat), .A2(G204gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G197gat), .A2(G204gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n209), .B(KEYINPUT77), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(KEYINPUT77), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n204), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G226gat), .A2(G233gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT27), .B(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(G190gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT70), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT28), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n218), .A2(new_n221), .A3(new_n222), .A4(new_n219), .ZN(new_n226));
  AND3_X1   g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT71), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n228), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n230));
  AND3_X1   g029(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT71), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT72), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT69), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT26), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(G169gat), .B2(G176gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n238), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G169gat), .A2(G176gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT72), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n247), .A2(new_n248), .A3(new_n229), .A4(new_n234), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n236), .A2(new_n242), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n227), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n237), .A2(KEYINPUT23), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT23), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(G169gat), .B2(G176gat), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n254), .B(new_n256), .C1(new_n230), .C2(new_n231), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n258));
  NAND3_X1  g057(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT65), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n262), .A2(new_n225), .B1(new_n259), .B2(new_n260), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n257), .A2(new_n258), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n247), .A2(KEYINPUT67), .A3(new_n256), .A4(new_n254), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n253), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(new_n225), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n259), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n238), .A2(KEYINPUT23), .A3(new_n241), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n245), .A2(KEYINPUT68), .A3(new_n246), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT25), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n272), .B1(new_n273), .B2(new_n247), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n251), .B1(new_n266), .B2(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(KEYINPUT78), .B(KEYINPUT29), .Z(new_n277));
  AOI21_X1  g076(.A(new_n217), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n257), .A2(new_n258), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n261), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(new_n265), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n252), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n271), .A2(new_n274), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n282), .A2(new_n283), .B1(new_n250), .B2(new_n227), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(new_n216), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n202), .B(new_n215), .C1(new_n278), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n276), .A2(new_n217), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n284), .A2(KEYINPUT29), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n214), .B(new_n287), .C1(new_n288), .C2(new_n217), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n277), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n216), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n287), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n202), .B1(new_n293), .B2(new_n215), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT37), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G8gat), .B(G36gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT80), .ZN(new_n297));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n215), .B1(new_n278), .B2(new_n285), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT79), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT37), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n302), .A2(new_n303), .A3(new_n289), .A4(new_n286), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n295), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT38), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n303), .B1(new_n293), .B2(new_n214), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n287), .B1(new_n288), .B2(new_n217), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n307), .B1(new_n214), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT38), .ZN(new_n310));
  XOR2_X1   g109(.A(new_n299), .B(KEYINPUT81), .Z(new_n311));
  NAND4_X1  g110(.A1(new_n304), .A2(new_n309), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT86), .B(KEYINPUT5), .ZN(new_n313));
  INV_X1    g112(.A(G113gat), .ZN(new_n314));
  INV_X1    g113(.A(G120gat), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT1), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G127gat), .B(G134gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT73), .B(G120gat), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n316), .B(new_n317), .C1(new_n318), .C2(new_n314), .ZN(new_n319));
  INV_X1    g118(.A(G134gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G127gat), .ZN(new_n321));
  INV_X1    g120(.A(G127gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G134gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n314), .A2(new_n315), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n326), .B1(G113gat), .B2(G120gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n324), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n319), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT83), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT2), .ZN(new_n332));
  INV_X1    g131(.A(G141gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(G148gat), .ZN(new_n334));
  INV_X1    g133(.A(G148gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n335), .A2(G141gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n332), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  XOR2_X1   g136(.A(G155gat), .B(G162gat), .Z(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT82), .B1(new_n333), .B2(G148gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT82), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(new_n335), .A3(G141gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n333), .A2(G148gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n340), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G155gat), .ZN(new_n345));
  INV_X1    g144(.A(G162gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n332), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n339), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n319), .A2(KEYINPUT83), .A3(new_n328), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n331), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT85), .B1(new_n351), .B2(new_n329), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n324), .A2(new_n327), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n315), .A2(KEYINPUT73), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n315), .A2(KEYINPUT73), .ZN(new_n357));
  OAI21_X1  g156(.A(G113gat), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n316), .B1(new_n314), .B2(new_n315), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n355), .A2(new_n358), .B1(new_n359), .B2(new_n324), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n337), .A2(new_n338), .B1(new_n344), .B2(new_n349), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT85), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n353), .A2(new_n354), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n313), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n351), .A2(KEYINPUT3), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n361), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n368), .A2(new_n370), .A3(new_n331), .A4(new_n352), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT4), .B1(new_n354), .B2(new_n363), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n351), .A2(new_n329), .ZN(new_n373));
  XOR2_X1   g172(.A(KEYINPUT84), .B(KEYINPUT4), .Z(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n365), .B(new_n371), .C1(new_n372), .C2(new_n375), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n371), .A2(new_n365), .A3(new_n313), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n354), .A2(KEYINPUT4), .A3(new_n363), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT87), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n373), .A2(new_n379), .A3(new_n374), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n360), .A2(new_n361), .ZN(new_n381));
  INV_X1    g180(.A(new_n374), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT87), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n378), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n367), .A2(new_n376), .B1(new_n377), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G1gat), .B(G29gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT0), .ZN(new_n387));
  XNOR2_X1  g186(.A(G57gat), .B(G85gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT6), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n367), .A2(new_n376), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n384), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n389), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(KEYINPUT6), .A3(new_n389), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n302), .A2(new_n289), .A3(new_n286), .A4(new_n299), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n306), .A2(new_n312), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(G228gat), .ZN(new_n401));
  INV_X1    g200(.A(G233gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n214), .A2(new_n277), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n361), .B1(new_n405), .B2(new_n369), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n291), .B1(new_n361), .B2(new_n369), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n214), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n404), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT3), .B1(new_n214), .B2(new_n410), .ZN(new_n411));
  OAI221_X1 g210(.A(new_n403), .B1(new_n214), .B2(new_n407), .C1(new_n411), .C2(new_n361), .ZN(new_n412));
  XNOR2_X1  g211(.A(G78gat), .B(G106gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT88), .ZN(new_n414));
  XOR2_X1   g213(.A(KEYINPUT31), .B(G50gat), .Z(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(KEYINPUT89), .A2(G22gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(G22gat), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n418), .B1(new_n419), .B2(new_n416), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n409), .A2(new_n412), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n421), .B1(new_n409), .B2(new_n412), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n365), .B1(new_n384), .B2(new_n371), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT90), .B(KEYINPUT39), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n389), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT91), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT39), .B1(new_n364), .B2(new_n366), .ZN(new_n430));
  OAI22_X1  g229(.A1(new_n428), .A2(new_n429), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  AOI211_X1 g230(.A(KEYINPUT91), .B(new_n389), .C1(new_n426), .C2(new_n427), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT92), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT40), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT40), .ZN(new_n435));
  OAI211_X1 g234(.A(KEYINPUT92), .B(new_n435), .C1(new_n431), .C2(new_n432), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n395), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT30), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n311), .B1(new_n290), .B2(new_n294), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n438), .B1(new_n439), .B2(new_n398), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n398), .A2(new_n438), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n400), .B(new_n425), .C1(new_n437), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n439), .A2(new_n398), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT30), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n396), .A2(new_n397), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n447), .A3(new_n441), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n281), .A2(new_n252), .B1(new_n271), .B2(new_n274), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n450));
  INV_X1    g249(.A(new_n242), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n247), .A2(new_n234), .A3(new_n229), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n451), .B1(new_n452), .B2(KEYINPUT72), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n450), .B1(new_n453), .B2(new_n249), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n360), .B1(new_n449), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(G227gat), .A2(G233gat), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n251), .B(new_n329), .C1(new_n275), .C2(new_n266), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n455), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT32), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(KEYINPUT74), .B(G71gat), .Z(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(G99gat), .ZN(new_n466));
  XOR2_X1   g265(.A(G15gat), .B(G43gat), .Z(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n457), .B1(new_n455), .B2(new_n458), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT34), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(new_n456), .B2(KEYINPUT75), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  AOI211_X1 g274(.A(new_n457), .B(new_n473), .C1(new_n455), .C2(new_n458), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n470), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n468), .B1(new_n459), .B2(new_n463), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n471), .A2(new_n474), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(new_n476), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n462), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n478), .A2(new_n462), .A3(new_n481), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(KEYINPUT36), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT36), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n478), .A2(new_n462), .A3(new_n481), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n486), .B1(new_n487), .B2(new_n482), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n448), .A2(new_n424), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n483), .A2(new_n425), .A3(new_n484), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT35), .B1(new_n448), .B2(new_n490), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n487), .A2(new_n482), .A3(new_n424), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT35), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n492), .A2(new_n443), .A3(new_n493), .A4(new_n447), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n444), .A2(new_n489), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT18), .ZN(new_n496));
  INV_X1    g295(.A(G1gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT16), .ZN(new_n498));
  INV_X1    g297(.A(G15gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(G22gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n419), .A2(G15gat), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(G1gat), .B1(new_n500), .B2(new_n501), .ZN(new_n503));
  OAI21_X1  g302(.A(G8gat), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n505));
  INV_X1    g304(.A(G8gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(G15gat), .B(G22gat), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n505), .B(new_n506), .C1(G1gat), .C2(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G50gat), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(KEYINPUT94), .A3(G43gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT15), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT94), .ZN(new_n514));
  XNOR2_X1  g313(.A(G43gat), .B(G50gat), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT14), .ZN(new_n517));
  INV_X1    g316(.A(G29gat), .ZN(new_n518));
  INV_X1    g317(.A(G36gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n510), .A2(G43gat), .ZN(new_n523));
  INV_X1    g322(.A(G43gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(G50gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n525), .A3(KEYINPUT15), .ZN(new_n526));
  NAND2_X1  g325(.A1(G29gat), .A2(G36gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n522), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n516), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n520), .A2(KEYINPUT93), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT93), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n531), .A2(new_n517), .A3(new_n518), .A4(new_n519), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n532), .A3(new_n521), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n526), .B1(new_n533), .B2(new_n527), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n529), .A2(new_n534), .A3(KEYINPUT17), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n536));
  NOR3_X1   g335(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n521), .B1(new_n537), .B2(new_n531), .ZN(new_n538));
  INV_X1    g337(.A(new_n532), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n527), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n526), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n523), .A2(new_n525), .A3(new_n514), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n543), .A2(new_n512), .A3(new_n511), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n544), .A2(new_n526), .A3(new_n527), .A4(new_n522), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n536), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n509), .B1(new_n535), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n542), .A2(new_n545), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n504), .A2(new_n508), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n548), .A2(new_n549), .B1(G229gat), .B2(G233gat), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n496), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT17), .B1(new_n529), .B2(new_n534), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n542), .A2(new_n536), .A3(new_n545), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n522), .A2(new_n526), .A3(new_n527), .ZN(new_n556));
  AOI22_X1  g355(.A1(new_n541), .A2(new_n540), .B1(new_n556), .B2(new_n544), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n555), .B1(new_n557), .B2(new_n509), .ZN(new_n558));
  NOR3_X1   g357(.A1(new_n554), .A2(KEYINPUT18), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n548), .A2(new_n549), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n542), .A2(new_n545), .A3(new_n504), .A4(new_n508), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n555), .B(KEYINPUT13), .Z(new_n563));
  AOI21_X1  g362(.A(KEYINPUT95), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT95), .ZN(new_n565));
  INV_X1    g364(.A(new_n563), .ZN(new_n566));
  AOI211_X1 g365(.A(new_n565), .B(new_n566), .C1(new_n560), .C2(new_n561), .ZN(new_n567));
  OAI22_X1  g366(.A1(new_n551), .A2(new_n559), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G113gat), .B(G141gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(G197gat), .ZN(new_n570));
  XOR2_X1   g369(.A(KEYINPUT11), .B(G169gat), .Z(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT12), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT96), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n547), .A2(new_n496), .A3(new_n550), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT18), .B1(new_n554), .B2(new_n558), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NOR3_X1   g378(.A1(new_n549), .A2(new_n529), .A3(new_n534), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n542), .A2(new_n545), .B1(new_n504), .B2(new_n508), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n563), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n565), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n562), .A2(KEYINPUT95), .A3(new_n563), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n579), .A2(new_n585), .A3(new_n573), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n575), .A2(new_n576), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n568), .A2(KEYINPUT96), .A3(new_n574), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n495), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(G57gat), .ZN(new_n595));
  INV_X1    g394(.A(G64gat), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n592), .B1(KEYINPUT9), .B2(new_n593), .ZN(new_n600));
  OAI21_X1  g399(.A(G64gat), .B1(new_n595), .B2(KEYINPUT97), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT97), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(new_n596), .A3(G57gat), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n599), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT98), .ZN(new_n608));
  XNOR2_X1  g407(.A(G127gat), .B(G155gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT99), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n608), .B(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n509), .B1(new_n606), .B2(new_n605), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT100), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n613), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n616));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(G183gat), .B(G211gat), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n614), .A2(new_n615), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n620), .B1(new_n614), .B2(new_n615), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(G99gat), .B(G106gat), .Z(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G85gat), .A2(G92gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT7), .ZN(new_n627));
  NOR2_X1   g426(.A1(G85gat), .A2(G92gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(G99gat), .A2(G106gat), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n628), .B1(KEYINPUT8), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n625), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n625), .B1(new_n627), .B2(new_n630), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(G232gat), .A2(G233gat), .ZN(new_n635));
  AOI22_X1  g434(.A1(new_n634), .A2(new_n548), .B1(KEYINPUT41), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n535), .A2(new_n546), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n636), .B1(new_n637), .B2(new_n634), .ZN(new_n638));
  XOR2_X1   g437(.A(G190gat), .B(G218gat), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n635), .A2(KEYINPUT41), .ZN(new_n641));
  XNOR2_X1  g440(.A(G134gat), .B(G162gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n640), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n605), .B1(new_n632), .B2(new_n633), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n593), .A2(KEYINPUT9), .ZN(new_n647));
  AOI22_X1  g446(.A1(new_n591), .A2(new_n647), .B1(new_n601), .B2(new_n603), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n597), .A2(new_n598), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(new_n649), .B2(new_n594), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n627), .A2(new_n630), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n624), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n650), .A2(new_n631), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT10), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n646), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n634), .A2(KEYINPUT10), .A3(new_n650), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(G230gat), .A2(G233gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT101), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n653), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n659), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G120gat), .B(G148gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT102), .ZN(new_n666));
  XNOR2_X1  g465(.A(G176gat), .B(G204gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n661), .A2(new_n663), .A3(new_n668), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n623), .A2(new_n645), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n590), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n447), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(new_n497), .ZN(G1324gat));
  NOR2_X1   g477(.A1(new_n676), .A2(new_n443), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT103), .B1(new_n679), .B2(new_n506), .ZN(new_n680));
  OR3_X1    g479(.A1(new_n679), .A2(KEYINPUT103), .A3(new_n506), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT16), .B(G8gat), .Z(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n683), .A2(KEYINPUT42), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(KEYINPUT42), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n680), .B(new_n681), .C1(new_n684), .C2(new_n685), .ZN(G1325gat));
  INV_X1    g485(.A(new_n676), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n487), .A2(new_n482), .ZN(new_n688));
  AOI21_X1  g487(.A(G15gat), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n485), .A2(new_n488), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n499), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT104), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n689), .B1(new_n687), .B2(new_n692), .ZN(G1326gat));
  NOR2_X1   g492(.A1(new_n676), .A2(new_n425), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT43), .B(G22gat), .Z(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  INV_X1    g495(.A(new_n623), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n673), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n698), .A2(new_n645), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n590), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n447), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n518), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT45), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n444), .A2(new_n489), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n491), .A2(new_n494), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n707), .A2(KEYINPUT44), .A3(new_n644), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n709), .B1(new_n495), .B2(new_n645), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n586), .A2(new_n576), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n573), .B1(new_n579), .B2(new_n585), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n588), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n711), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n587), .A2(KEYINPUT105), .A3(new_n588), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n698), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n708), .A2(new_n710), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT106), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n708), .A2(new_n710), .A3(new_n722), .A4(new_n719), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n721), .A2(new_n702), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n704), .B1(new_n518), .B2(new_n724), .ZN(G1328gat));
  NOR2_X1   g524(.A1(new_n443), .A2(G36gat), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  OR3_X1    g526(.A1(new_n700), .A2(KEYINPUT107), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT107), .B1(new_n700), .B2(new_n727), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n728), .A2(KEYINPUT46), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT46), .B1(new_n728), .B2(new_n729), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n443), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n721), .A2(new_n733), .A3(new_n723), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n721), .A2(KEYINPUT108), .A3(new_n733), .A4(new_n723), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n736), .A2(G36gat), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n732), .A2(new_n738), .ZN(G1329gat));
  OAI21_X1  g538(.A(G43gat), .B1(new_n720), .B2(new_n690), .ZN(new_n740));
  INV_X1    g539(.A(new_n688), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(G43gat), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n701), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n740), .A2(KEYINPUT47), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n690), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n721), .A2(new_n745), .A3(new_n723), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n746), .A2(G43gat), .B1(new_n701), .B2(new_n742), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n744), .B1(new_n747), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g547(.A1(new_n700), .A2(G50gat), .A3(new_n425), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n721), .A2(new_n424), .A3(new_n723), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n749), .B1(new_n750), .B2(G50gat), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n720), .A2(new_n425), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n510), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT48), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  OAI22_X1  g554(.A1(new_n751), .A2(KEYINPUT48), .B1(new_n753), .B2(new_n755), .ZN(G1331gat));
  NAND4_X1  g555(.A1(new_n718), .A2(new_n623), .A3(new_n645), .A4(new_n672), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT109), .Z(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n707), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n447), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(new_n595), .ZN(G1332gat));
  NOR2_X1   g560(.A1(new_n759), .A2(new_n443), .ZN(new_n762));
  NOR2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  AND2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n762), .B2(new_n763), .ZN(G1333gat));
  OAI21_X1  g565(.A(G71gat), .B1(new_n759), .B2(new_n690), .ZN(new_n767));
  INV_X1    g566(.A(G71gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n688), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n759), .B2(new_n769), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g570(.A1(new_n759), .A2(new_n425), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n772), .B(G78gat), .Z(G1335gat));
  AOI21_X1  g572(.A(new_n645), .B1(new_n705), .B2(new_n706), .ZN(new_n774));
  INV_X1    g573(.A(new_n718), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n623), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT51), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  INV_X1    g578(.A(new_n776), .ZN(new_n780));
  NOR4_X1   g579(.A1(new_n495), .A2(new_n779), .A3(new_n780), .A4(new_n645), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n778), .A2(new_n782), .A3(KEYINPUT111), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n777), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n447), .A2(G85gat), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n783), .A2(new_n672), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n708), .A2(new_n710), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n780), .A2(new_n673), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n702), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT110), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G85gat), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n790), .A2(KEYINPUT110), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n787), .B1(new_n792), .B2(new_n793), .ZN(G1336gat));
  NAND3_X1  g593(.A1(new_n788), .A2(new_n733), .A3(new_n789), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G92gat), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n443), .A2(G92gat), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n672), .B(new_n797), .C1(new_n777), .C2(new_n781), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT52), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n672), .A3(new_n785), .A4(new_n797), .ZN(new_n801));
  XOR2_X1   g600(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n796), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n800), .A2(new_n803), .ZN(G1337gat));
  NOR3_X1   g603(.A1(new_n741), .A2(G99gat), .A3(new_n673), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n783), .A2(new_n785), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n788), .A2(new_n745), .A3(new_n789), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G99gat), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(G1338gat));
  NAND4_X1  g608(.A1(new_n708), .A2(new_n710), .A3(new_n424), .A4(new_n789), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G106gat), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n425), .A2(G106gat), .A3(new_n673), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n777), .B2(new_n781), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT114), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n810), .A2(KEYINPUT113), .A3(G106gat), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n818), .B(new_n814), .C1(new_n777), .C2(new_n781), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n813), .A2(new_n816), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT53), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n783), .A2(new_n785), .A3(new_n814), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n810), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(G106gat), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n824), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n822), .B(new_n823), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n821), .A2(new_n828), .ZN(G1339gat));
  NAND3_X1  g628(.A1(new_n655), .A2(new_n656), .A3(new_n659), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n661), .A2(KEYINPUT54), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n659), .B1(new_n655), .B2(new_n656), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n668), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(KEYINPUT55), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n671), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT55), .B1(new_n831), .B2(new_n834), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n716), .A2(new_n717), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n555), .B1(new_n547), .B2(new_n560), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n562), .A2(new_n563), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n572), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n586), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n840), .B1(new_n845), .B2(new_n672), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n673), .A2(new_n844), .A3(KEYINPUT116), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n644), .B1(new_n839), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n644), .A2(new_n838), .A3(new_n845), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n697), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n775), .A2(new_n674), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n424), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n733), .A2(new_n447), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(new_n688), .A3(new_n856), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n857), .A2(new_n314), .A3(new_n589), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n587), .A2(KEYINPUT105), .A3(new_n588), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT105), .B1(new_n587), .B2(new_n588), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n836), .A2(new_n837), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n846), .A2(new_n847), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n645), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n623), .B1(new_n864), .B2(new_n850), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n702), .B(new_n492), .C1(new_n865), .C2(new_n853), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n447), .B1(new_n852), .B2(new_n854), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(KEYINPUT117), .A3(new_n492), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n733), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n775), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n858), .B1(new_n872), .B2(new_n314), .ZN(G1340gat));
  NAND3_X1  g672(.A1(new_n871), .A2(new_n318), .A3(new_n672), .ZN(new_n874));
  OAI21_X1  g673(.A(G120gat), .B1(new_n857), .B2(new_n673), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1341gat));
  NOR3_X1   g675(.A1(new_n857), .A2(new_n322), .A3(new_n697), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT118), .ZN(new_n878));
  AOI21_X1  g677(.A(G127gat), .B1(new_n871), .B2(new_n623), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(G1342gat));
  INV_X1    g679(.A(KEYINPUT56), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n645), .A2(G134gat), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT117), .B1(new_n869), .B2(new_n492), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n443), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(KEYINPUT119), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n887), .B1(new_n871), .B2(new_n882), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n881), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(G134gat), .B1(new_n857), .B2(new_n645), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n885), .A2(KEYINPUT119), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n871), .A2(new_n887), .A3(new_n882), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(KEYINPUT56), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n889), .A2(new_n890), .A3(new_n893), .ZN(G1343gat));
  AND4_X1   g693(.A1(new_n443), .A2(new_n869), .A3(new_n424), .A4(new_n690), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n589), .A2(G141gat), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT58), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n425), .B1(new_n852), .B2(new_n854), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT57), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n856), .A2(new_n690), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n845), .A2(new_n672), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(new_n861), .B2(new_n589), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n645), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n623), .B1(new_n904), .B2(new_n850), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n424), .B1(new_n905), .B2(new_n853), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n901), .B1(new_n906), .B2(KEYINPUT57), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n900), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(G141gat), .B1(new_n908), .B2(new_n589), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n897), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n900), .A2(KEYINPUT120), .A3(new_n907), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n913), .A3(new_n775), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n914), .A2(G141gat), .B1(new_n895), .B2(new_n896), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n910), .B1(new_n915), .B2(new_n916), .ZN(G1344gat));
  NOR2_X1   g716(.A1(new_n335), .A2(KEYINPUT59), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n912), .A2(new_n913), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n673), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n714), .A2(new_n715), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n838), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n644), .B1(new_n922), .B2(new_n902), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n697), .B1(new_n923), .B2(new_n851), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n675), .A2(new_n589), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n425), .A2(KEYINPUT57), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n672), .B(new_n928), .C1(new_n898), .C2(new_n899), .ZN(new_n929));
  OAI21_X1  g728(.A(G148gat), .B1(new_n929), .B2(new_n901), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT59), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n920), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n895), .A2(new_n335), .A3(new_n672), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1345gat));
  OAI21_X1  g733(.A(G155gat), .B1(new_n919), .B2(new_n697), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n895), .A2(new_n345), .A3(new_n623), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1346gat));
  OAI21_X1  g736(.A(G162gat), .B1(new_n919), .B2(new_n645), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n895), .A2(new_n346), .A3(new_n644), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1347gat));
  AOI21_X1  g739(.A(new_n702), .B1(new_n852), .B2(new_n854), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n941), .A2(new_n733), .A3(new_n492), .ZN(new_n942));
  AOI21_X1  g741(.A(G169gat), .B1(new_n942), .B2(new_n775), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n741), .A2(new_n443), .A3(new_n702), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n855), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n921), .A2(G169gat), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(G1348gat));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n672), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n673), .A2(G176gat), .ZN(new_n949));
  AOI22_X1  g748(.A1(new_n948), .A2(G176gat), .B1(new_n942), .B2(new_n949), .ZN(new_n950));
  XOR2_X1   g749(.A(new_n950), .B(KEYINPUT121), .Z(G1349gat));
  NAND3_X1  g750(.A1(new_n855), .A2(new_n623), .A3(new_n944), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n952), .A2(KEYINPUT122), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(KEYINPUT122), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(G183gat), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n942), .A2(new_n218), .A3(new_n623), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(KEYINPUT60), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT60), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n955), .A2(new_n959), .A3(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(G1350gat));
  NAND3_X1  g760(.A1(new_n942), .A2(new_n219), .A3(new_n644), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n644), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G190gat), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n964), .A2(KEYINPUT61), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n964), .A2(KEYINPUT61), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(G1351gat));
  INV_X1    g766(.A(new_n927), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n968), .B1(new_n924), .B2(new_n925), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n424), .B1(new_n865), .B2(new_n853), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n969), .B1(new_n970), .B2(KEYINPUT57), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n443), .A2(new_n702), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(new_n690), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n921), .A2(G197gat), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n745), .A2(new_n443), .A3(new_n425), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n941), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n978), .A2(new_n718), .ZN(new_n979));
  OAI22_X1  g778(.A1(new_n975), .A2(new_n976), .B1(G197gat), .B2(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(G1352gat));
  INV_X1    g780(.A(KEYINPUT123), .ZN(new_n982));
  NAND4_X1  g781(.A1(new_n971), .A2(new_n982), .A3(new_n672), .A4(new_n974), .ZN(new_n983));
  OAI21_X1  g782(.A(KEYINPUT123), .B1(new_n929), .B2(new_n973), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n983), .A2(new_n984), .A3(G204gat), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n673), .A2(G204gat), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n941), .A2(new_n977), .A3(new_n986), .ZN(new_n987));
  XOR2_X1   g786(.A(new_n987), .B(KEYINPUT62), .Z(new_n988));
  NAND2_X1  g787(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(KEYINPUT124), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT124), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n985), .A2(new_n991), .A3(new_n988), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n992), .ZN(G1353gat));
  INV_X1    g792(.A(G211gat), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT63), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n994), .B1(KEYINPUT126), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n996), .B1(new_n975), .B2(new_n697), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT126), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n997), .A2(new_n998), .A3(KEYINPUT63), .ZN(new_n999));
  OAI221_X1 g798(.A(new_n996), .B1(KEYINPUT126), .B2(new_n995), .C1(new_n975), .C2(new_n697), .ZN(new_n1000));
  NOR3_X1   g799(.A1(new_n978), .A2(G211gat), .A3(new_n697), .ZN(new_n1001));
  XNOR2_X1  g800(.A(new_n1001), .B(KEYINPUT125), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(G1354gat));
  NAND2_X1  g802(.A1(new_n975), .A2(KEYINPUT127), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1004), .A2(new_n644), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n975), .A2(KEYINPUT127), .ZN(new_n1006));
  OAI21_X1  g805(.A(G218gat), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OR3_X1    g806(.A1(new_n978), .A2(G218gat), .A3(new_n645), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1007), .A2(new_n1008), .ZN(G1355gat));
endmodule


