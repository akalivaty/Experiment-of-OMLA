//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n565, new_n566, new_n567,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n616, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1119;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n467), .B(KEYINPUT66), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n469), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n471), .A2(G2105), .B1(G101), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G112), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n466), .A2(G136), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n465), .A2(new_n472), .ZN(new_n482));
  AOI211_X1 g057(.A(new_n479), .B(new_n481), .C1(G124), .C2(new_n482), .ZN(G162));
  INV_X1    g058(.A(G138), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n466), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n466), .B(new_n486), .C1(new_n485), .C2(KEYINPUT4), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n482), .B2(G126), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n489), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n499), .A2(new_n501), .B1(new_n498), .B2(G543), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n504), .A2(KEYINPUT68), .A3(KEYINPUT6), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n502), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n505), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n509), .A2(new_n510), .ZN(new_n520));
  INV_X1    g095(.A(new_n506), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n520), .A2(G51), .A3(G543), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n498), .A2(G543), .ZN(new_n523));
  AND2_X1   g098(.A1(G63), .A2(G651), .ZN(new_n524));
  INV_X1    g099(.A(new_n501), .ZN(new_n525));
  AOI21_X1  g100(.A(KEYINPUT69), .B1(new_n500), .B2(KEYINPUT5), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n523), .B(new_n524), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT70), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT70), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n522), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n502), .A2(new_n511), .A3(G89), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n519), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n533), .A2(new_n535), .ZN(new_n538));
  AOI211_X1 g113(.A(KEYINPUT71), .B(new_n538), .C1(new_n529), .C2(new_n531), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  AOI22_X1  g116(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n504), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  INV_X1    g119(.A(G52), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n512), .A2(new_n544), .B1(new_n514), .B2(new_n545), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n543), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  AOI22_X1  g123(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(KEYINPUT72), .B1(new_n549), .B2(new_n504), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n502), .A2(new_n511), .A3(G81), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n511), .A2(G43), .A3(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  OAI211_X1 g129(.A(G56), .B(new_n523), .C1(new_n525), .C2(new_n526), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT72), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n557), .A2(new_n558), .A3(G651), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n550), .A2(new_n554), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT73), .Z(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g139(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n565));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  XNOR2_X1  g143(.A(KEYINPUT75), .B(G65), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n523), .B(new_n569), .C1(new_n525), .C2(new_n526), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n504), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n502), .A2(new_n511), .A3(G91), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n520), .A2(G53), .A3(G543), .A4(new_n521), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT9), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n511), .A2(new_n577), .A3(G53), .A4(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n574), .A2(KEYINPUT76), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(KEYINPUT76), .B1(new_n574), .B2(new_n579), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n580), .A2(new_n581), .ZN(G299));
  INV_X1    g157(.A(new_n512), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G87), .ZN(new_n584));
  INV_X1    g159(.A(new_n514), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G49), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(G288));
  AOI22_X1  g163(.A1(new_n502), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n504), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n511), .A2(G48), .A3(G543), .ZN(new_n591));
  INV_X1    g166(.A(G86), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n512), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(G85), .A2(new_n583), .B1(new_n585), .B2(G47), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n504), .B2(new_n597), .ZN(G290));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NOR2_X1   g174(.A1(G301), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n583), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n502), .A2(new_n511), .A3(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n502), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G54), .ZN(new_n607));
  OAI22_X1  g182(.A1(new_n606), .A2(new_n504), .B1(new_n607), .B2(new_n514), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT77), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n600), .B1(new_n611), .B2(new_n599), .ZN(G284));
  AOI21_X1  g187(.A(new_n600), .B1(new_n611), .B2(new_n599), .ZN(G321));
  MUX2_X1   g188(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g189(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n611), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n560), .A2(new_n599), .ZN(new_n618));
  INV_X1    g193(.A(new_n611), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n619), .A2(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n618), .B1(new_n620), .B2(new_n599), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n466), .A2(G135), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n482), .A2(G123), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n472), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND3_X1  g203(.A1(new_n472), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n628), .A2(new_n633), .A3(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT78), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2430), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(KEYINPUT14), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n642), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2443), .B(G2446), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT79), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT80), .Z(new_n652));
  OAI21_X1  g227(.A(G14), .B1(new_n647), .B2(new_n650), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  XOR2_X1   g230(.A(KEYINPUT81), .B(KEYINPUT17), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  NAND3_X1  g235(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT82), .Z(new_n662));
  INV_X1    g237(.A(new_n655), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n663), .A2(new_n658), .A3(new_n660), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT18), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n657), .A2(new_n659), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n660), .B1(new_n659), .B2(new_n655), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2096), .B(G2100), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1956), .B(G2474), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1961), .B(G1966), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n673), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(new_n676), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT20), .Z(new_n680));
  AOI211_X1 g255(.A(new_n678), .B(new_n680), .C1(new_n673), .C2(new_n677), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G229));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G22), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G166), .B2(new_n688), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(G1971), .Z(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(G6), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(new_n594), .B2(new_n688), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT32), .B(G1981), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n688), .A2(G23), .ZN(new_n696));
  INV_X1    g271(.A(G288), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n688), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT33), .B(G1976), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT86), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n691), .A2(new_n695), .A3(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(KEYINPUT34), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(KEYINPUT34), .ZN(new_n704));
  NOR2_X1   g279(.A1(G16), .A2(G24), .ZN(new_n705));
  XOR2_X1   g280(.A(G290), .B(KEYINPUT85), .Z(new_n706));
  AOI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(G16), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(G1986), .Z(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G25), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT83), .ZN(new_n711));
  AOI22_X1  g286(.A1(G119), .A2(new_n482), .B1(new_n466), .B2(G131), .ZN(new_n712));
  OAI21_X1  g287(.A(KEYINPUT84), .B1(G95), .B2(G2105), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NOR3_X1   g289(.A1(KEYINPUT84), .A2(G95), .A3(G2105), .ZN(new_n715));
  OAI221_X1 g290(.A(G2104), .B1(G107), .B2(new_n472), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n711), .B1(new_n717), .B2(G29), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT35), .B(G1991), .Z(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n718), .B(new_n720), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n703), .A2(new_n704), .A3(new_n708), .A4(new_n721), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT36), .Z(new_n723));
  XOR2_X1   g298(.A(KEYINPUT31), .B(G11), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT92), .ZN(new_n725));
  INV_X1    g300(.A(G28), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(KEYINPUT30), .ZN(new_n727));
  AOI21_X1  g302(.A(G29), .B1(new_n726), .B2(KEYINPUT30), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(G164), .A2(G29), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G27), .B2(G29), .ZN(new_n731));
  INV_X1    g306(.A(G2078), .ZN(new_n732));
  OAI221_X1 g307(.A(new_n729), .B1(new_n709), .B2(new_n627), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n709), .A2(G35), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT93), .Z(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G162), .B2(new_n709), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT29), .B(G2090), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n733), .B(new_n738), .C1(new_n732), .C2(new_n731), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n709), .A2(G26), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT28), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n466), .A2(G140), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n482), .A2(G128), .ZN(new_n743));
  OR2_X1    g318(.A1(G104), .A2(G2105), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n744), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n741), .B1(new_n747), .B2(new_n709), .ZN(new_n748));
  INV_X1    g323(.A(G2067), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n709), .A2(G32), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n482), .A2(G129), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT91), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n473), .A2(G105), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT26), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n754), .B(new_n756), .C1(G141), .C2(new_n466), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n751), .B1(new_n758), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT27), .B(G1996), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n750), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n759), .B2(new_n760), .ZN(new_n762));
  NOR2_X1   g337(.A1(G171), .A2(new_n688), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G5), .B2(new_n688), .ZN(new_n764));
  INV_X1    g339(.A(G1961), .ZN(new_n765));
  NAND2_X1  g340(.A1(G115), .A2(G2104), .ZN(new_n766));
  INV_X1    g341(.A(G127), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n465), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n472), .B1(new_n768), .B2(KEYINPUT90), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(KEYINPUT90), .B2(new_n768), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT25), .ZN(new_n771));
  NAND2_X1  g346(.A1(G103), .A2(G2104), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G2105), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n472), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n466), .A2(G139), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(new_n709), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n709), .B2(G33), .ZN(new_n779));
  INV_X1    g354(.A(G2072), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n764), .A2(new_n765), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n739), .A2(new_n762), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n688), .A2(G19), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT89), .Z(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n561), .B2(new_n688), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1341), .ZN(new_n786));
  INV_X1    g361(.A(G34), .ZN(new_n787));
  AOI21_X1  g362(.A(G29), .B1(new_n787), .B2(KEYINPUT24), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(KEYINPUT24), .B2(new_n787), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n475), .B2(new_n709), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2084), .ZN(new_n791));
  OAI221_X1 g366(.A(new_n791), .B1(new_n779), .B2(new_n780), .C1(new_n765), .C2(new_n764), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n782), .A2(new_n786), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G21), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G168), .B2(G16), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1966), .Z(new_n796));
  NOR2_X1   g371(.A1(G4), .A2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT87), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n619), .B2(new_n688), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT88), .B(G1348), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(G299), .A2(G16), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n688), .A2(G20), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT23), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1956), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n793), .A2(new_n796), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n723), .A2(new_n808), .ZN(G311));
  INV_X1    g384(.A(G311), .ZN(G150));
  NAND2_X1  g385(.A1(new_n502), .A2(G67), .ZN(new_n811));
  INV_X1    g386(.A(G80), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(new_n500), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G651), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n502), .A2(new_n511), .A3(G93), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT94), .B(G55), .Z(new_n816));
  NAND3_X1  g391(.A1(new_n511), .A2(G543), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT95), .ZN(new_n818));
  AND3_X1   g393(.A1(new_n815), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n818), .B1(new_n815), .B2(new_n817), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n814), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G860), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT37), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n611), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n815), .A2(new_n817), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(KEYINPUT95), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n815), .A2(new_n817), .A3(new_n818), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n557), .A2(G651), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n553), .B1(new_n830), .B2(KEYINPUT72), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n829), .A2(new_n831), .A3(new_n559), .A4(new_n814), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n821), .A2(new_n560), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n825), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT96), .Z(new_n838));
  NOR2_X1   g413(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n839), .A2(G860), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n823), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT97), .Z(G145));
  XOR2_X1   g417(.A(new_n495), .B(KEYINPUT98), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n747), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(new_n758), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n777), .A2(KEYINPUT99), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n758), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n482), .A2(G130), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n472), .A2(G118), .ZN(new_n850));
  OAI21_X1  g425(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(G142), .B2(new_n466), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n630), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n848), .B(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n777), .A2(KEYINPUT99), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(new_n717), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n855), .B(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(G162), .B(new_n627), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n475), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(G37), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n858), .B2(new_n861), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT40), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(G395));
  NAND2_X1  g442(.A1(new_n821), .A2(new_n599), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n620), .B(new_n835), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n610), .B1(new_n580), .B2(new_n581), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT76), .ZN(new_n871));
  INV_X1    g446(.A(new_n579), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n502), .A2(new_n569), .B1(G78), .B2(G543), .ZN(new_n873));
  INV_X1    g448(.A(G91), .ZN(new_n874));
  OAI22_X1  g449(.A1(new_n873), .A2(new_n504), .B1(new_n874), .B2(new_n512), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n871), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n608), .B1(new_n604), .B2(new_n601), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n574), .A2(KEYINPUT76), .A3(new_n579), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n870), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n870), .A2(KEYINPUT100), .A3(new_n879), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n869), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT41), .B1(new_n870), .B2(new_n879), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n870), .A2(KEYINPUT41), .A3(new_n879), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n884), .B(new_n885), .C1(new_n869), .C2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n886), .A2(new_n892), .A3(KEYINPUT102), .ZN(new_n893));
  XNOR2_X1  g468(.A(G290), .B(new_n594), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n697), .B(G303), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n894), .B(new_n895), .Z(new_n896));
  XOR2_X1   g471(.A(new_n896), .B(KEYINPUT42), .Z(new_n897));
  NAND2_X1  g472(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT102), .B1(new_n886), .B2(new_n892), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n898), .B(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n868), .B1(new_n900), .B2(new_n599), .ZN(G295));
  OAI21_X1  g476(.A(new_n868), .B1(new_n900), .B2(new_n599), .ZN(G331));
  AND3_X1   g477(.A1(new_n522), .A2(new_n530), .A3(new_n527), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n530), .B1(new_n522), .B2(new_n527), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n536), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT71), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n536), .B(new_n519), .C1(new_n903), .C2(new_n904), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n906), .A2(new_n907), .A3(G301), .ZN(new_n908));
  AOI21_X1  g483(.A(G301), .B1(new_n906), .B2(new_n907), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n908), .A2(new_n834), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(G171), .B1(new_n537), .B2(new_n539), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n906), .A2(new_n907), .A3(G301), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n911), .A2(new_n912), .B1(new_n833), .B2(new_n832), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n870), .A2(KEYINPUT41), .A3(new_n879), .ZN(new_n914));
  OAI22_X1  g489(.A1(new_n910), .A2(new_n913), .B1(new_n914), .B2(new_n887), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n835), .A2(new_n912), .A3(new_n911), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n834), .B1(new_n908), .B2(new_n909), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n880), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(KEYINPUT104), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n890), .B(new_n920), .C1(new_n910), .C2(new_n913), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n919), .A2(new_n921), .A3(KEYINPUT105), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n896), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n896), .B1(new_n919), .B2(new_n921), .ZN(new_n927));
  XNOR2_X1  g502(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n926), .A2(new_n863), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n915), .ZN(new_n932));
  AND4_X1   g507(.A1(new_n882), .A2(new_n916), .A3(new_n883), .A4(new_n917), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n896), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n934), .A2(new_n863), .ZN(new_n935));
  INV_X1    g510(.A(new_n896), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n922), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(KEYINPUT107), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT107), .B1(new_n935), .B2(new_n937), .ZN(new_n940));
  OAI211_X1 g515(.A(KEYINPUT44), .B(new_n931), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n942));
  AND4_X1   g517(.A1(new_n863), .A2(new_n937), .A3(new_n934), .A4(new_n928), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n936), .B1(new_n922), .B2(new_n923), .ZN(new_n945));
  AOI211_X1 g520(.A(G37), .B(new_n927), .C1(new_n945), .C2(new_n925), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n944), .B1(new_n946), .B2(new_n928), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n942), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n926), .A2(new_n863), .A3(new_n937), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n943), .B1(new_n950), .B2(new_n929), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n951), .A2(KEYINPUT106), .A3(KEYINPUT44), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n941), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(KEYINPUT108), .B(new_n941), .C1(new_n949), .C2(new_n952), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(G397));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n843), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n468), .A2(G40), .A3(new_n474), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  OR3_X1    g538(.A1(new_n961), .A2(G1996), .A3(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT46), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n961), .A2(new_n963), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n746), .B(new_n749), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n968), .A2(new_n753), .A3(new_n757), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n965), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n970), .B(KEYINPUT126), .Z(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(KEYINPUT47), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n966), .A2(G1996), .A3(new_n758), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n973), .B(KEYINPUT109), .Z(new_n974));
  OAI21_X1  g549(.A(new_n968), .B1(G1996), .B2(new_n758), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n974), .B1(new_n966), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n717), .A2(new_n720), .ZN(new_n977));
  AOI22_X1  g552(.A1(new_n976), .A2(new_n977), .B1(new_n749), .B2(new_n747), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n967), .A2(G1986), .A3(G290), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT127), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT48), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n719), .B1(new_n712), .B2(new_n716), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n966), .B1(new_n977), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n976), .A2(new_n983), .ZN(new_n984));
  OAI22_X1  g559(.A1(new_n978), .A2(new_n967), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n972), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n495), .A2(new_n958), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n960), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n963), .B1(KEYINPUT110), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n960), .A2(G1384), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n843), .A2(new_n990), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n988), .A2(KEYINPUT110), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n989), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(KEYINPUT111), .B(G1971), .Z(new_n994));
  AND2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n987), .A2(KEYINPUT50), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n987), .A2(KEYINPUT50), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n962), .A3(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(G2090), .ZN(new_n999));
  OAI21_X1  g574(.A(G8), .B1(new_n995), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G303), .A2(G8), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1001), .B(KEYINPUT55), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n963), .A2(new_n987), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n697), .A2(G1976), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT52), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT112), .B1(new_n697), .B2(G1976), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1007), .B(new_n1010), .C1(KEYINPUT52), .C2(new_n1008), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT113), .B(G1981), .Z(new_n1015));
  NAND2_X1  g590(.A1(new_n594), .A2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g591(.A(KEYINPUT114), .B(G86), .Z(new_n1017));
  OAI21_X1  g592(.A(new_n591), .B1(new_n512), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n1020), .A2(new_n1021), .A3(new_n590), .ZN(new_n1022));
  INV_X1    g597(.A(G1981), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1016), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT49), .ZN(new_n1025));
  OR2_X1    g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(new_n1007), .A3(new_n1027), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1014), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1976), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1028), .A2(new_n1030), .A3(new_n697), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n1016), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n1004), .A2(new_n1029), .B1(new_n1007), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1014), .A2(new_n1034), .A3(new_n1028), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1003), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1029), .A2(new_n1034), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n495), .A2(new_n990), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n962), .A2(new_n988), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT117), .B(G2084), .ZN(new_n1043));
  OAI22_X1  g618(.A1(new_n1042), .A2(G1966), .B1(new_n998), .B2(new_n1043), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1044), .A2(G8), .A3(G168), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT63), .B1(new_n1039), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1003), .A2(KEYINPUT63), .A3(new_n1045), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1029), .A2(new_n1036), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1029), .A2(new_n1036), .A3(KEYINPUT118), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1047), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1033), .B1(new_n1046), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(G286), .A2(G8), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1054), .B(KEYINPUT122), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(G8), .B2(new_n1044), .ZN(new_n1056));
  XOR2_X1   g631(.A(new_n1056), .B(KEYINPUT51), .Z(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1044), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1058), .A2(KEYINPUT123), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(KEYINPUT123), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1057), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT62), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT62), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1057), .B(new_n1063), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n998), .B(KEYINPUT121), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n765), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n993), .B2(G2078), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(G2078), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1042), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1066), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1071), .A2(G171), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1062), .A2(new_n1064), .A3(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n993), .A2(G1996), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT58), .B(G1341), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1005), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n561), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1065), .A2(new_n800), .B1(new_n749), .B2(new_n1005), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1080), .A2(KEYINPUT60), .A3(new_n610), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT56), .B(G2072), .Z(new_n1084));
  INV_X1    g659(.A(new_n998), .ZN(new_n1085));
  OAI22_X1  g660(.A1(new_n993), .A2(new_n1084), .B1(G1956), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n574), .A2(KEYINPUT57), .A3(new_n579), .ZN(new_n1087));
  XOR2_X1   g662(.A(new_n1087), .B(KEYINPUT120), .Z(new_n1088));
  AND2_X1   g663(.A1(new_n872), .A2(KEYINPUT119), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n574), .B1(new_n872), .B2(KEYINPUT119), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1088), .B1(KEYINPUT57), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1086), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1086), .A2(new_n1093), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT61), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1094), .A2(KEYINPUT61), .A3(new_n1095), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1083), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n610), .B1(new_n1080), .B2(KEYINPUT60), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(KEYINPUT60), .B2(new_n1080), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1095), .B1(new_n1080), .B2(new_n610), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1098), .A2(new_n1100), .B1(new_n1101), .B2(new_n1094), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1103), .B1(new_n961), .B2(new_n962), .ZN(new_n1104));
  AOI211_X1 g679(.A(KEYINPUT124), .B(new_n963), .C1(new_n959), .C2(new_n960), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n991), .B(new_n1069), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(KEYINPUT125), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1108));
  XNOR2_X1  g683(.A(G301), .B(KEYINPUT54), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1107), .A2(new_n1110), .B1(new_n1071), .B2(new_n1109), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1061), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1073), .B1(new_n1102), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1053), .B1(new_n1113), .B2(new_n1039), .ZN(new_n1114));
  XOR2_X1   g689(.A(G290), .B(G1986), .Z(new_n1115));
  OAI211_X1 g690(.A(new_n976), .B(new_n983), .C1(new_n967), .C2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n986), .B1(new_n1114), .B2(new_n1116), .ZN(G329));
  assign    G231 = 1'b0;
  OR4_X1    g692(.A1(new_n461), .A2(G229), .A3(G401), .A4(G227), .ZN(new_n1119));
  NOR3_X1   g693(.A1(new_n865), .A2(new_n1119), .A3(new_n951), .ZN(G308));
  INV_X1    g694(.A(G308), .ZN(G225));
endmodule


