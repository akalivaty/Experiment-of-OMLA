//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT32), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT2), .B(G113), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT69), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT69), .A2(G119), .ZN(new_n194));
  INV_X1    g008(.A(G116), .ZN(new_n195));
  NOR3_X1   g009(.A1(new_n193), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G116), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n191), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  XOR2_X1   g013(.A(KEYINPUT2), .B(G113), .Z(new_n200));
  INV_X1    g014(.A(KEYINPUT69), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(new_n197), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(G116), .A3(new_n192), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n200), .B(new_n203), .C1(G116), .C2(new_n197), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n199), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G143), .B(G146), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT0), .A3(G128), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT0), .B(G128), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  INV_X1    g026(.A(G134), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT65), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G134), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G137), .ZN(new_n218));
  AOI21_X1  g032(.A(KEYINPUT11), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n214), .A2(new_n216), .A3(new_n220), .A4(G137), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT11), .ZN(new_n224));
  NOR3_X1   g038(.A1(new_n224), .A2(new_n213), .A3(G137), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n214), .A2(new_n216), .A3(G137), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(KEYINPUT66), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n212), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT65), .B(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n224), .B1(new_n229), .B2(G137), .ZN(new_n230));
  AND4_X1   g044(.A1(new_n212), .A2(new_n227), .A3(new_n221), .A4(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n211), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(G137), .B1(new_n214), .B2(new_n216), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n234), .B1(new_n213), .B2(G137), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n229), .B2(G137), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n235), .A2(new_n237), .A3(G131), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G143), .ZN(new_n241));
  INV_X1    g055(.A(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G146), .ZN(new_n243));
  AOI21_X1  g057(.A(G128), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(KEYINPUT1), .A3(G146), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT68), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n245), .B(new_n248), .C1(new_n207), .C2(G128), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n207), .A2(new_n251), .A3(G128), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n227), .A2(new_n212), .A3(new_n221), .A4(new_n230), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n239), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n232), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n206), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n232), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n226), .A2(KEYINPUT66), .ZN(new_n261));
  INV_X1    g075(.A(new_n225), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n221), .B1(new_n233), .B2(KEYINPUT11), .ZN(new_n264));
  OAI21_X1  g078(.A(G131), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n210), .B1(new_n265), .B2(new_n254), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT70), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n268));
  INV_X1    g082(.A(G128), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(KEYINPUT1), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n247), .A2(new_n249), .B1(new_n207), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(new_n238), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n268), .B1(new_n272), .B2(new_n254), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n260), .A2(new_n267), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n258), .A2(new_n274), .ZN(new_n275));
  XOR2_X1   g089(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n276));
  NOR2_X1   g090(.A1(G237), .A2(G953), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G210), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n276), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT26), .B(G101), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n265), .A2(new_n254), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT70), .B1(new_n283), .B2(new_n211), .ZN(new_n284));
  AOI211_X1 g098(.A(new_n259), .B(new_n210), .C1(new_n265), .C2(new_n254), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n231), .A2(new_n271), .A3(new_n238), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(new_n205), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n282), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT72), .B(KEYINPUT31), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n275), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT31), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(new_n275), .B2(new_n289), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT28), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n295), .B1(new_n256), .B2(new_n205), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n256), .A2(new_n205), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n288), .A2(new_n260), .A3(new_n267), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n296), .B(new_n297), .C1(new_n298), .C2(new_n295), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n282), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT73), .B1(new_n294), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n255), .A2(KEYINPUT30), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n302), .A2(new_n284), .A3(new_n285), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n257), .B1(new_n287), .B2(new_n266), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n205), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n298), .A2(new_n281), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT31), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n275), .A2(new_n289), .A3(new_n290), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n308), .A2(new_n300), .A3(KEYINPUT73), .A4(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n190), .B1(new_n301), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G902), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n284), .A2(new_n285), .A3(new_n287), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n298), .B1(new_n314), .B2(new_n206), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT28), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n316), .A2(KEYINPUT29), .A3(new_n296), .A4(new_n281), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n275), .A2(new_n298), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n282), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n299), .A2(new_n282), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n313), .B(new_n317), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G472), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n308), .A2(new_n300), .A3(new_n309), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n188), .B1(new_n327), .B2(new_n310), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n312), .B(new_n324), .C1(KEYINPUT32), .C2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT5), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n196), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n203), .B1(G116), .B2(new_n197), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n331), .B(G113), .C1(new_n332), .C2(new_n330), .ZN(new_n333));
  INV_X1    g147(.A(G104), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT3), .B1(new_n334), .B2(G107), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n336));
  INV_X1    g150(.A(G107), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(G104), .ZN(new_n338));
  INV_X1    g152(.A(G101), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n334), .A2(G107), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n335), .A2(new_n338), .A3(new_n339), .A4(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n334), .A2(G107), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n337), .A2(G104), .ZN(new_n343));
  OAI21_X1  g157(.A(G101), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n333), .A2(new_n204), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n335), .A2(new_n338), .A3(new_n340), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n335), .A2(new_n338), .A3(KEYINPUT79), .A4(new_n340), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(G101), .A3(new_n351), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n341), .A2(KEYINPUT4), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n339), .A2(KEYINPUT4), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n350), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n205), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n347), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G110), .B(G122), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n347), .B(new_n359), .C1(new_n354), .C2(new_n357), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(KEYINPUT6), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n210), .A2(G125), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n364), .B1(new_n253), .B2(G125), .ZN(new_n365));
  INV_X1    g179(.A(G224), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(G953), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n365), .B(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT6), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n358), .A2(new_n369), .A3(new_n360), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n363), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT84), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n363), .A2(new_n368), .A3(KEYINPUT84), .A4(new_n370), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT7), .ZN(new_n376));
  OR3_X1    g190(.A1(new_n365), .A2(new_n376), .A3(new_n367), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n359), .B(KEYINPUT8), .ZN(new_n378));
  INV_X1    g192(.A(new_n347), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n346), .B1(new_n333), .B2(new_n204), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n365), .B1(new_n376), .B2(new_n367), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n377), .A2(new_n381), .A3(new_n362), .A4(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n313), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n375), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(G210), .B1(G237), .B2(G902), .ZN(new_n387));
  XOR2_X1   g201(.A(new_n387), .B(KEYINPUT85), .Z(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n384), .B1(new_n373), .B2(new_n374), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n387), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(G214), .B1(G237), .B2(G902), .ZN(new_n393));
  XOR2_X1   g207(.A(new_n393), .B(KEYINPUT82), .Z(new_n394));
  XOR2_X1   g208(.A(new_n394), .B(KEYINPUT83), .Z(new_n395));
  INV_X1    g209(.A(G952), .ZN(new_n396));
  AOI211_X1 g210(.A(G953), .B(new_n396), .C1(G234), .C2(G237), .ZN(new_n397));
  INV_X1    g211(.A(G953), .ZN(new_n398));
  AOI211_X1 g212(.A(new_n313), .B(new_n398), .C1(G234), .C2(G237), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT21), .B(G898), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n395), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n392), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G475), .ZN(new_n404));
  INV_X1    g218(.A(G140), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G125), .ZN(new_n406));
  INV_X1    g220(.A(G125), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G140), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n408), .A3(KEYINPUT76), .ZN(new_n409));
  OR3_X1    g223(.A1(new_n405), .A2(KEYINPUT76), .A3(G125), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT16), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT16), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n406), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n240), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n240), .B1(new_n411), .B2(new_n413), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n242), .A2(KEYINPUT86), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n242), .A2(KEYINPUT86), .ZN(new_n419));
  OAI211_X1 g233(.A(G214), .B(new_n277), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G237), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(new_n398), .A3(G214), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(KEYINPUT86), .B2(new_n242), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n212), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT17), .ZN(new_n425));
  INV_X1    g239(.A(new_n424), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT86), .B(G143), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n423), .B(new_n212), .C1(new_n422), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n417), .B(new_n425), .C1(KEYINPUT17), .C2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n423), .B1(new_n422), .B2(new_n427), .ZN(new_n431));
  AND2_X1   g245(.A1(KEYINPUT18), .A2(G131), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT87), .ZN(new_n434));
  XNOR2_X1  g248(.A(G125), .B(G140), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n240), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n409), .A2(new_n410), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n434), .B(new_n436), .C1(new_n437), .C2(new_n240), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT87), .A4(G146), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n433), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n430), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G113), .B(G122), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT90), .B(G104), .ZN(new_n445));
  XOR2_X1   g259(.A(new_n444), .B(new_n445), .Z(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(KEYINPUT91), .ZN(new_n447));
  AOI21_X1  g261(.A(G902), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n442), .B1(KEYINPUT91), .B2(new_n446), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n404), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n437), .A2(KEYINPUT19), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n435), .A2(KEYINPUT19), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(G146), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT88), .B1(new_n454), .B2(new_n416), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n411), .A2(new_n413), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G146), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT88), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT19), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(new_n409), .B2(new_n410), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n240), .B1(new_n460), .B2(new_n452), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n455), .A2(new_n429), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n441), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT89), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n446), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n433), .A2(new_n440), .ZN(new_n467));
  INV_X1    g281(.A(new_n428), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(new_n424), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n457), .A2(new_n461), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(KEYINPUT88), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n467), .B1(new_n471), .B2(new_n462), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT89), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n466), .A2(new_n473), .B1(new_n446), .B2(new_n443), .ZN(new_n474));
  NOR2_X1   g288(.A1(G475), .A2(G902), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT20), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n443), .A2(new_n446), .ZN(new_n478));
  INV_X1    g292(.A(new_n446), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(new_n472), .B2(KEYINPUT89), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n464), .A2(new_n465), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT20), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n475), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n450), .B1(new_n477), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G469), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n352), .A2(new_n353), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n211), .A3(new_n356), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT10), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n345), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n244), .A2(new_n246), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n252), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n346), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n253), .A2(new_n490), .B1(new_n493), .B2(new_n489), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n283), .A2(KEYINPUT80), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT80), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n496), .B1(new_n265), .B2(new_n254), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n488), .B(new_n494), .C1(new_n495), .C2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT12), .ZN(new_n499));
  OR2_X1    g313(.A1(new_n499), .A2(KEYINPUT81), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(KEYINPUT81), .ZN(new_n501));
  INV_X1    g315(.A(new_n283), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n345), .B1(new_n252), .B2(new_n491), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(new_n271), .B2(new_n345), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n500), .B(new_n501), .C1(new_n502), .C2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n493), .B1(new_n253), .B2(new_n346), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n506), .A2(KEYINPUT81), .A3(new_n499), .A4(new_n283), .ZN(new_n507));
  XNOR2_X1  g321(.A(G110), .B(G140), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n398), .A2(G227), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n498), .A2(new_n505), .A3(new_n507), .A4(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n494), .A2(new_n488), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n283), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n511), .B1(new_n515), .B2(new_n498), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n486), .B(new_n313), .C1(new_n513), .C2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n486), .A2(new_n313), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n498), .A2(new_n507), .A3(new_n505), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n510), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n515), .A2(new_n498), .A3(new_n511), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n517), .B(new_n519), .C1(new_n486), .C2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT92), .B1(new_n242), .B2(G128), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT92), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n269), .A3(G143), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n242), .A2(G128), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n229), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT93), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT13), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n242), .A2(KEYINPUT13), .A3(G128), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n528), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G134), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT93), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n528), .A2(new_n537), .A3(new_n229), .A4(new_n529), .ZN(new_n538));
  INV_X1    g352(.A(G122), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G116), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n195), .A2(G122), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G107), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n540), .A2(new_n541), .A3(new_n337), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n531), .A2(new_n536), .A3(new_n538), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT94), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n535), .A2(G134), .B1(new_n543), .B2(new_n544), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT94), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n548), .A2(new_n549), .A3(new_n538), .A4(new_n531), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n528), .A2(new_n529), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n217), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n553), .A2(new_n530), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n337), .B1(new_n540), .B2(KEYINPUT14), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(new_n542), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT9), .B(G234), .ZN(new_n560));
  INV_X1    g374(.A(G217), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n560), .A2(new_n561), .A3(G953), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n557), .B1(new_n547), .B2(new_n550), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n562), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n313), .ZN(new_n568));
  INV_X1    g382(.A(G478), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n569), .A2(KEYINPUT15), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n567), .B(new_n313), .C1(KEYINPUT15), .C2(new_n569), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(G221), .B1(new_n560), .B2(G902), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n485), .A2(new_n524), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n403), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n197), .A2(G128), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT23), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n202), .A2(G128), .A3(new_n192), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(KEYINPUT74), .A3(KEYINPUT23), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n202), .A2(new_n192), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n269), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT74), .B1(new_n580), .B2(KEYINPUT23), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n579), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n582), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n578), .B1(new_n587), .B2(G128), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT24), .B(G110), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OAI22_X1  g404(.A1(new_n586), .A2(G110), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n591), .A2(new_n457), .A3(new_n436), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n590), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n415), .B2(new_n416), .ZN(new_n594));
  INV_X1    g408(.A(G110), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT75), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n595), .B1(new_n586), .B2(new_n596), .ZN(new_n597));
  OAI211_X1 g411(.A(KEYINPUT75), .B(new_n579), .C1(new_n584), .C2(new_n585), .ZN(new_n598));
  AOI211_X1 g412(.A(KEYINPUT77), .B(new_n594), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT77), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n586), .A2(new_n596), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(new_n598), .A3(G110), .ZN(new_n602));
  INV_X1    g416(.A(new_n594), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n592), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT22), .B(G137), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n398), .A2(G221), .A3(G234), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n606), .B(new_n607), .Z(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n592), .B(new_n608), .C1(new_n599), .C2(new_n604), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n561), .B1(G234), .B2(new_n313), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(G902), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT78), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n610), .A2(new_n313), .A3(new_n611), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT25), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n610), .A2(KEYINPUT25), .A3(new_n313), .A4(new_n611), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n617), .B1(new_n622), .B2(new_n613), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n329), .A2(new_n577), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  NAND2_X1  g439(.A1(new_n327), .A2(new_n310), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n313), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n328), .B1(new_n627), .B2(G472), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n524), .A2(new_n575), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n623), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT95), .ZN(new_n633));
  INV_X1    g447(.A(new_n387), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n386), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT95), .B1(new_n390), .B2(new_n387), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n391), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n394), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n401), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT98), .B(G478), .Z(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n567), .B2(new_n313), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT33), .B1(new_n565), .B2(KEYINPUT96), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n565), .A2(new_n562), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n565), .A2(new_n562), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT96), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n559), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n564), .A2(new_n648), .A3(KEYINPUT33), .A4(new_n566), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n569), .A2(G902), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT97), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n646), .A2(new_n649), .A3(new_n653), .A4(new_n650), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n642), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n485), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n639), .A2(new_n640), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n632), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT99), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT34), .B(G104), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  INV_X1    g475(.A(new_n450), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n474), .A2(KEYINPUT20), .A3(new_n476), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n483), .B1(new_n482), .B2(new_n475), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n573), .B(new_n662), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n401), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n666), .A2(new_n638), .A3(new_n637), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n628), .A3(new_n631), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT35), .B(G107), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G9));
  OAI21_X1  g484(.A(new_n605), .B1(KEYINPUT36), .B2(new_n609), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n609), .A2(KEYINPUT36), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n592), .B(new_n672), .C1(new_n599), .C2(new_n604), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  AOI22_X1  g489(.A1(new_n622), .A2(new_n613), .B1(new_n615), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n628), .A2(new_n577), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  XOR2_X1   g494(.A(new_n397), .B(KEYINPUT100), .Z(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(G900), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n682), .B1(new_n683), .B2(new_n399), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n485), .A2(new_n573), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n676), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n329), .A2(new_n639), .A3(new_n687), .A4(new_n630), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n626), .A2(new_n187), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n189), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n626), .A2(new_n190), .B1(new_n323), .B2(G472), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n629), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n694), .A2(KEYINPUT101), .A3(new_n639), .A4(new_n687), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G128), .ZN(G30));
  XOR2_X1   g511(.A(new_n684), .B(KEYINPUT39), .Z(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n629), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT40), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n485), .A2(new_n574), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n676), .A2(new_n638), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n392), .B(KEYINPUT38), .ZN(new_n704));
  INV_X1    g518(.A(G472), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n275), .A2(new_n289), .ZN(new_n706));
  INV_X1    g520(.A(new_n315), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n706), .B1(new_n707), .B2(new_n281), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n705), .B1(new_n708), .B2(new_n313), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n709), .B1(new_n626), .B2(new_n190), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n692), .A2(new_n710), .ZN(new_n711));
  AND4_X1   g525(.A1(new_n701), .A2(new_n703), .A3(new_n704), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n242), .ZN(G45));
  OAI21_X1  g527(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n652), .A2(new_n654), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n714), .B(new_n685), .C1(new_n715), .C2(new_n642), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n676), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(new_n329), .A3(new_n630), .A4(new_n639), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  AND2_X1   g533(.A1(new_n515), .A2(new_n498), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n512), .B1(new_n720), .B2(new_n511), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n313), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(G469), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n723), .A2(new_n575), .A3(new_n517), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n329), .A2(new_n623), .A3(new_n724), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n725), .A2(new_n657), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NAND4_X1  g542(.A1(new_n667), .A2(new_n329), .A3(new_n623), .A4(new_n724), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  AND3_X1   g544(.A1(new_n637), .A2(new_n638), .A3(new_n724), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n485), .A2(new_n574), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n676), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n329), .A2(new_n731), .A3(new_n640), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G119), .ZN(G21));
  NAND3_X1  g549(.A1(new_n637), .A2(new_n702), .A3(new_n638), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n316), .A2(new_n296), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n282), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n188), .B1(new_n739), .B2(new_n294), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(new_n627), .B2(G472), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n724), .A2(new_n640), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n737), .A2(new_n741), .A3(new_n743), .A4(new_n623), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G122), .ZN(G24));
  INV_X1    g559(.A(new_n716), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n731), .A2(new_n741), .A3(new_n677), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G125), .ZN(G27));
  NAND3_X1  g562(.A1(new_n389), .A2(new_n391), .A3(new_n638), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n521), .A2(KEYINPUT102), .A3(G469), .A4(new_n522), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n517), .A2(new_n750), .A3(new_n519), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n498), .A2(new_n511), .ZN(new_n752));
  AOI22_X1  g566(.A1(new_n752), .A2(new_n515), .B1(new_n520), .B2(new_n510), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT102), .B1(new_n753), .B2(G469), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n575), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n749), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n329), .A2(new_n623), .A3(new_n746), .A4(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT42), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n691), .A2(KEYINPUT103), .A3(new_n189), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT103), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n761), .B1(new_n328), .B2(KEYINPUT32), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n693), .A3(new_n762), .ZN(new_n763));
  NOR4_X1   g577(.A1(new_n716), .A2(new_n749), .A3(new_n758), .A4(new_n755), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n764), .A3(new_n623), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n759), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  INV_X1    g581(.A(new_n686), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n329), .A2(new_n623), .A3(new_n768), .A4(new_n756), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  OAI21_X1  g584(.A(G469), .B1(new_n753), .B2(KEYINPUT45), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n521), .A2(KEYINPUT45), .A3(new_n522), .ZN(new_n772));
  OR3_X1    g586(.A1(new_n771), .A2(new_n772), .A3(KEYINPUT104), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT104), .B1(new_n771), .B2(new_n772), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n518), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n775), .A2(KEYINPUT46), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n517), .B1(new_n775), .B2(KEYINPUT46), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n575), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n778), .A2(new_n699), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n655), .A2(new_n714), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT43), .ZN(new_n782));
  AOI21_X1  g596(.A(G902), .B1(new_n327), .B2(new_n310), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n691), .B1(new_n705), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(new_n784), .A3(new_n677), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT44), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n749), .B(KEYINPUT105), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n780), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  XNOR2_X1  g603(.A(new_n778), .B(KEYINPUT47), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  NOR4_X1   g605(.A1(new_n329), .A2(new_n623), .A3(new_n716), .A4(new_n749), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  NOR2_X1   g608(.A1(G952), .A2(G953), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n729), .A2(new_n734), .ZN(new_n796));
  INV_X1    g610(.A(new_n740), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n623), .B(new_n797), .C1(new_n705), .C2(new_n783), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n798), .A2(new_n736), .A3(new_n742), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n665), .B1(new_n655), .B2(new_n485), .ZN(new_n800));
  INV_X1    g614(.A(new_n402), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n801), .B1(new_n389), .B2(new_n391), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n623), .A2(new_n630), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n784), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n799), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n624), .A2(new_n678), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n796), .A2(new_n726), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n749), .A2(new_n684), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n329), .A2(new_n630), .A3(new_n733), .A4(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n741), .A2(new_n677), .A3(new_n746), .A4(new_n756), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n769), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n766), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT107), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n769), .A2(new_n810), .A3(new_n811), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n765), .B2(new_n759), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n628), .A2(new_n631), .A3(new_n802), .A4(new_n800), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n729), .A2(new_n734), .A3(new_n744), .A4(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n678), .B(new_n624), .C1(new_n725), .C2(new_n657), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT107), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n816), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n718), .A2(new_n747), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n684), .B(KEYINPUT108), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n677), .A2(new_n755), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n711), .A3(new_n737), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n696), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n696), .A2(KEYINPUT52), .A3(new_n823), .A4(new_n826), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n814), .A2(new_n822), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT53), .ZN(new_n832));
  XOR2_X1   g646(.A(KEYINPUT109), .B(KEYINPUT54), .Z(new_n833));
  NAND3_X1  g647(.A1(new_n816), .A2(new_n820), .A3(KEYINPUT53), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n829), .B2(new_n830), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n829), .A2(new_n830), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n808), .A2(new_n813), .A3(KEYINPUT107), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n821), .B1(new_n816), .B2(new_n820), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n835), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n832), .A2(KEYINPUT54), .B1(new_n833), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n782), .A2(new_n682), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n724), .A2(new_n389), .A3(new_n391), .A4(new_n638), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n763), .A2(new_n623), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g661(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n845), .A2(KEYINPUT110), .A3(KEYINPUT48), .A4(new_n846), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n843), .A2(new_n798), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n731), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n623), .A2(new_n397), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n711), .A2(new_n844), .A3(new_n853), .ZN(new_n854));
  AOI211_X1 g668(.A(new_n396), .B(G953), .C1(new_n854), .C2(new_n656), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n849), .A2(new_n850), .A3(new_n852), .A4(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT111), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n851), .A2(new_n787), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n723), .A2(new_n517), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT106), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n575), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n858), .B1(new_n790), .B2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n741), .A2(new_n677), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n655), .A2(new_n485), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n845), .A2(new_n864), .B1(new_n854), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n704), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n867), .A2(new_n394), .A3(new_n724), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n851), .A2(KEYINPUT50), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT50), .B1(new_n851), .B2(new_n868), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n872));
  OR3_X1    g686(.A1(new_n863), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n872), .B1(new_n863), .B2(new_n871), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n857), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n795), .B1(new_n842), .B2(new_n875), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n860), .B(KEYINPUT49), .Z(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(new_n692), .A3(new_n867), .A4(new_n710), .ZN(new_n878));
  INV_X1    g692(.A(new_n623), .ZN(new_n879));
  INV_X1    g693(.A(new_n395), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n781), .A2(new_n880), .A3(new_n575), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT112), .B1(new_n876), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n839), .A2(new_n840), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n831), .A2(KEYINPUT53), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT54), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n841), .A2(new_n833), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n875), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(G952), .B2(G953), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT112), .ZN(new_n890));
  INV_X1    g704(.A(new_n882), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n883), .A2(new_n892), .ZN(G75));
  NAND2_X1  g707(.A1(new_n363), .A2(new_n370), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(new_n368), .Z(new_n895));
  XNOR2_X1  g709(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n895), .B(new_n896), .ZN(new_n897));
  XNOR2_X1  g711(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n834), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n836), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(new_n831), .B2(KEYINPUT53), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n902), .A2(G902), .A3(new_n388), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT115), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n903), .A2(new_n904), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n899), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n398), .A2(G952), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT114), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n902), .A2(G210), .A3(G902), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT56), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n911), .B1(new_n914), .B2(new_n897), .ZN(new_n915));
  INV_X1    g729(.A(new_n897), .ZN(new_n916));
  AOI211_X1 g730(.A(KEYINPUT114), .B(new_n916), .C1(new_n912), .C2(new_n913), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n910), .A2(new_n918), .ZN(G51));
  XNOR2_X1  g733(.A(new_n841), .B(new_n833), .ZN(new_n920));
  XNOR2_X1  g734(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n518), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n721), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n902), .A2(G902), .A3(new_n773), .A4(new_n774), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT118), .Z(new_n926));
  AOI21_X1  g740(.A(new_n908), .B1(new_n924), .B2(new_n926), .ZN(G54));
  AND4_X1   g741(.A1(KEYINPUT58), .A2(new_n902), .A3(G475), .A4(G902), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n909), .B1(new_n928), .B2(new_n482), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(new_n482), .B2(new_n928), .ZN(G60));
  AND2_X1   g744(.A1(new_n646), .A2(new_n649), .ZN(new_n931));
  NAND2_X1  g745(.A1(G478), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT59), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n920), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n886), .A2(new_n887), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n931), .B1(new_n935), .B2(new_n933), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n934), .A2(new_n908), .A3(new_n936), .ZN(G63));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n938));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT60), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n938), .B1(new_n841), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n940), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n902), .A2(KEYINPUT119), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n908), .B1(new_n944), .B2(new_n675), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n941), .A2(new_n612), .A3(new_n943), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT120), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n941), .A2(KEYINPUT120), .A3(new_n612), .A4(new_n943), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n945), .A2(new_n948), .A3(KEYINPUT61), .A4(new_n949), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n902), .A2(KEYINPUT119), .A3(new_n942), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT119), .B1(new_n902), .B2(new_n942), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n675), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n953), .A2(new_n909), .A3(new_n946), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n950), .A2(new_n956), .ZN(G66));
  OAI21_X1  g771(.A(G953), .B1(new_n400), .B2(new_n366), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT121), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n820), .B2(G953), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n894), .B1(G898), .B2(new_n398), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(G69));
  NAND3_X1  g776(.A1(new_n788), .A2(new_n766), .A3(new_n769), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n780), .A2(new_n737), .A3(new_n846), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n964), .A2(new_n696), .A3(new_n823), .ZN(new_n965));
  AOI211_X1 g779(.A(new_n963), .B(new_n965), .C1(new_n791), .C2(new_n792), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n398), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n274), .A2(new_n304), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n460), .A2(new_n452), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(new_n970));
  XNOR2_X1  g784(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(G900), .B2(G953), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n967), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n975));
  INV_X1    g789(.A(new_n712), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(new_n696), .A3(new_n823), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT62), .Z(new_n978));
  NOR3_X1   g792(.A1(new_n749), .A2(new_n629), .A3(new_n699), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n329), .A2(new_n623), .A3(new_n800), .A4(new_n979), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT124), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n788), .A2(new_n978), .A3(new_n793), .A4(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n972), .B1(new_n982), .B2(G953), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n974), .A2(new_n975), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n398), .B1(G227), .B2(G900), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n985), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n974), .A2(new_n975), .A3(new_n987), .A4(new_n983), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n986), .A2(new_n988), .ZN(G72));
  XOR2_X1   g803(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n990));
  NOR2_X1   g804(.A1(new_n705), .A2(new_n313), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(new_n982), .B2(new_n820), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n318), .B(KEYINPUT127), .Z(new_n994));
  NOR3_X1   g808(.A1(new_n993), .A2(new_n282), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n992), .B1(new_n966), .B2(new_n820), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n282), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n909), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n992), .B1(new_n319), .B2(new_n706), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n832), .A2(new_n999), .ZN(new_n1000));
  NOR3_X1   g814(.A1(new_n995), .A2(new_n998), .A3(new_n1000), .ZN(G57));
endmodule


