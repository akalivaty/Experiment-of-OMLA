//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n795, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT90), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT14), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n208), .B(new_n209), .C1(G29gat), .C2(G36gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G29gat), .ZN(new_n213));
  INV_X1    g012(.A(G36gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT90), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n214), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n209), .B1(new_n216), .B2(new_n208), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n212), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219));
  INV_X1    g018(.A(G50gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT91), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT91), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G50gat), .ZN(new_n223));
  AOI21_X1  g022(.A(G43gat), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G43gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(G50gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n219), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n220), .A2(G43gat), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT89), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G43gat), .B(G50gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT89), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n219), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n218), .A2(new_n227), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n220), .A2(G43gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n225), .A2(G50gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(new_n235), .A3(new_n231), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n229), .A2(KEYINPUT15), .A3(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n208), .B1(G29gat), .B2(G36gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n215), .A2(new_n238), .A3(KEYINPUT14), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(new_n211), .A3(new_n210), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n233), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G8gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(G15gat), .B(G22gat), .ZN(new_n244));
  INV_X1    g043(.A(G1gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT16), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n244), .A2(G1gat), .ZN(new_n248));
  OAI211_X1 g047(.A(KEYINPUT92), .B(new_n243), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n244), .A2(G1gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n244), .A2(new_n246), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n243), .A2(KEYINPUT92), .ZN(new_n252));
  OR2_X1    g051(.A1(new_n243), .A2(KEYINPUT92), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n250), .A2(new_n251), .A3(new_n252), .A4(new_n253), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n242), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G229gat), .A2(G233gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT17), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n233), .B2(new_n241), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n222), .A2(G50gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n220), .A2(KEYINPUT91), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n225), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT15), .B1(new_n264), .B2(new_n234), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n237), .B1(new_n265), .B2(new_n240), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n218), .A2(new_n229), .A3(new_n232), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(KEYINPUT17), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n261), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n255), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT93), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT93), .ZN(new_n272));
  AOI211_X1 g071(.A(new_n272), .B(new_n255), .C1(new_n261), .C2(new_n268), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n259), .B(KEYINPUT18), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n242), .B(new_n255), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n257), .B(KEYINPUT13), .Z(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n233), .A2(new_n260), .A3(new_n241), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT17), .B1(new_n266), .B2(new_n267), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n270), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n272), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n269), .A2(KEYINPUT93), .A3(new_n270), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT18), .B1(new_n284), .B2(new_n259), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n207), .B1(new_n278), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n258), .B1(new_n282), .B2(new_n283), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT94), .B1(new_n287), .B2(KEYINPUT18), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n259), .B1(new_n271), .B2(new_n273), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT94), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT18), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n274), .A2(new_n277), .A3(new_n206), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n286), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT95), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n274), .A2(new_n277), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n297), .A2(new_n288), .A3(new_n206), .A4(new_n292), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT95), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(new_n286), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT85), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT3), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT22), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT72), .B(G218gat), .ZN(new_n305));
  INV_X1    g104(.A(G211gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n308));
  XNOR2_X1  g107(.A(G197gat), .B(G204gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT73), .B(G211gat), .ZN(new_n312));
  INV_X1    g111(.A(G218gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n307), .A2(new_n309), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(new_n308), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n310), .A2(new_n314), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n303), .B1(new_n320), .B2(KEYINPUT29), .ZN(new_n321));
  INV_X1    g120(.A(G141gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G148gat), .ZN(new_n323));
  INV_X1    g122(.A(G148gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G141gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n323), .A2(new_n325), .B1(KEYINPUT2), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G155gat), .ZN(new_n328));
  INV_X1    g127(.A(G162gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n326), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT81), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT81), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n327), .A2(new_n334), .A3(new_n331), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n330), .B(KEYINPUT80), .ZN(new_n336));
  INV_X1    g135(.A(new_n326), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n327), .A2(new_n337), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n333), .A2(new_n335), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(new_n336), .ZN(new_n342));
  INV_X1    g141(.A(new_n335), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n334), .B1(new_n327), .B2(new_n331), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT82), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n321), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n345), .A2(KEYINPUT3), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT77), .B(KEYINPUT29), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n320), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT84), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(G228gat), .ZN(new_n356));
  INV_X1    g155(.A(G233gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n320), .B(KEYINPUT84), .C1(new_n350), .C2(new_n352), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n349), .A2(new_n355), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n353), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n316), .B(new_n351), .C1(new_n318), .C2(new_n319), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n339), .B1(new_n362), .B2(new_n303), .ZN(new_n363));
  OAI22_X1  g162(.A1(new_n361), .A2(new_n363), .B1(new_n356), .B2(new_n357), .ZN(new_n364));
  INV_X1    g163(.A(G22gat), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n360), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n365), .B1(new_n360), .B2(new_n364), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n302), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n360), .A2(new_n364), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G22gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n360), .A2(new_n364), .A3(new_n365), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(KEYINPUT85), .A3(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G78gat), .B(G106gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT31), .B(G50gat), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n373), .B(new_n374), .Z(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n368), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n366), .A2(new_n367), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n378), .A2(KEYINPUT85), .A3(new_n375), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(G190gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT27), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G183gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT67), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT27), .B(G183gat), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n381), .B(new_n385), .C1(new_n386), .C2(new_n384), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT68), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT28), .ZN(new_n390));
  AOI21_X1  g189(.A(G190gat), .B1(new_n383), .B2(new_n384), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n391), .B(KEYINPUT68), .C1(new_n384), .C2(new_n386), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n386), .A2(KEYINPUT28), .A3(new_n381), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n396), .A2(KEYINPUT26), .ZN(new_n397));
  INV_X1    g196(.A(G169gat), .ZN(new_n398));
  INV_X1    g197(.A(G176gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n396), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n395), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT76), .ZN(new_n406));
  INV_X1    g205(.A(new_n396), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT23), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n407), .B1(new_n400), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(new_n408), .B2(new_n407), .ZN(new_n410));
  NAND3_X1  g209(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(G183gat), .B2(G190gat), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT66), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT24), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n413), .A2(new_n414), .B1(G183gat), .B2(G190gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n412), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT25), .B1(new_n410), .B2(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(KEYINPUT65), .B(G169gat), .Z(new_n419));
  NAND3_X1  g218(.A1(new_n419), .A2(KEYINPUT23), .A3(new_n399), .ZN(new_n420));
  INV_X1    g219(.A(G183gat), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n414), .B1(new_n421), .B2(new_n381), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n381), .A3(KEYINPUT64), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT64), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n424), .B1(G183gat), .B2(G190gat), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n422), .A2(new_n411), .A3(new_n423), .A4(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT25), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n420), .A2(new_n426), .A3(new_n427), .A4(new_n409), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n418), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n405), .A2(new_n406), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G226gat), .A2(G233gat), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n432), .B(KEYINPUT75), .Z(new_n433));
  AOI21_X1  g232(.A(new_n403), .B1(new_n393), .B2(new_n394), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT76), .B1(new_n434), .B2(new_n429), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n431), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n320), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n434), .A2(new_n429), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n432), .B1(new_n438), .B2(KEYINPUT29), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n438), .A2(new_n432), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n431), .A2(new_n435), .A3(new_n351), .ZN(new_n442));
  INV_X1    g241(.A(new_n433), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n440), .B1(new_n444), .B2(new_n437), .ZN(new_n445));
  XOR2_X1   g244(.A(G8gat), .B(G36gat), .Z(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(KEYINPUT78), .ZN(new_n447));
  XNOR2_X1  g246(.A(G64gat), .B(G92gat), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n447), .B(new_n448), .Z(new_n449));
  NAND2_X1  g248(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT79), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n445), .A2(KEYINPUT79), .A3(new_n449), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n442), .A2(new_n443), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n320), .B1(new_n455), .B2(new_n441), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT30), .ZN(new_n457));
  INV_X1    g256(.A(new_n449), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n456), .A2(new_n457), .A3(new_n458), .A4(new_n440), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n458), .B(new_n440), .C1(new_n444), .C2(new_n437), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT30), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n454), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G1gat), .B(G29gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(KEYINPUT0), .ZN(new_n465));
  XNOR2_X1  g264(.A(G57gat), .B(G85gat), .ZN(new_n466));
  XOR2_X1   g265(.A(new_n465), .B(new_n466), .Z(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(G225gat), .A2(G233gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(G113gat), .B(G120gat), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n470), .A2(KEYINPUT1), .ZN(new_n471));
  XOR2_X1   g270(.A(G127gat), .B(G134gat), .Z(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n350), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n341), .A2(new_n346), .A3(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n339), .A2(KEYINPUT4), .A3(new_n473), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT4), .B1(new_n339), .B2(new_n473), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n469), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT39), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n468), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OR2_X1    g281(.A1(new_n480), .A2(new_n481), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n339), .A2(new_n473), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n469), .B(new_n484), .C1(new_n347), .C2(new_n473), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(KEYINPUT86), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n482), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT40), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n476), .A2(new_n479), .A3(KEYINPUT5), .A4(new_n469), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n476), .A2(new_n469), .A3(new_n479), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT5), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n484), .B1(new_n347), .B2(new_n473), .ZN(new_n493));
  INV_X1    g292(.A(new_n469), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n490), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT87), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(KEYINPUT87), .B(new_n490), .C1(new_n491), .C2(new_n495), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n468), .A3(new_n499), .ZN(new_n500));
  OAI211_X1 g299(.A(KEYINPUT40), .B(new_n482), .C1(new_n483), .C2(new_n486), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n489), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n380), .B1(new_n463), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n445), .A2(KEYINPUT37), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT37), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n505), .B(new_n440), .C1(new_n444), .C2(new_n437), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n449), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT38), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT88), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n468), .B(new_n490), .C1(new_n491), .C2(new_n495), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n467), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT83), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n496), .A2(KEYINPUT83), .A3(new_n467), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n500), .A2(new_n516), .A3(new_n511), .A4(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n460), .ZN(new_n519));
  INV_X1    g318(.A(new_n507), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n437), .B1(new_n455), .B2(new_n441), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n436), .A2(new_n320), .A3(new_n439), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n522), .A2(KEYINPUT37), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT38), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n519), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n509), .A2(new_n513), .A3(new_n518), .A4(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT88), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n527), .B(KEYINPUT38), .C1(new_n504), .C2(new_n507), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n503), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n405), .A2(new_n430), .A3(new_n473), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT69), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT69), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n438), .A2(new_n533), .A3(new_n473), .ZN(new_n534));
  NAND2_X1  g333(.A1(G227gat), .A2(G233gat), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n471), .B(new_n472), .Z(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(new_n434), .B2(new_n429), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n532), .A2(new_n534), .A3(new_n535), .A4(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT34), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT32), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n532), .A2(new_n534), .A3(new_n537), .ZN(new_n541));
  INV_X1    g340(.A(new_n535), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT33), .B1(new_n541), .B2(new_n542), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT70), .B(G71gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(G99gat), .ZN(new_n546));
  XOR2_X1   g345(.A(G15gat), .B(G43gat), .Z(new_n547));
  XOR2_X1   g346(.A(new_n546), .B(new_n547), .Z(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NOR3_X1   g348(.A1(new_n543), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  AOI221_X4 g349(.A(new_n540), .B1(KEYINPUT33), .B2(new_n548), .C1(new_n541), .C2(new_n542), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n539), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n544), .A2(new_n549), .ZN(new_n553));
  INV_X1    g352(.A(new_n543), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n539), .ZN(new_n556));
  INV_X1    g355(.A(new_n551), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(KEYINPUT36), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n552), .A2(KEYINPUT71), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n555), .A2(new_n557), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT71), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n563), .A3(new_n539), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n561), .A2(new_n564), .A3(new_n558), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n560), .B1(KEYINPUT36), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n452), .A2(new_n453), .B1(new_n459), .B2(new_n461), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n517), .A2(new_n511), .ZN(new_n568));
  INV_X1    g367(.A(new_n510), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT83), .B1(new_n496), .B2(new_n467), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n567), .B1(new_n571), .B2(new_n512), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n380), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n530), .A2(new_n566), .A3(new_n573), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n518), .A2(new_n513), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n377), .A2(new_n552), .A3(new_n558), .A4(new_n379), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT35), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n567), .A2(new_n577), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n558), .B1(new_n552), .B2(KEYINPUT71), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n563), .B1(new_n562), .B2(new_n539), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR4_X1   g381(.A1(new_n366), .A2(new_n367), .A3(new_n302), .A4(new_n376), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n375), .B1(new_n378), .B2(KEYINPUT85), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n583), .B1(new_n584), .B2(new_n368), .ZN(new_n585));
  INV_X1    g384(.A(new_n571), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(new_n513), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n582), .A2(new_n585), .A3(new_n567), .A4(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n579), .B1(new_n588), .B2(KEYINPUT35), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n301), .B1(new_n574), .B2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(KEYINPUT41), .ZN(new_n592));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT8), .ZN(new_n598));
  NAND2_X1  g397(.A1(G85gat), .A2(G92gat), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT7), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(G85gat), .ZN(new_n602));
  INV_X1    g401(.A(G92gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n598), .A2(new_n601), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G99gat), .B(G106gat), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  AND3_X1   g408(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g411(.A1(KEYINPUT8), .A2(new_n597), .B1(new_n602), .B2(new_n603), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n607), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n596), .B1(new_n609), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n606), .A2(new_n608), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n612), .A2(new_n607), .A3(new_n613), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(KEYINPUT99), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n269), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n621));
  INV_X1    g420(.A(new_n619), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n622), .A2(new_n242), .B1(KEYINPUT41), .B2(new_n591), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n620), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n621), .B1(new_n620), .B2(new_n623), .ZN(new_n626));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n627), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n620), .A2(new_n623), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT100), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n629), .B1(new_n631), .B2(new_n624), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n595), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n627), .B1(new_n625), .B2(new_n626), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n631), .A2(new_n624), .A3(new_n629), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n635), .A3(new_n594), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G71gat), .B(G78gat), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n640));
  AND2_X1   g439(.A1(G57gat), .A2(G64gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(G57gat), .A2(G64gat), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT96), .B1(G71gat), .B2(G78gat), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n639), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G71gat), .A2(G78gat), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT9), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OR2_X1    g448(.A1(G57gat), .A2(G64gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(G57gat), .A2(G64gat), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(new_n638), .A3(new_n644), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(KEYINPUT21), .ZN(new_n655));
  XNOR2_X1  g454(.A(G127gat), .B(G155gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n255), .B1(KEYINPUT21), .B2(new_n654), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n657), .B(new_n658), .Z(new_n659));
  NAND2_X1  g458(.A1(G231gat), .A2(G233gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT97), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(G183gat), .B(G211gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT98), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n663), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n659), .B(new_n666), .Z(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT101), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n637), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n633), .A2(new_n636), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT101), .B1(new_n671), .B2(new_n667), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT10), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n674), .B1(new_n646), .B2(new_n653), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(new_n615), .A3(new_n618), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n675), .A2(new_n615), .A3(KEYINPUT103), .A4(new_n618), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(new_n609), .B2(new_n614), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n652), .A2(new_n638), .A3(new_n644), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n638), .B1(new_n652), .B2(new_n644), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n616), .A2(KEYINPUT102), .A3(new_n617), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n682), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n616), .A2(new_n617), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n654), .A2(new_n681), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n674), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n680), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(G230gat), .A2(G233gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT104), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n687), .A2(new_n694), .A3(new_n689), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(G120gat), .B(G148gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(G176gat), .B(G204gat), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n699), .B(new_n700), .Z(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n696), .A2(new_n697), .A3(new_n701), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n673), .A2(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n590), .A2(new_n587), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT105), .B(G1gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1324gat));
  NOR2_X1   g509(.A1(new_n590), .A2(new_n707), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n243), .B1(new_n711), .B2(new_n463), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT16), .B(G8gat), .ZN(new_n713));
  NOR4_X1   g512(.A1(new_n590), .A2(new_n567), .A3(new_n707), .A4(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT42), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(KEYINPUT42), .B2(new_n714), .ZN(G1325gat));
  INV_X1    g515(.A(G15gat), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n711), .A2(new_n717), .A3(new_n552), .A4(new_n558), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT36), .B1(new_n580), .B2(new_n581), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n559), .A2(KEYINPUT36), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n720), .B1(new_n719), .B2(new_n721), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n590), .A2(new_n707), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n718), .B1(new_n717), .B2(new_n725), .ZN(G1326gat));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n380), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT43), .B(G22gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1327gat));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n573), .A2(new_n719), .A3(new_n721), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n585), .A2(new_n561), .A3(new_n564), .A4(new_n558), .ZN(new_n732));
  OAI21_X1  g531(.A(KEYINPUT35), .B1(new_n732), .B2(new_n572), .ZN(new_n733));
  OR3_X1    g532(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n731), .A2(new_n530), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n730), .B1(new_n735), .B2(new_n637), .ZN(new_n736));
  INV_X1    g535(.A(new_n587), .ZN(new_n737));
  OAI211_X1 g536(.A(KEYINPUT44), .B(new_n671), .C1(new_n574), .C2(new_n589), .ZN(new_n738));
  INV_X1    g537(.A(new_n295), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n739), .A2(new_n668), .A3(new_n705), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n736), .A2(new_n737), .A3(new_n738), .A4(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n213), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n742), .B2(new_n741), .ZN(new_n744));
  INV_X1    g543(.A(new_n590), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n668), .A2(new_n705), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n671), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n745), .A2(new_n213), .A3(new_n737), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT45), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n744), .A2(new_n750), .ZN(G1328gat));
  NAND4_X1  g550(.A1(new_n736), .A2(new_n463), .A3(new_n738), .A4(new_n740), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n214), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n753), .B2(new_n752), .ZN(new_n755));
  NOR4_X1   g554(.A1(new_n590), .A2(G36gat), .A3(new_n567), .A4(new_n747), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT46), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(G1329gat));
  NOR2_X1   g557(.A1(new_n590), .A2(new_n747), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n559), .A2(G43gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n719), .A2(new_n721), .ZN(new_n762));
  AND4_X1   g561(.A1(new_n762), .A2(new_n736), .A3(new_n738), .A4(new_n740), .ZN(new_n763));
  OAI211_X1 g562(.A(KEYINPUT47), .B(new_n761), .C1(new_n763), .C2(new_n225), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(KEYINPUT106), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n719), .A2(new_n721), .A3(new_n720), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n736), .A2(new_n767), .A3(new_n738), .A4(new_n740), .ZN(new_n768));
  AOI22_X1  g567(.A1(new_n768), .A2(G43gat), .B1(new_n759), .B2(new_n760), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n764), .B1(new_n769), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g569(.A1(new_n745), .A2(new_n380), .A3(new_n748), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n262), .A2(new_n263), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n585), .A2(new_n772), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n736), .A2(new_n738), .A3(new_n740), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT48), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT48), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n773), .A2(new_n778), .A3(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1331gat));
  NAND3_X1  g579(.A1(new_n673), .A2(new_n739), .A3(new_n705), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n735), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n737), .ZN(new_n783));
  XOR2_X1   g582(.A(KEYINPUT109), .B(G57gat), .Z(new_n784));
  XNOR2_X1  g583(.A(new_n783), .B(new_n784), .ZN(G1332gat));
  NOR3_X1   g584(.A1(new_n735), .A2(new_n567), .A3(new_n781), .ZN(new_n786));
  NOR2_X1   g585(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n787));
  AND2_X1   g586(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n786), .B2(new_n787), .ZN(G1333gat));
  NAND2_X1  g589(.A1(new_n782), .A2(new_n767), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n559), .A2(G71gat), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n791), .A2(G71gat), .B1(new_n782), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g593(.A1(new_n782), .A2(new_n380), .ZN(new_n795));
  XNOR2_X1  g594(.A(KEYINPUT110), .B(G78gat), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n795), .B(new_n796), .ZN(G1335gat));
  NOR3_X1   g596(.A1(new_n668), .A2(new_n295), .A3(new_n706), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n736), .A2(new_n737), .A3(new_n738), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(G85gat), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n587), .A2(G85gat), .A3(new_n706), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n530), .A2(new_n566), .A3(new_n573), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n733), .A2(new_n734), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n637), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n668), .A2(new_n295), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n804), .A2(KEYINPUT51), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT51), .B1(new_n804), .B2(new_n805), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n801), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n800), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n800), .A2(new_n808), .A3(KEYINPUT111), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(G1336gat));
  NAND4_X1  g612(.A1(new_n736), .A2(new_n463), .A3(new_n738), .A4(new_n798), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G92gat), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n567), .A2(G92gat), .A3(new_n706), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n806), .B2(new_n807), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT52), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n815), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(G1337gat));
  XOR2_X1   g621(.A(KEYINPUT112), .B(G99gat), .Z(new_n823));
  NAND3_X1  g622(.A1(new_n736), .A2(new_n738), .A3(new_n798), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(new_n724), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n559), .A2(new_n706), .A3(new_n823), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n826), .B1(new_n806), .B2(new_n807), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(G1338gat));
  NAND4_X1  g627(.A1(new_n736), .A2(new_n380), .A3(new_n738), .A4(new_n798), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(G106gat), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n585), .A2(G106gat), .A3(new_n706), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n806), .B2(new_n807), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT53), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n830), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(G1339gat));
  AOI21_X1  g636(.A(new_n694), .B1(new_n680), .B2(new_n691), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n680), .A2(new_n691), .A3(new_n694), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n843));
  AOI211_X1 g642(.A(new_n843), .B(new_n701), .C1(new_n838), .C2(new_n839), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n692), .A2(new_n839), .A3(new_n695), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT113), .B1(new_n845), .B2(new_n702), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n842), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n704), .ZN(new_n850));
  AOI211_X1 g649(.A(KEYINPUT54), .B(new_n694), .C1(new_n680), .C2(new_n691), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n843), .B1(new_n851), .B2(new_n701), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n845), .A2(KEYINPUT113), .A3(new_n702), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n848), .B1(new_n840), .B2(new_n841), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n850), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n295), .A2(new_n849), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n257), .B1(new_n284), .B2(new_n256), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n275), .A2(new_n276), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n205), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n705), .B(new_n860), .C1(new_n293), .C2(new_n294), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n671), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n855), .B1(new_n844), .B2(new_n846), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n852), .A2(new_n853), .B1(new_n841), .B2(new_n840), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n863), .B(new_n704), .C1(new_n864), .C2(KEYINPUT55), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n298), .A2(new_n860), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n865), .A2(new_n637), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n667), .B1(new_n862), .B2(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n670), .A2(new_n739), .A3(new_n672), .A4(new_n706), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n576), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n587), .A2(new_n463), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n301), .ZN(new_n877));
  OAI21_X1  g676(.A(G113gat), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n587), .B1(new_n868), .B2(new_n869), .ZN(new_n879));
  INV_X1    g678(.A(new_n732), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(new_n463), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n739), .A2(G113gat), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT114), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n878), .A2(new_n885), .ZN(G1340gat));
  AOI21_X1  g685(.A(G120gat), .B1(new_n882), .B2(new_n705), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n705), .A2(G120gat), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n875), .B2(new_n888), .ZN(G1341gat));
  OAI21_X1  g688(.A(G127gat), .B1(new_n876), .B2(new_n667), .ZN(new_n890));
  INV_X1    g689(.A(G127gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n882), .A2(new_n891), .A3(new_n668), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1342gat));
  OR4_X1    g692(.A1(G134gat), .A2(new_n881), .A3(new_n463), .A4(new_n637), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n894), .A2(KEYINPUT56), .ZN(new_n895));
  OAI21_X1  g694(.A(G134gat), .B1(new_n876), .B2(new_n637), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(KEYINPUT56), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G1343gat));
  INV_X1    g697(.A(KEYINPUT116), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n861), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n298), .A2(KEYINPUT116), .A3(new_n705), .A4(new_n860), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n847), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n856), .A3(KEYINPUT118), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n298), .A2(new_n299), .A3(new_n286), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n299), .B1(new_n298), .B2(new_n286), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT118), .B1(new_n904), .B2(new_n856), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n902), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n867), .B1(new_n910), .B2(new_n637), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n869), .B1(new_n911), .B2(new_n668), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n380), .A2(KEYINPUT57), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g714(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n917), .B1(new_n870), .B2(new_n380), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n874), .A2(new_n762), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n920), .A2(KEYINPUT122), .A3(new_n301), .A4(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n903), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n863), .B(new_n704), .C1(new_n864), .C2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT118), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n301), .A2(new_n926), .A3(new_n905), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n671), .B1(new_n927), .B2(new_n902), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n667), .B1(new_n928), .B2(new_n867), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n913), .B1(new_n929), .B2(new_n869), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n301), .B(new_n921), .C1(new_n930), .C2(new_n918), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n922), .A2(new_n933), .A3(G141gat), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n765), .A2(new_n380), .A3(new_n766), .ZN(new_n936));
  INV_X1    g735(.A(new_n879), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n724), .A2(KEYINPUT121), .A3(new_n380), .A4(new_n879), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n938), .A2(new_n567), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n301), .A2(new_n322), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT120), .Z(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT58), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n934), .A2(new_n944), .ZN(new_n945));
  NOR4_X1   g744(.A1(new_n936), .A2(new_n937), .A3(new_n942), .A4(new_n463), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n918), .B1(new_n912), .B2(new_n914), .ZN(new_n947));
  INV_X1    g746(.A(new_n921), .ZN(new_n948));
  OAI21_X1  g747(.A(KEYINPUT119), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT119), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n950), .B(new_n921), .C1(new_n930), .C2(new_n918), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n949), .A2(new_n295), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n946), .B1(new_n952), .B2(G141gat), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT58), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n945), .B1(new_n953), .B2(new_n954), .ZN(G1344gat));
  NAND3_X1  g754(.A1(new_n949), .A2(new_n705), .A3(new_n951), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G148gat), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT59), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(KEYINPUT123), .B1(new_n865), .B2(new_n637), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n671), .A2(new_n849), .A3(new_n856), .A4(new_n961), .ZN(new_n962));
  AND4_X1   g761(.A1(new_n298), .A2(new_n960), .A3(new_n860), .A4(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n667), .B1(new_n928), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n964), .B1(new_n301), .B2(new_n707), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT57), .B1(new_n965), .B2(new_n380), .ZN(new_n966));
  AOI211_X1 g765(.A(new_n585), .B(new_n916), .C1(new_n868), .C2(new_n869), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n705), .B(new_n921), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n958), .A2(new_n324), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n706), .A2(G148gat), .ZN(new_n970));
  AOI22_X1  g769(.A1(new_n968), .A2(new_n969), .B1(new_n940), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n959), .A2(new_n971), .ZN(G1345gat));
  NAND2_X1  g771(.A1(new_n949), .A2(new_n951), .ZN(new_n973));
  OAI21_X1  g772(.A(G155gat), .B1(new_n973), .B2(new_n667), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n940), .A2(new_n328), .A3(new_n668), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1346gat));
  OAI21_X1  g775(.A(G162gat), .B1(new_n973), .B2(new_n637), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n463), .A2(G162gat), .A3(new_n637), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n938), .A2(new_n939), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1347gat));
  NOR2_X1   g779(.A1(new_n737), .A2(new_n567), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n870), .A2(new_n871), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(G169gat), .B1(new_n982), .B2(new_n877), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT125), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n870), .A2(new_n587), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT124), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n567), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n870), .A2(KEYINPUT124), .A3(new_n587), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(new_n880), .ZN(new_n990));
  INV_X1    g789(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n295), .A2(new_n419), .ZN(new_n992));
  INV_X1    g791(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n984), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  NOR3_X1   g793(.A1(new_n990), .A2(KEYINPUT125), .A3(new_n992), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n983), .B1(new_n994), .B2(new_n995), .ZN(G1348gat));
  OAI21_X1  g795(.A(G176gat), .B1(new_n982), .B2(new_n706), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n705), .A2(new_n399), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n997), .B1(new_n990), .B2(new_n998), .ZN(G1349gat));
  OAI21_X1  g798(.A(G183gat), .B1(new_n982), .B2(new_n667), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n668), .A2(new_n386), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n1000), .B1(new_n990), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1002), .A2(KEYINPUT60), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT60), .ZN(new_n1004));
  OAI211_X1 g803(.A(new_n1004), .B(new_n1000), .C1(new_n990), .C2(new_n1001), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1003), .A2(new_n1005), .ZN(G1350gat));
  OAI21_X1  g805(.A(G190gat), .B1(new_n982), .B2(new_n637), .ZN(new_n1007));
  XNOR2_X1  g806(.A(new_n1007), .B(KEYINPUT61), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n671), .A2(new_n381), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n1008), .B1(new_n990), .B2(new_n1009), .ZN(G1351gat));
  INV_X1    g809(.A(new_n936), .ZN(new_n1011));
  AND2_X1   g810(.A1(new_n989), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g811(.A(G197gat), .B1(new_n1012), .B2(new_n295), .ZN(new_n1013));
  OR2_X1    g812(.A1(new_n966), .A2(new_n967), .ZN(new_n1014));
  AND2_X1   g813(.A1(new_n724), .A2(new_n981), .ZN(new_n1015));
  AND2_X1   g814(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AND2_X1   g815(.A1(new_n301), .A2(G197gat), .ZN(new_n1017));
  AOI21_X1  g816(.A(new_n1013), .B1(new_n1016), .B2(new_n1017), .ZN(G1352gat));
  NAND2_X1  g817(.A1(new_n989), .A2(new_n1011), .ZN(new_n1019));
  OR2_X1    g818(.A1(new_n706), .A2(G204gat), .ZN(new_n1020));
  OR3_X1    g819(.A1(new_n1019), .A2(KEYINPUT62), .A3(new_n1020), .ZN(new_n1021));
  OAI211_X1 g820(.A(new_n705), .B(new_n1015), .C1(new_n966), .C2(new_n967), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1022), .A2(G204gat), .ZN(new_n1023));
  OAI21_X1  g822(.A(KEYINPUT62), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1024));
  NAND3_X1  g823(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .ZN(G1353gat));
  OAI211_X1 g824(.A(new_n668), .B(new_n1015), .C1(new_n966), .C2(new_n967), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1026), .A2(G211gat), .ZN(new_n1027));
  NAND2_X1  g826(.A1(new_n1027), .A2(KEYINPUT63), .ZN(new_n1028));
  NOR2_X1   g827(.A1(new_n667), .A2(G211gat), .ZN(new_n1029));
  NAND3_X1  g828(.A1(new_n989), .A2(new_n1011), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g829(.A1(new_n1030), .A2(KEYINPUT126), .ZN(new_n1031));
  INV_X1    g830(.A(KEYINPUT126), .ZN(new_n1032));
  NAND4_X1  g831(.A1(new_n989), .A2(new_n1032), .A3(new_n1011), .A4(new_n1029), .ZN(new_n1033));
  NAND2_X1  g832(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g833(.A(KEYINPUT63), .ZN(new_n1035));
  NAND3_X1  g834(.A1(new_n1026), .A2(new_n1035), .A3(G211gat), .ZN(new_n1036));
  NAND3_X1  g835(.A1(new_n1028), .A2(new_n1034), .A3(new_n1036), .ZN(G1354gat));
  NOR2_X1   g836(.A1(new_n637), .A2(new_n305), .ZN(new_n1038));
  OAI211_X1 g837(.A(new_n1015), .B(new_n1038), .C1(new_n966), .C2(new_n967), .ZN(new_n1039));
  NAND4_X1  g838(.A1(new_n987), .A2(new_n1011), .A3(new_n671), .A4(new_n988), .ZN(new_n1040));
  NAND2_X1  g839(.A1(new_n1040), .A2(new_n313), .ZN(new_n1041));
  NAND2_X1  g840(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g841(.A1(new_n1042), .A2(KEYINPUT127), .ZN(new_n1043));
  INV_X1    g842(.A(KEYINPUT127), .ZN(new_n1044));
  NAND3_X1  g843(.A1(new_n1039), .A2(new_n1044), .A3(new_n1041), .ZN(new_n1045));
  NAND2_X1  g844(.A1(new_n1043), .A2(new_n1045), .ZN(G1355gat));
endmodule


