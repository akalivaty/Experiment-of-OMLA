

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783;

  NAND2_X1 U365 ( .A1(n360), .A2(n359), .ZN(n417) );
  NOR2_X1 U366 ( .A1(n592), .A2(n591), .ZN(n593) );
  OR2_X1 U367 ( .A1(n646), .A2(G902), .ZN(n355) );
  XNOR2_X1 U368 ( .A(n517), .B(n402), .ZN(n699) );
  BUF_X1 U369 ( .A(G143), .Z(n344) );
  XNOR2_X1 U370 ( .A(n490), .B(n521), .ZN(n668) );
  INV_X1 U371 ( .A(G953), .ZN(n769) );
  NOR2_X2 U372 ( .A1(n622), .A2(n579), .ZN(n581) );
  NAND2_X2 U373 ( .A1(n385), .A2(n608), .ZN(n354) );
  AND2_X2 U374 ( .A1(n662), .A2(n645), .ZN(n475) );
  BUF_X1 U375 ( .A(G113), .Z(n379) );
  OR2_X1 U376 ( .A1(n426), .A2(KEYINPUT110), .ZN(n345) );
  XNOR2_X2 U377 ( .A(n520), .B(n519), .ZN(n735) );
  NOR2_X2 U378 ( .A1(n782), .A2(n637), .ZN(n373) );
  NAND2_X1 U379 ( .A1(n512), .A2(n765), .ZN(n460) );
  NOR2_X1 U380 ( .A1(G953), .A2(G237), .ZN(n524) );
  NAND2_X1 U381 ( .A1(n398), .A2(n396), .ZN(n783) );
  XNOR2_X1 U382 ( .A(n505), .B(n504), .ZN(n709) );
  INV_X1 U383 ( .A(KEYINPUT3), .ZN(n469) );
  AND2_X1 U384 ( .A1(n424), .A2(n422), .ZN(n450) );
  AND2_X1 U385 ( .A1(n425), .A2(n345), .ZN(n424) );
  NAND2_X1 U386 ( .A1(n367), .A2(n441), .ZN(n378) );
  NOR2_X1 U387 ( .A1(n442), .A2(n443), .ZN(n367) );
  NAND2_X1 U388 ( .A1(n431), .A2(n428), .ZN(n427) );
  OR2_X1 U389 ( .A1(n568), .A2(n432), .ZN(n431) );
  XNOR2_X1 U390 ( .A(n421), .B(n565), .ZN(n611) );
  NAND2_X1 U391 ( .A1(n364), .A2(n564), .ZN(n421) );
  XNOR2_X1 U392 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U393 ( .A(n470), .B(n469), .ZN(n472) );
  NAND2_X1 U394 ( .A1(n414), .A2(n413), .ZN(n628) );
  XNOR2_X2 U395 ( .A(n366), .B(n644), .ZN(n772) );
  XNOR2_X2 U396 ( .A(n573), .B(n452), .ZN(n575) );
  NOR2_X1 U397 ( .A1(n563), .A2(n571), .ZN(n363) );
  XNOR2_X2 U398 ( .A(n515), .B(n406), .ZN(n766) );
  XNOR2_X1 U399 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n669) );
  AND2_X1 U400 ( .A1(n419), .A2(n762), .ZN(n418) );
  NAND2_X1 U401 ( .A1(n764), .A2(n615), .ZN(n419) );
  INV_X1 U402 ( .A(n569), .ZN(n430) );
  XNOR2_X1 U403 ( .A(n611), .B(KEYINPUT109), .ZN(n568) );
  XNOR2_X1 U404 ( .A(n669), .B(G101), .ZN(n512) );
  AND2_X1 U405 ( .A1(n356), .A2(n418), .ZN(n361) );
  INV_X1 U406 ( .A(n373), .ZN(n371) );
  INV_X1 U407 ( .A(KEYINPUT44), .ZN(n370) );
  AND2_X1 U408 ( .A1(n706), .A2(n705), .ZN(n619) );
  AND2_X1 U409 ( .A1(n429), .A2(n706), .ZN(n428) );
  NAND2_X1 U410 ( .A1(n567), .A2(n430), .ZN(n429) );
  NOR2_X1 U411 ( .A1(n571), .A2(n713), .ZN(n383) );
  NAND2_X1 U412 ( .A1(n368), .A2(n705), .ZN(n622) );
  AND2_X1 U413 ( .A1(n559), .A2(n482), .ZN(n483) );
  XNOR2_X1 U414 ( .A(n503), .B(n502), .ZN(n504) );
  INV_X1 U415 ( .A(KEYINPUT25), .ZN(n502) );
  XNOR2_X1 U416 ( .A(KEYINPUT5), .B(G137), .ZN(n510) );
  XNOR2_X1 U417 ( .A(KEYINPUT98), .B(KEYINPUT23), .ZN(n492) );
  NAND2_X1 U418 ( .A1(n411), .A2(G475), .ZN(n408) );
  XNOR2_X1 U419 ( .A(n527), .B(n526), .ZN(n534) );
  NAND2_X1 U420 ( .A1(n459), .A2(n460), .ZN(n485) );
  XOR2_X1 U421 ( .A(G137), .B(G140), .Z(n490) );
  NAND2_X1 U422 ( .A1(n757), .A2(n401), .ZN(n399) );
  XNOR2_X1 U423 ( .A(n377), .B(KEYINPUT39), .ZN(n616) );
  NOR2_X1 U424 ( .A1(n592), .A2(n584), .ZN(n377) );
  BUF_X1 U425 ( .A(n709), .Z(n376) );
  XOR2_X1 U426 ( .A(KEYINPUT68), .B(KEYINPUT48), .Z(n608) );
  INV_X1 U427 ( .A(KEYINPUT67), .ZN(n488) );
  INV_X1 U428 ( .A(n725), .ZN(n451) );
  XNOR2_X1 U429 ( .A(n553), .B(KEYINPUT6), .ZN(n563) );
  XNOR2_X1 U430 ( .A(G110), .B(KEYINPUT97), .ZN(n494) );
  INV_X1 U431 ( .A(G128), .ZN(n464) );
  XNOR2_X1 U432 ( .A(n379), .B(n344), .ZN(n528) );
  XNOR2_X1 U433 ( .A(n525), .B(n455), .ZN(n526) );
  INV_X1 U434 ( .A(KEYINPUT106), .ZN(n452) );
  INV_X1 U435 ( .A(KEYINPUT103), .ZN(n362) );
  XNOR2_X1 U436 ( .A(n614), .B(KEYINPUT38), .ZN(n721) );
  XNOR2_X1 U437 ( .A(n508), .B(n507), .ZN(n708) );
  BUF_X1 U438 ( .A(n563), .Z(n630) );
  XNOR2_X1 U439 ( .A(n448), .B(G107), .ZN(n765) );
  XNOR2_X1 U440 ( .A(G104), .B(G110), .ZN(n448) );
  XNOR2_X1 U441 ( .A(n473), .B(G122), .ZN(n406) );
  XOR2_X1 U442 ( .A(G107), .B(KEYINPUT7), .Z(n540) );
  XNOR2_X1 U443 ( .A(n405), .B(n404), .ZN(n662) );
  XNOR2_X1 U444 ( .A(n485), .B(n407), .ZN(n404) );
  XNOR2_X1 U445 ( .A(n766), .B(n468), .ZN(n405) );
  XNOR2_X1 U446 ( .A(n463), .B(KEYINPUT72), .ZN(n407) );
  NAND2_X1 U447 ( .A1(n418), .A2(n350), .ZN(n359) );
  INV_X1 U448 ( .A(n590), .ZN(n444) );
  AND2_X1 U449 ( .A1(n624), .A2(KEYINPUT34), .ZN(n443) );
  NAND2_X1 U450 ( .A1(n446), .A2(n447), .ZN(n441) );
  NOR2_X1 U451 ( .A1(n735), .A2(KEYINPUT34), .ZN(n447) );
  XNOR2_X1 U452 ( .A(n620), .B(n621), .ZN(n625) );
  XNOR2_X1 U453 ( .A(n358), .B(n357), .ZN(n582) );
  INV_X1 U454 ( .A(KEYINPUT30), .ZN(n357) );
  OR2_X1 U455 ( .A1(n572), .A2(n353), .ZN(n597) );
  INV_X1 U456 ( .A(KEYINPUT28), .ZN(n382) );
  XNOR2_X1 U457 ( .A(n535), .B(KEYINPUT13), .ZN(n536) );
  INV_X1 U458 ( .A(G475), .ZN(n535) );
  XNOR2_X1 U459 ( .A(n517), .B(n516), .ZN(n646) );
  NAND2_X1 U460 ( .A1(n411), .A2(G472), .ZN(n409) );
  XNOR2_X1 U461 ( .A(G119), .B(G128), .ZN(n498) );
  OR2_X2 U462 ( .A1(n704), .A2(n645), .ZN(n412) );
  XNOR2_X1 U463 ( .A(n653), .B(n652), .ZN(n654) );
  INV_X1 U464 ( .A(n412), .ZN(n696) );
  XNOR2_X1 U465 ( .A(n485), .B(n403), .ZN(n402) );
  XNOR2_X1 U466 ( .A(n486), .B(KEYINPUT72), .ZN(n403) );
  NAND2_X1 U467 ( .A1(n411), .A2(G210), .ZN(n410) );
  NAND2_X1 U468 ( .A1(n393), .A2(n390), .ZN(n780) );
  NAND2_X1 U469 ( .A1(n392), .A2(n391), .ZN(n390) );
  AND2_X1 U470 ( .A1(n395), .A2(n394), .ZN(n393) );
  NOR2_X1 U471 ( .A1(n597), .A2(n578), .ZN(n391) );
  OR2_X1 U472 ( .A1(n616), .A2(n397), .ZN(n396) );
  AND2_X1 U473 ( .A1(n400), .A2(n399), .ZN(n398) );
  NAND2_X1 U474 ( .A1(n564), .A2(KEYINPUT40), .ZN(n397) );
  NAND2_X1 U475 ( .A1(n423), .A2(n346), .ZN(n422) );
  INV_X1 U476 ( .A(n625), .ZN(n760) );
  INV_X1 U477 ( .A(n376), .ZN(n413) );
  INV_X1 U478 ( .A(KEYINPUT87), .ZN(n415) );
  INV_X1 U479 ( .A(n757), .ZN(n564) );
  AND2_X1 U480 ( .A1(n426), .A2(KEYINPUT110), .ZN(n346) );
  AND2_X1 U481 ( .A1(n380), .A2(n627), .ZN(n347) );
  XOR2_X1 U482 ( .A(n497), .B(n496), .Z(n348) );
  NOR2_X1 U483 ( .A1(n727), .A2(n735), .ZN(n349) );
  NAND2_X1 U484 ( .A1(n449), .A2(KEYINPUT85), .ZN(n350) );
  AND2_X1 U485 ( .A1(n575), .A2(n451), .ZN(n351) );
  INV_X1 U486 ( .A(KEYINPUT40), .ZN(n401) );
  INV_X1 U487 ( .A(KEYINPUT110), .ZN(n434) );
  XNOR2_X1 U488 ( .A(KEYINPUT15), .B(G902), .ZN(n645) );
  NAND2_X1 U489 ( .A1(n352), .A2(n594), .ZN(n375) );
  XNOR2_X1 U490 ( .A(n352), .B(n781), .ZN(G45) );
  XNOR2_X1 U491 ( .A(n593), .B(KEYINPUT105), .ZN(n352) );
  XNOR2_X1 U492 ( .A(n368), .B(KEYINPUT1), .ZN(n706) );
  INV_X1 U493 ( .A(n368), .ZN(n353) );
  XNOR2_X2 U494 ( .A(n440), .B(G469), .ZN(n368) );
  NAND2_X1 U495 ( .A1(n354), .A2(n356), .ZN(n420) );
  NAND2_X1 U496 ( .A1(n361), .A2(n354), .ZN(n360) );
  XNOR2_X2 U497 ( .A(n355), .B(G472), .ZN(n553) );
  NAND2_X1 U498 ( .A1(n387), .A2(n450), .ZN(n356) );
  NAND2_X1 U499 ( .A1(n553), .A2(n720), .ZN(n358) );
  NAND2_X1 U500 ( .A1(n365), .A2(n372), .ZN(n643) );
  NAND2_X1 U501 ( .A1(n371), .A2(n369), .ZN(n365) );
  NAND2_X1 U502 ( .A1(n439), .A2(n643), .ZN(n366) );
  AND2_X1 U503 ( .A1(n639), .A2(n370), .ZN(n369) );
  NAND2_X1 U504 ( .A1(n373), .A2(n642), .ZN(n372) );
  NAND2_X1 U505 ( .A1(n438), .A2(n374), .ZN(n439) );
  NAND2_X1 U506 ( .A1(n436), .A2(n347), .ZN(n374) );
  INV_X1 U507 ( .A(n450), .ZN(n607) );
  NAND2_X1 U508 ( .A1(n386), .A2(n450), .ZN(n385) );
  NOR2_X2 U509 ( .A1(n772), .A2(n674), .ZN(n384) );
  NAND2_X2 U510 ( .A1(n417), .A2(n416), .ZN(n674) );
  XNOR2_X1 U511 ( .A(n375), .B(KEYINPUT83), .ZN(n603) );
  OR2_X2 U512 ( .A1(n420), .A2(KEYINPUT85), .ZN(n416) );
  NOR2_X2 U513 ( .A1(n783), .A2(n780), .ZN(n586) );
  XNOR2_X2 U514 ( .A(n378), .B(n549), .ZN(n638) );
  INV_X1 U515 ( .A(n427), .ZN(n423) );
  XNOR2_X1 U516 ( .A(n636), .B(KEYINPUT32), .ZN(n782) );
  OR2_X1 U517 ( .A1(n626), .A2(n725), .ZN(n380) );
  NAND2_X1 U518 ( .A1(n381), .A2(n603), .ZN(n604) );
  NAND2_X1 U519 ( .A1(n602), .A2(n601), .ZN(n381) );
  XNOR2_X1 U520 ( .A(n383), .B(n382), .ZN(n572) );
  NOR2_X2 U521 ( .A1(n597), .A2(n596), .ZN(n755) );
  INV_X1 U522 ( .A(n512), .ZN(n458) );
  XNOR2_X2 U523 ( .A(n384), .B(KEYINPUT2), .ZN(n704) );
  AND2_X1 U524 ( .A1(n606), .A2(n605), .ZN(n386) );
  AND2_X1 U525 ( .A1(n606), .A2(n388), .ZN(n387) );
  AND2_X1 U526 ( .A1(n605), .A2(n389), .ZN(n388) );
  INV_X1 U527 ( .A(n608), .ZN(n389) );
  INV_X1 U528 ( .A(n736), .ZN(n392) );
  NAND2_X1 U529 ( .A1(n597), .A2(n578), .ZN(n394) );
  NAND2_X1 U530 ( .A1(n736), .A2(n578), .ZN(n395) );
  NAND2_X1 U531 ( .A1(n616), .A2(n401), .ZN(n400) );
  XNOR2_X2 U532 ( .A(n577), .B(n576), .ZN(n736) );
  XNOR2_X2 U533 ( .A(n472), .B(n471), .ZN(n515) );
  OR2_X1 U534 ( .A1(n704), .A2(n408), .ZN(n655) );
  OR2_X1 U535 ( .A1(n704), .A2(n409), .ZN(n648) );
  OR2_X1 U536 ( .A1(n704), .A2(n410), .ZN(n664) );
  INV_X1 U537 ( .A(n645), .ZN(n411) );
  NOR2_X1 U538 ( .A1(n412), .A2(n547), .ZN(n693) );
  INV_X1 U539 ( .A(n628), .ZN(n743) );
  NAND2_X1 U540 ( .A1(n628), .A2(KEYINPUT88), .ZN(n437) );
  XNOR2_X1 U541 ( .A(n618), .B(n415), .ZN(n414) );
  XNOR2_X1 U542 ( .A(n500), .B(n499), .ZN(n688) );
  XOR2_X2 U543 ( .A(G146), .B(G125), .Z(n489) );
  XNOR2_X2 U544 ( .A(KEYINPUT10), .B(n489), .ZN(n521) );
  XNOR2_X1 U545 ( .A(n552), .B(n551), .ZN(n635) );
  INV_X1 U546 ( .A(n437), .ZN(n436) );
  NAND2_X1 U547 ( .A1(n427), .A2(n434), .ZN(n425) );
  NAND2_X1 U548 ( .A1(n568), .A2(n430), .ZN(n426) );
  NAND2_X1 U549 ( .A1(n433), .A2(n569), .ZN(n432) );
  INV_X1 U550 ( .A(n567), .ZN(n433) );
  NAND2_X1 U551 ( .A1(n435), .A2(n629), .ZN(n438) );
  NAND2_X1 U552 ( .A1(n347), .A2(n628), .ZN(n435) );
  NAND2_X1 U553 ( .A1(n699), .A2(n546), .ZN(n440) );
  NAND2_X1 U554 ( .A1(n445), .A2(n444), .ZN(n442) );
  NAND2_X1 U555 ( .A1(n735), .A2(KEYINPUT34), .ZN(n445) );
  INV_X1 U556 ( .A(n624), .ZN(n446) );
  XNOR2_X2 U557 ( .A(n484), .B(KEYINPUT0), .ZN(n624) );
  INV_X1 U558 ( .A(n764), .ZN(n449) );
  XNOR2_X2 U559 ( .A(n672), .B(G146), .ZN(n517) );
  NOR2_X2 U560 ( .A1(n709), .A2(n708), .ZN(n705) );
  AND2_X1 U561 ( .A1(n538), .A2(G221), .ZN(n453) );
  AND2_X1 U562 ( .A1(G227), .A2(n769), .ZN(n454) );
  AND2_X1 U563 ( .A1(G214), .A2(n524), .ZN(n455) );
  NAND2_X1 U564 ( .A1(n557), .A2(n556), .ZN(n757) );
  OR2_X1 U565 ( .A1(n724), .A2(n708), .ZN(n456) );
  INV_X1 U566 ( .A(KEYINPUT85), .ZN(n615) );
  INV_X1 U567 ( .A(KEYINPUT88), .ZN(n629) );
  XNOR2_X1 U568 ( .A(n490), .B(n454), .ZN(n486) );
  INV_X1 U569 ( .A(n721), .ZN(n584) );
  INV_X1 U570 ( .A(KEYINPUT77), .ZN(n580) );
  XNOR2_X1 U571 ( .A(n668), .B(n453), .ZN(n500) );
  XNOR2_X1 U572 ( .A(n537), .B(n536), .ZN(n588) );
  INV_X1 U573 ( .A(n765), .ZN(n457) );
  NAND2_X1 U574 ( .A1(n458), .A2(n457), .ZN(n459) );
  XOR2_X1 U575 ( .A(KEYINPUT18), .B(KEYINPUT95), .Z(n462) );
  XNOR2_X1 U576 ( .A(KEYINPUT79), .B(KEYINPUT17), .ZN(n461) );
  XNOR2_X1 U577 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X2 U578 ( .A(KEYINPUT82), .B(G143), .ZN(n465) );
  XNOR2_X2 U579 ( .A(n465), .B(n464), .ZN(n487) );
  NAND2_X1 U580 ( .A1(G224), .A2(n769), .ZN(n466) );
  XNOR2_X1 U581 ( .A(n466), .B(n489), .ZN(n467) );
  XNOR2_X1 U582 ( .A(n487), .B(n467), .ZN(n468) );
  XOR2_X1 U583 ( .A(KEYINPUT74), .B(KEYINPUT16), .Z(n473) );
  XNOR2_X2 U584 ( .A(G116), .B(G113), .ZN(n470) );
  XOR2_X1 U585 ( .A(KEYINPUT70), .B(G119), .Z(n471) );
  OR2_X1 U586 ( .A1(G237), .A2(G902), .ZN(n476) );
  AND2_X1 U587 ( .A1(n476), .A2(G210), .ZN(n474) );
  XNOR2_X2 U588 ( .A(n475), .B(n474), .ZN(n614) );
  NAND2_X1 U589 ( .A1(G214), .A2(n476), .ZN(n720) );
  INV_X1 U590 ( .A(n720), .ZN(n609) );
  NOR2_X1 U591 ( .A1(n614), .A2(n609), .ZN(n477) );
  XNOR2_X1 U592 ( .A(n477), .B(KEYINPUT91), .ZN(n566) );
  XNOR2_X1 U593 ( .A(n566), .B(KEYINPUT19), .ZN(n595) );
  NAND2_X1 U594 ( .A1(G234), .A2(G237), .ZN(n478) );
  XNOR2_X1 U595 ( .A(n478), .B(KEYINPUT14), .ZN(n731) );
  INV_X1 U596 ( .A(G902), .ZN(n546) );
  NAND2_X1 U597 ( .A1(G953), .A2(n546), .ZN(n479) );
  NAND2_X1 U598 ( .A1(n731), .A2(n479), .ZN(n481) );
  NOR2_X1 U599 ( .A1(G953), .A2(G952), .ZN(n480) );
  NOR2_X1 U600 ( .A1(n481), .A2(n480), .ZN(n559) );
  NAND2_X1 U601 ( .A1(G953), .A2(G898), .ZN(n482) );
  NAND2_X1 U602 ( .A1(n595), .A2(n483), .ZN(n484) );
  XNOR2_X2 U603 ( .A(n487), .B(G134), .ZN(n543) );
  XNOR2_X1 U604 ( .A(n488), .B(G131), .ZN(n530) );
  XNOR2_X2 U605 ( .A(n543), .B(n530), .ZN(n672) );
  NAND2_X1 U606 ( .A1(n769), .A2(G234), .ZN(n491) );
  XOR2_X1 U607 ( .A(KEYINPUT8), .B(n491), .Z(n538) );
  XOR2_X1 U608 ( .A(KEYINPUT24), .B(KEYINPUT71), .Z(n493) );
  XNOR2_X1 U609 ( .A(n493), .B(n492), .ZN(n497) );
  XOR2_X1 U610 ( .A(KEYINPUT96), .B(KEYINPUT78), .Z(n495) );
  XNOR2_X1 U611 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U612 ( .A(n348), .B(n498), .ZN(n499) );
  NOR2_X1 U613 ( .A1(G902), .A2(n688), .ZN(n505) );
  NAND2_X1 U614 ( .A1(G234), .A2(n645), .ZN(n501) );
  XNOR2_X1 U615 ( .A(KEYINPUT20), .B(n501), .ZN(n506) );
  NAND2_X1 U616 ( .A1(n506), .A2(G217), .ZN(n503) );
  XOR2_X1 U617 ( .A(KEYINPUT99), .B(KEYINPUT21), .Z(n508) );
  NAND2_X1 U618 ( .A1(G221), .A2(n506), .ZN(n507) );
  NAND2_X1 U619 ( .A1(n524), .A2(G210), .ZN(n509) );
  XNOR2_X1 U620 ( .A(n509), .B(KEYINPUT76), .ZN(n511) );
  XNOR2_X1 U621 ( .A(n511), .B(n510), .ZN(n513) );
  XNOR2_X1 U622 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U623 ( .A(n515), .B(n514), .ZN(n516) );
  INV_X1 U624 ( .A(n630), .ZN(n518) );
  NAND2_X1 U625 ( .A1(n619), .A2(n518), .ZN(n520) );
  XNOR2_X1 U626 ( .A(KEYINPUT93), .B(KEYINPUT33), .ZN(n519) );
  INV_X1 U627 ( .A(n521), .ZN(n527) );
  XOR2_X1 U628 ( .A(KEYINPUT12), .B(KEYINPUT101), .Z(n523) );
  XNOR2_X1 U629 ( .A(G140), .B(KEYINPUT11), .ZN(n522) );
  XNOR2_X1 U630 ( .A(n523), .B(n522), .ZN(n525) );
  XOR2_X1 U631 ( .A(G104), .B(G122), .Z(n529) );
  XNOR2_X1 U632 ( .A(n529), .B(n528), .ZN(n532) );
  XOR2_X1 U633 ( .A(KEYINPUT102), .B(n530), .Z(n531) );
  XNOR2_X1 U634 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U635 ( .A(n534), .B(n533), .ZN(n653) );
  NOR2_X1 U636 ( .A1(G902), .A2(n653), .ZN(n537) );
  INV_X1 U637 ( .A(n588), .ZN(n557) );
  NAND2_X1 U638 ( .A1(G217), .A2(n538), .ZN(n539) );
  XNOR2_X1 U639 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U640 ( .A(n541), .B(KEYINPUT9), .Z(n545) );
  XNOR2_X1 U641 ( .A(G116), .B(G122), .ZN(n542) );
  XNOR2_X1 U642 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U643 ( .A(n545), .B(n544), .ZN(n694) );
  NAND2_X1 U644 ( .A1(n694), .A2(n546), .ZN(n548) );
  INV_X1 U645 ( .A(G478), .ZN(n547) );
  XNOR2_X1 U646 ( .A(n548), .B(n547), .ZN(n556) );
  INV_X1 U647 ( .A(n556), .ZN(n587) );
  NAND2_X1 U648 ( .A1(n557), .A2(n587), .ZN(n590) );
  XNOR2_X1 U649 ( .A(KEYINPUT80), .B(KEYINPUT35), .ZN(n549) );
  XNOR2_X1 U650 ( .A(G122), .B(KEYINPUT127), .ZN(n550) );
  XNOR2_X1 U651 ( .A(n638), .B(n550), .ZN(G24) );
  NAND2_X1 U652 ( .A1(n556), .A2(n588), .ZN(n724) );
  NOR2_X1 U653 ( .A1(n624), .A2(n456), .ZN(n552) );
  XNOR2_X1 U654 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n551) );
  INV_X1 U655 ( .A(n553), .ZN(n713) );
  NAND2_X1 U656 ( .A1(n376), .A2(n713), .ZN(n554) );
  OR2_X1 U657 ( .A1(n706), .A2(n554), .ZN(n555) );
  NOR2_X1 U658 ( .A1(n635), .A2(n555), .ZN(n637) );
  XOR2_X1 U659 ( .A(G110), .B(n637), .Z(G12) );
  NAND2_X1 U660 ( .A1(G953), .A2(G900), .ZN(n558) );
  NAND2_X1 U661 ( .A1(n559), .A2(n558), .ZN(n579) );
  NOR2_X1 U662 ( .A1(n708), .A2(n579), .ZN(n561) );
  INV_X1 U663 ( .A(KEYINPUT69), .ZN(n560) );
  XNOR2_X1 U664 ( .A(n561), .B(n560), .ZN(n562) );
  NAND2_X1 U665 ( .A1(n709), .A2(n562), .ZN(n571) );
  INV_X1 U666 ( .A(KEYINPUT104), .ZN(n565) );
  BUF_X1 U667 ( .A(n566), .Z(n567) );
  XOR2_X1 U668 ( .A(KEYINPUT90), .B(KEYINPUT36), .Z(n569) );
  INV_X1 U669 ( .A(n706), .ZN(n632) );
  XNOR2_X1 U670 ( .A(G125), .B(KEYINPUT37), .ZN(n570) );
  XNOR2_X1 U671 ( .A(n607), .B(n570), .ZN(G27) );
  XOR2_X1 U672 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n578) );
  NAND2_X1 U673 ( .A1(n721), .A2(n720), .ZN(n573) );
  INV_X1 U674 ( .A(n724), .ZN(n574) );
  NAND2_X1 U675 ( .A1(n575), .A2(n574), .ZN(n577) );
  XNOR2_X1 U676 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n576) );
  XNOR2_X1 U677 ( .A(n581), .B(n580), .ZN(n583) );
  NAND2_X1 U678 ( .A1(n583), .A2(n582), .ZN(n592) );
  XNOR2_X1 U679 ( .A(KEYINPUT86), .B(KEYINPUT46), .ZN(n585) );
  XNOR2_X1 U680 ( .A(n586), .B(n585), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n588), .A2(n587), .ZN(n759) );
  AND2_X1 U682 ( .A1(n757), .A2(n759), .ZN(n725) );
  NAND2_X1 U683 ( .A1(KEYINPUT47), .A2(n725), .ZN(n589) );
  XNOR2_X1 U684 ( .A(n589), .B(KEYINPUT84), .ZN(n594) );
  OR2_X1 U685 ( .A1(n590), .A2(n614), .ZN(n591) );
  NAND2_X1 U686 ( .A1(n759), .A2(n757), .ZN(n598) );
  INV_X1 U687 ( .A(n595), .ZN(n596) );
  NAND2_X1 U688 ( .A1(n598), .A2(n755), .ZN(n600) );
  INV_X1 U689 ( .A(KEYINPUT47), .ZN(n599) );
  NAND2_X1 U690 ( .A1(n600), .A2(n599), .ZN(n602) );
  NAND2_X1 U691 ( .A1(n755), .A2(KEYINPUT47), .ZN(n601) );
  XNOR2_X1 U692 ( .A(n604), .B(KEYINPUT75), .ZN(n605) );
  NOR2_X1 U693 ( .A1(n706), .A2(n609), .ZN(n610) );
  NAND2_X1 U694 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U695 ( .A(n612), .B(KEYINPUT43), .ZN(n613) );
  AND2_X1 U696 ( .A1(n614), .A2(n613), .ZN(n764) );
  OR2_X1 U697 ( .A1(n616), .A2(n759), .ZN(n762) );
  NAND2_X1 U698 ( .A1(n632), .A2(n630), .ZN(n617) );
  NOR2_X1 U699 ( .A1(n635), .A2(n617), .ZN(n618) );
  XOR2_X1 U700 ( .A(KEYINPUT100), .B(KEYINPUT31), .Z(n621) );
  NAND2_X1 U701 ( .A1(n619), .A2(n553), .ZN(n716) );
  NOR2_X1 U702 ( .A1(n624), .A2(n716), .ZN(n620) );
  OR2_X1 U703 ( .A1(n553), .A2(n622), .ZN(n623) );
  NOR2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n744) );
  NOR2_X1 U705 ( .A1(n625), .A2(n744), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n638), .A2(KEYINPUT44), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n630), .A2(n376), .ZN(n631) );
  NOR2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U709 ( .A(n633), .B(KEYINPUT81), .ZN(n634) );
  NOR2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n636) );
  INV_X1 U711 ( .A(n638), .ZN(n641) );
  NAND2_X1 U712 ( .A1(n641), .A2(KEYINPUT89), .ZN(n639) );
  NOR2_X1 U713 ( .A1(KEYINPUT89), .A2(KEYINPUT44), .ZN(n640) );
  NAND2_X1 U714 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U715 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n644) );
  XOR2_X1 U716 ( .A(KEYINPUT62), .B(n646), .Z(n647) );
  XNOR2_X1 U717 ( .A(n648), .B(n647), .ZN(n650) );
  INV_X1 U718 ( .A(G952), .ZN(n649) );
  NAND2_X1 U719 ( .A1(n649), .A2(G953), .ZN(n691) );
  NAND2_X1 U720 ( .A1(n650), .A2(n691), .ZN(n651) );
  XNOR2_X1 U721 ( .A(n651), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U722 ( .A(KEYINPUT94), .B(KEYINPUT59), .ZN(n652) );
  XNOR2_X1 U723 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U724 ( .A1(n656), .A2(n691), .ZN(n659) );
  XNOR2_X1 U725 ( .A(KEYINPUT119), .B(KEYINPUT60), .ZN(n657) );
  XNOR2_X1 U726 ( .A(n657), .B(KEYINPUT66), .ZN(n658) );
  XNOR2_X1 U727 ( .A(n659), .B(n658), .ZN(G60) );
  XNOR2_X1 U728 ( .A(KEYINPUT92), .B(KEYINPUT54), .ZN(n660) );
  XOR2_X1 U729 ( .A(n660), .B(KEYINPUT55), .Z(n661) );
  XNOR2_X1 U730 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U732 ( .A1(n665), .A2(n691), .ZN(n667) );
  INV_X1 U733 ( .A(KEYINPUT56), .ZN(n666) );
  XNOR2_X1 U734 ( .A(n667), .B(n666), .ZN(G51) );
  XNOR2_X1 U735 ( .A(n668), .B(KEYINPUT123), .ZN(n670) );
  XNOR2_X1 U736 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U737 ( .A(n672), .B(n671), .ZN(n676) );
  XOR2_X1 U738 ( .A(KEYINPUT124), .B(n676), .Z(n673) );
  XNOR2_X1 U739 ( .A(n674), .B(n673), .ZN(n682) );
  NOR2_X1 U740 ( .A1(n682), .A2(KEYINPUT125), .ZN(n675) );
  NOR2_X1 U741 ( .A1(n675), .A2(G953), .ZN(n681) );
  XOR2_X1 U742 ( .A(G227), .B(n676), .Z(n679) );
  NOR2_X1 U743 ( .A1(n769), .A2(KEYINPUT125), .ZN(n677) );
  NAND2_X1 U744 ( .A1(n677), .A2(G900), .ZN(n678) );
  NOR2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U746 ( .A1(n681), .A2(n680), .ZN(n686) );
  INV_X1 U747 ( .A(n682), .ZN(n684) );
  INV_X1 U748 ( .A(KEYINPUT125), .ZN(n683) );
  NOR2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U750 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U751 ( .A(KEYINPUT126), .B(n687), .Z(G72) );
  NAND2_X1 U752 ( .A1(n696), .A2(G217), .ZN(n690) );
  XNOR2_X1 U753 ( .A(n688), .B(KEYINPUT120), .ZN(n689) );
  XNOR2_X1 U754 ( .A(n690), .B(n689), .ZN(n692) );
  INV_X1 U755 ( .A(n691), .ZN(n702) );
  NOR2_X1 U756 ( .A1(n692), .A2(n702), .ZN(G66) );
  XNOR2_X1 U757 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X1 U758 ( .A1(n695), .A2(n702), .ZN(G63) );
  NAND2_X1 U759 ( .A1(n696), .A2(G469), .ZN(n701) );
  XNOR2_X1 U760 ( .A(KEYINPUT118), .B(KEYINPUT57), .ZN(n697) );
  XNOR2_X1 U761 ( .A(n697), .B(KEYINPUT58), .ZN(n698) );
  XNOR2_X1 U762 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U763 ( .A(n701), .B(n700), .ZN(n703) );
  NOR2_X1 U764 ( .A1(n703), .A2(n702), .ZN(G54) );
  BUF_X1 U765 ( .A(n704), .Z(n741) );
  NOR2_X1 U766 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U767 ( .A(n707), .B(KEYINPUT50), .ZN(n712) );
  NAND2_X1 U768 ( .A1(n376), .A2(n708), .ZN(n710) );
  XNOR2_X1 U769 ( .A(KEYINPUT49), .B(n710), .ZN(n711) );
  NOR2_X1 U770 ( .A1(n712), .A2(n711), .ZN(n714) );
  NAND2_X1 U771 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U772 ( .A(n715), .B(KEYINPUT114), .ZN(n717) );
  AND2_X1 U773 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U774 ( .A(KEYINPUT51), .B(n718), .Z(n719) );
  NOR2_X1 U775 ( .A1(n736), .A2(n719), .ZN(n728) );
  NOR2_X1 U776 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U777 ( .A(KEYINPUT115), .B(n722), .Z(n723) );
  NOR2_X1 U778 ( .A1(n724), .A2(n723), .ZN(n726) );
  NOR2_X1 U779 ( .A1(n726), .A2(n351), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n728), .A2(n349), .ZN(n729) );
  XNOR2_X1 U781 ( .A(KEYINPUT52), .B(n729), .ZN(n730) );
  XNOR2_X1 U782 ( .A(KEYINPUT116), .B(n730), .ZN(n733) );
  NAND2_X1 U783 ( .A1(G952), .A2(n731), .ZN(n732) );
  NOR2_X1 U784 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U785 ( .A1(n734), .A2(G953), .ZN(n739) );
  NOR2_X1 U786 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U787 ( .A(n737), .B(KEYINPUT117), .ZN(n738) );
  AND2_X1 U788 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U789 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U790 ( .A(KEYINPUT53), .B(n742), .Z(G75) );
  XOR2_X1 U791 ( .A(n743), .B(G101), .Z(G3) );
  INV_X1 U792 ( .A(n744), .ZN(n746) );
  NOR2_X1 U793 ( .A1(n746), .A2(n757), .ZN(n745) );
  XOR2_X1 U794 ( .A(G104), .B(n745), .Z(G6) );
  NOR2_X1 U795 ( .A1(n746), .A2(n759), .ZN(n750) );
  XOR2_X1 U796 ( .A(KEYINPUT111), .B(KEYINPUT26), .Z(n748) );
  XNOR2_X1 U797 ( .A(G107), .B(KEYINPUT27), .ZN(n747) );
  XNOR2_X1 U798 ( .A(n748), .B(n747), .ZN(n749) );
  XNOR2_X1 U799 ( .A(n750), .B(n749), .ZN(G9) );
  XOR2_X1 U800 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n753) );
  INV_X1 U801 ( .A(n759), .ZN(n751) );
  NAND2_X1 U802 ( .A1(n755), .A2(n751), .ZN(n752) );
  XNOR2_X1 U803 ( .A(n753), .B(n752), .ZN(n754) );
  XNOR2_X1 U804 ( .A(G128), .B(n754), .ZN(G30) );
  NAND2_X1 U805 ( .A1(n755), .A2(n564), .ZN(n756) );
  XNOR2_X1 U806 ( .A(n756), .B(G146), .ZN(G48) );
  NOR2_X1 U807 ( .A1(n760), .A2(n757), .ZN(n758) );
  XOR2_X1 U808 ( .A(n379), .B(n758), .Z(G15) );
  NOR2_X1 U809 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U810 ( .A(G116), .B(n761), .Z(G18) );
  INV_X1 U811 ( .A(n762), .ZN(n763) );
  XOR2_X1 U812 ( .A(G134), .B(n763), .Z(G36) );
  XOR2_X1 U813 ( .A(G140), .B(n764), .Z(G42) );
  XOR2_X1 U814 ( .A(KEYINPUT122), .B(n765), .Z(n768) );
  XNOR2_X1 U815 ( .A(n766), .B(G101), .ZN(n767) );
  XNOR2_X1 U816 ( .A(n768), .B(n767), .ZN(n771) );
  NOR2_X1 U817 ( .A1(G898), .A2(n769), .ZN(n770) );
  NOR2_X1 U818 ( .A1(n771), .A2(n770), .ZN(n779) );
  OR2_X1 U819 ( .A1(n772), .A2(G953), .ZN(n777) );
  NAND2_X1 U820 ( .A1(G953), .A2(G224), .ZN(n773) );
  XNOR2_X1 U821 ( .A(KEYINPUT61), .B(n773), .ZN(n774) );
  NAND2_X1 U822 ( .A1(n774), .A2(G898), .ZN(n775) );
  XOR2_X1 U823 ( .A(KEYINPUT121), .B(n775), .Z(n776) );
  NAND2_X1 U824 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U825 ( .A(n779), .B(n778), .ZN(G69) );
  XOR2_X1 U826 ( .A(n780), .B(G137), .Z(G39) );
  XOR2_X1 U827 ( .A(n344), .B(KEYINPUT113), .Z(n781) );
  XOR2_X1 U828 ( .A(n782), .B(G119), .Z(G21) );
  XOR2_X1 U829 ( .A(G131), .B(n783), .Z(G33) );
endmodule

