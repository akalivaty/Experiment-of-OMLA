//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT29), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT65), .A3(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  OR3_X1    g012(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n198), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n192), .A2(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n198), .A2(new_n195), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G143), .B(G146), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT66), .A3(new_n198), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n196), .A2(new_n201), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT11), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G137), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT11), .A3(G134), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(G137), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G131), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT68), .ZN(new_n217));
  INV_X1    g031(.A(G131), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n211), .A2(new_n213), .A3(new_n218), .A4(new_n214), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n217), .B1(new_n216), .B2(new_n219), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n208), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n210), .A2(G137), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n212), .A2(G134), .ZN(new_n224));
  OAI21_X1  g038(.A(G131), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n219), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n206), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n192), .A2(G146), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n230), .B1(new_n191), .B2(new_n193), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n227), .B1(new_n195), .B2(KEYINPUT1), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n229), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT69), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n226), .A2(new_n233), .A3(new_n236), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n222), .A2(KEYINPUT30), .A3(new_n235), .A4(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G113), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT2), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT2), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G113), .ZN(new_n242));
  INV_X1    g056(.A(G116), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(G119), .ZN(new_n244));
  INV_X1    g058(.A(G119), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G116), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n240), .B(new_n242), .C1(new_n244), .C2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n240), .A2(new_n242), .ZN(new_n248));
  XNOR2_X1  g062(.A(G116), .B(G119), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT67), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n247), .A2(new_n250), .A3(KEYINPUT67), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n216), .A2(new_n219), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n205), .A2(new_n207), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n196), .A2(new_n201), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n234), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT30), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n255), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n238), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n254), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT67), .B1(new_n247), .B2(new_n250), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n256), .A2(KEYINPUT68), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n266), .B1(new_n269), .B2(new_n208), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n235), .A2(new_n237), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n263), .A2(new_n272), .ZN(new_n273));
  XOR2_X1   g087(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n274));
  XNOR2_X1  g088(.A(new_n274), .B(KEYINPUT71), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT26), .B(G101), .ZN(new_n276));
  NOR2_X1   g090(.A1(G237), .A2(G953), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G210), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n276), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n275), .B(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n222), .A2(new_n255), .A3(new_n234), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT28), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n255), .B1(new_n234), .B2(new_n259), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n286), .B1(new_n270), .B2(new_n271), .ZN(new_n287));
  XOR2_X1   g101(.A(KEYINPUT73), .B(KEYINPUT28), .Z(new_n288));
  OAI21_X1  g102(.A(new_n285), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n280), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n188), .B1(new_n282), .B2(new_n291), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n283), .A2(KEYINPUT75), .A3(new_n284), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT75), .B1(new_n283), .B2(new_n284), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n222), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n235), .A2(new_n237), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n266), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n284), .B1(new_n298), .B2(new_n272), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n280), .A2(new_n188), .ZN(new_n301));
  AOI21_X1  g115(.A(G902), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n187), .B1(new_n292), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n280), .B1(new_n270), .B2(new_n271), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT31), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n263), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n305), .A2(new_n263), .A3(KEYINPUT72), .A4(new_n306), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n305), .A2(new_n263), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n289), .A2(new_n280), .B1(new_n312), .B2(KEYINPUT31), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G902), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n314), .A2(KEYINPUT32), .A3(new_n187), .A4(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(G902), .B1(new_n311), .B2(new_n313), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT32), .B1(new_n319), .B2(new_n187), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n314), .A2(new_n187), .A3(new_n315), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT32), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(KEYINPUT74), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n304), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G234), .ZN(new_n327));
  OAI21_X1  g141(.A(G217), .B1(new_n327), .B2(G902), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT76), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(G902), .ZN(new_n330));
  XOR2_X1   g144(.A(KEYINPUT22), .B(G137), .Z(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT80), .ZN(new_n332));
  INV_X1    g146(.A(G221), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n333), .A2(new_n327), .A3(G953), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n332), .B(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G140), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G125), .ZN(new_n337));
  INV_X1    g151(.A(G125), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G140), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(new_n339), .A3(KEYINPUT16), .ZN(new_n340));
  OR3_X1    g154(.A1(new_n338), .A2(KEYINPUT16), .A3(G140), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n190), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n340), .A2(new_n341), .A3(G146), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT77), .B1(new_n245), .B2(G128), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT23), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n227), .A2(G119), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT23), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(KEYINPUT77), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n245), .A2(G128), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G110), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n348), .A2(new_n351), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT24), .B(G110), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n345), .B(new_n353), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n355), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n357), .B1(new_n352), .B2(G110), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n337), .A2(new_n339), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n337), .A2(new_n339), .A3(KEYINPUT78), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(new_n190), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n358), .A2(new_n359), .A3(new_n344), .A4(new_n364), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n356), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n358), .A2(new_n344), .A3(new_n364), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT79), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n335), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n365), .A3(new_n356), .ZN(new_n370));
  INV_X1    g184(.A(new_n335), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n330), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT25), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n374), .B(new_n315), .C1(new_n369), .C2(new_n372), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n329), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n366), .A2(new_n368), .A3(new_n335), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n370), .A2(new_n371), .ZN(new_n378));
  AOI21_X1  g192(.A(G902), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(new_n374), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n373), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n360), .A2(G146), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n364), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G237), .ZN(new_n385));
  INV_X1    g199(.A(G953), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(G214), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n192), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n277), .A2(G143), .A3(G214), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g204(.A(KEYINPUT18), .B(G131), .C1(new_n390), .C2(KEYINPUT88), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT88), .ZN(new_n392));
  NAND2_X1  g206(.A1(KEYINPUT18), .A2(G131), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n388), .A2(new_n392), .A3(new_n393), .A4(new_n389), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n384), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT89), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT89), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n384), .A2(new_n391), .A3(new_n397), .A4(new_n394), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G113), .B(G122), .ZN(new_n400));
  INV_X1    g214(.A(G104), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT90), .ZN(new_n403));
  INV_X1    g217(.A(new_n344), .ZN(new_n404));
  AOI21_X1  g218(.A(G146), .B1(new_n340), .B2(new_n341), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n343), .A2(KEYINPUT90), .A3(new_n344), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT17), .ZN(new_n408));
  AOI211_X1 g222(.A(new_n408), .B(new_n218), .C1(new_n388), .C2(new_n389), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n406), .A2(new_n407), .A3(KEYINPUT91), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n390), .A2(G131), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n388), .A2(new_n218), .A3(new_n389), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n408), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT92), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n412), .A2(KEYINPUT92), .A3(new_n408), .A4(new_n413), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n411), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n409), .B1(new_n345), .B2(new_n403), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT91), .B1(new_n419), .B2(new_n407), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n399), .B(new_n402), .C1(new_n418), .C2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT93), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n406), .A2(new_n407), .A3(new_n410), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT91), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n426), .A2(new_n411), .A3(new_n416), .A4(new_n417), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n427), .A2(KEYINPUT93), .A3(new_n402), .A4(new_n399), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n404), .B1(new_n412), .B2(new_n413), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT19), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n360), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n362), .A2(new_n363), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n432), .B1(new_n433), .B2(new_n431), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n430), .B1(new_n434), .B2(G146), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n399), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n402), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n429), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n440));
  INV_X1    g254(.A(G475), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .A4(new_n315), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n423), .A2(new_n428), .B1(new_n437), .B2(new_n436), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n315), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT20), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G478), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(KEYINPUT15), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G122), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G116), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n243), .A2(G122), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G107), .ZN(new_n454));
  INV_X1    g268(.A(G107), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n227), .A2(G143), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT94), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n458), .B(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n192), .A2(G128), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n210), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(KEYINPUT13), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n457), .B(new_n462), .C1(new_n464), .C2(new_n210), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT9), .B(G234), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n467), .A2(G217), .A3(new_n386), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n456), .B(KEYINPUT95), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n210), .B1(new_n460), .B2(new_n461), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n458), .A2(new_n459), .ZN(new_n471));
  AOI21_X1  g285(.A(KEYINPUT94), .B1(new_n227), .B2(G143), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n461), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(G134), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n469), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT14), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(new_n243), .A3(G122), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT14), .B1(new_n450), .B2(G116), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n450), .A2(G116), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n480), .A2(KEYINPUT96), .A3(G107), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT96), .B1(new_n480), .B2(G107), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n465), .B(new_n468), .C1(new_n475), .C2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  OAI221_X1 g299(.A(new_n469), .B1(new_n481), .B2(new_n482), .C1(new_n474), .C2(new_n470), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n468), .B1(new_n486), .B2(new_n465), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n315), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT97), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n465), .B1(new_n475), .B2(new_n483), .ZN(new_n491));
  INV_X1    g305(.A(new_n468), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n484), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(KEYINPUT97), .A3(new_n315), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n449), .B1(new_n490), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n488), .A2(new_n449), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(G234), .A2(G237), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(G952), .A3(new_n386), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(G902), .A3(G953), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT21), .B(G898), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n499), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n402), .B1(new_n427), .B2(new_n399), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n508), .B1(new_n423), .B2(new_n428), .ZN(new_n509));
  OAI21_X1  g323(.A(G475), .B1(new_n509), .B2(G902), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n446), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(G110), .B(G140), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n386), .A2(G227), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n269), .A2(KEYINPUT85), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT85), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n267), .A2(new_n516), .A3(new_n268), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g332(.A1(KEYINPUT83), .A2(G101), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n401), .A2(G107), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT82), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n401), .A2(G107), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT3), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR4_X1   g338(.A1(new_n401), .A2(KEYINPUT82), .A3(KEYINPUT3), .A4(G107), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n520), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT81), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n527), .B(KEYINPUT3), .C1(new_n401), .C2(G107), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n455), .A2(G104), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n527), .B1(new_n530), .B2(KEYINPUT3), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n519), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT3), .B1(new_n401), .B2(G107), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT81), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n528), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n523), .A2(new_n455), .A3(G104), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT82), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n521), .A2(new_n523), .A3(new_n455), .A4(G104), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(G101), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n536), .A2(new_n540), .A3(new_n541), .A4(new_n520), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n533), .A2(KEYINPUT4), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n536), .A2(new_n540), .A3(new_n520), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT4), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n544), .A2(KEYINPUT83), .A3(new_n545), .A4(G101), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n543), .A2(new_n208), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n530), .A2(new_n520), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G101), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n542), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n233), .A2(KEYINPUT10), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n229), .B1(new_n232), .B2(new_n206), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n542), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT84), .B(KEYINPUT10), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n550), .A2(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n518), .A2(new_n547), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n553), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n233), .B1(new_n542), .B2(new_n549), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n269), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT12), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n553), .B1(new_n550), .B2(new_n233), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n560), .B1(new_n216), .B2(new_n219), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n559), .A2(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n514), .B1(new_n556), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G469), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n518), .A2(new_n547), .A3(new_n555), .ZN(new_n566));
  INV_X1    g380(.A(new_n514), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n555), .A2(new_n547), .ZN(new_n568));
  INV_X1    g382(.A(new_n269), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n566), .B(new_n567), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n564), .A2(new_n565), .A3(new_n315), .A4(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n565), .A2(new_n315), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n567), .B1(new_n556), .B2(new_n563), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n566), .B(new_n514), .C1(new_n568), .C2(new_n569), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n571), .B(new_n573), .C1(new_n565), .C2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n333), .B1(new_n467), .B2(new_n315), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(G214), .B1(G237), .B2(G902), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT5), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n239), .B1(new_n244), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n582), .A2(new_n584), .B1(new_n249), .B2(new_n248), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n542), .A2(new_n549), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT86), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT86), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n542), .A2(new_n588), .A3(new_n549), .A4(new_n585), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n543), .A2(new_n266), .A3(new_n546), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(G110), .B(G122), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(KEYINPUT6), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT6), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n592), .A2(new_n598), .A3(new_n594), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n258), .A2(new_n257), .A3(G125), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n233), .A2(new_n338), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n386), .A2(G224), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n597), .A2(new_n599), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(G210), .B1(G237), .B2(G902), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n593), .B(KEYINPUT8), .ZN(new_n607));
  INV_X1    g421(.A(new_n586), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n585), .B1(new_n542), .B2(new_n549), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n603), .A2(KEYINPUT7), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n600), .A2(new_n601), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n611), .ZN(new_n613));
  AOI21_X1  g427(.A(KEYINPUT87), .B1(new_n602), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT87), .ZN(new_n615));
  AOI211_X1 g429(.A(new_n615), .B(new_n611), .C1(new_n600), .C2(new_n601), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n610), .B(new_n612), .C1(new_n614), .C2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(G902), .B1(new_n618), .B2(new_n596), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n605), .A2(new_n606), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n606), .B1(new_n605), .B2(new_n619), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n581), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n511), .A2(new_n580), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n326), .A2(new_n382), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT98), .B(G101), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G3));
  INV_X1    g440(.A(new_n322), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n319), .A2(new_n187), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n627), .A2(new_n628), .A3(new_n381), .ZN(new_n629));
  INV_X1    g443(.A(new_n580), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(new_n631), .B(KEYINPUT99), .Z(new_n632));
  NAND2_X1  g446(.A1(new_n446), .A2(new_n510), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT33), .B1(new_n468), .B2(KEYINPUT100), .ZN(new_n634));
  OR2_X1    g448(.A1(new_n494), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n494), .A2(new_n634), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n447), .A2(G902), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT101), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT101), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n635), .A2(new_n640), .A3(new_n636), .A4(new_n637), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n490), .A2(new_n447), .A3(new_n495), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n639), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n633), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n621), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n605), .A2(new_n606), .A3(new_n619), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n506), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(new_n648), .A3(new_n581), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n632), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT102), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT34), .B(G104), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  NAND2_X1  g468(.A1(new_n510), .A2(KEYINPUT103), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n656), .B(G475), .C1(new_n509), .C2(G902), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n446), .A2(new_n499), .A3(new_n655), .A4(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n649), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n632), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NOR2_X1   g476(.A1(new_n335), .A2(KEYINPUT36), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(new_n368), .A3(new_n366), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n370), .B1(KEYINPUT36), .B2(new_n335), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n330), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n380), .ZN(new_n669));
  INV_X1    g483(.A(new_n329), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n379), .B2(new_n374), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n668), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n627), .A2(new_n628), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n623), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  XNOR2_X1  g490(.A(KEYINPUT104), .B(G900), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n502), .B1(new_n677), .B2(new_n504), .ZN(new_n678));
  OAI22_X1  g492(.A1(new_n376), .A2(new_n380), .B1(new_n667), .B2(new_n666), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n581), .B(new_n679), .C1(new_n620), .C2(new_n621), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n658), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n326), .A2(new_n630), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT105), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n322), .A2(new_n323), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n317), .A3(new_n316), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n324), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n580), .B1(new_n686), .B2(new_n304), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(new_n688), .A3(new_n681), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  XOR2_X1   g505(.A(new_n678), .B(KEYINPUT39), .Z(new_n692));
  NAND2_X1  g506(.A1(new_n630), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n693), .B(KEYINPUT40), .Z(new_n694));
  AOI21_X1  g508(.A(new_n290), .B1(new_n298), .B2(new_n272), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n263), .B2(new_n305), .ZN(new_n696));
  OAI21_X1  g510(.A(G472), .B1(new_n696), .B2(G902), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n686), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n647), .B(KEYINPUT38), .ZN(new_n699));
  INV_X1    g513(.A(new_n508), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n429), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n441), .B1(new_n701), .B2(new_n315), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n445), .B2(new_n442), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n496), .A2(new_n498), .ZN(new_n704));
  INV_X1    g518(.A(new_n581), .ZN(new_n705));
  NOR4_X1   g519(.A1(new_n703), .A2(new_n704), .A3(new_n705), .A4(new_n679), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n694), .A2(new_n698), .A3(new_n699), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G143), .ZN(G45));
  INV_X1    g522(.A(new_n678), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n633), .A2(new_n643), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n680), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n687), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G146), .ZN(G48));
  NAND3_X1  g527(.A1(new_n564), .A2(new_n315), .A3(new_n570), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(G469), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n571), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n578), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n326), .A2(new_n650), .A3(new_n382), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT41), .B(G113), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NAND4_X1  g534(.A1(new_n326), .A2(new_n659), .A3(new_n382), .A4(new_n717), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  NAND3_X1  g536(.A1(new_n703), .A2(new_n507), .A3(new_n679), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n717), .A2(new_n647), .A3(new_n581), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n326), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT106), .B(G119), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G21));
  NOR3_X1   g542(.A1(new_n703), .A2(new_n622), .A3(new_n704), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n312), .A2(KEYINPUT31), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n280), .B1(new_n295), .B2(new_n299), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n311), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n187), .A2(new_n315), .ZN(new_n733));
  OAI22_X1  g547(.A1(new_n732), .A2(new_n733), .B1(new_n319), .B2(new_n187), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n715), .A2(new_n648), .A3(new_n579), .A4(new_n571), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n734), .A2(new_n381), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n729), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  OAI221_X1 g552(.A(new_n679), .B1(new_n319), .B2(new_n187), .C1(new_n732), .C2(new_n733), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n710), .A2(new_n724), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n338), .ZN(G27));
  OR2_X1    g555(.A1(new_n316), .A2(KEYINPUT110), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n316), .A2(KEYINPUT110), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n742), .A2(new_n304), .A3(new_n684), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n382), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT42), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n620), .A2(new_n621), .A3(new_n705), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n571), .A2(new_n573), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n575), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n555), .ZN(new_n752));
  INV_X1    g566(.A(new_n547), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n269), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(KEYINPUT107), .A3(new_n566), .A4(new_n514), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n751), .A2(G469), .A3(new_n574), .A4(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n748), .B1(new_n749), .B2(new_n756), .ZN(new_n757));
  AND4_X1   g571(.A1(new_n748), .A2(new_n756), .A3(new_n571), .A4(new_n573), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n579), .B(new_n747), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NOR4_X1   g573(.A1(new_n745), .A2(new_n746), .A3(new_n710), .A4(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n710), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n645), .A2(new_n579), .A3(new_n581), .A4(new_n646), .ZN(new_n763));
  INV_X1    g577(.A(new_n757), .ZN(new_n764));
  INV_X1    g578(.A(new_n758), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n326), .A2(new_n762), .A3(new_n382), .A4(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n746), .B1(new_n767), .B2(new_n768), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n761), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G131), .ZN(G33));
  NOR2_X1   g587(.A1(new_n658), .A2(new_n678), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n326), .A2(new_n382), .A3(new_n774), .A4(new_n766), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  INV_X1    g590(.A(new_n747), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n679), .B1(new_n627), .B2(new_n628), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT112), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n703), .A2(new_n643), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT43), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT43), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n703), .A2(new_n782), .A3(new_n643), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n777), .B1(new_n785), .B2(KEYINPUT44), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n565), .B1(new_n576), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n751), .A2(KEYINPUT45), .A3(new_n574), .A4(new_n755), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n572), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OR3_X1    g604(.A1(new_n790), .A2(KEYINPUT111), .A3(KEYINPUT46), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT111), .B1(new_n790), .B2(KEYINPUT46), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(KEYINPUT46), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n791), .A2(new_n571), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n579), .A3(new_n692), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n786), .B(new_n796), .C1(KEYINPUT44), .C2(new_n785), .ZN(new_n797));
  XOR2_X1   g611(.A(KEYINPUT113), .B(G137), .Z(new_n798));
  XNOR2_X1  g612(.A(new_n797), .B(new_n798), .ZN(G39));
  NAND2_X1  g613(.A1(new_n794), .A2(new_n579), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT47), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n801), .A2(new_n802), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n794), .A2(new_n579), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n303), .B1(new_n685), .B2(new_n324), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n710), .A2(new_n382), .A3(new_n777), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n764), .A2(new_n765), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n679), .A2(new_n578), .A3(new_n678), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n698), .A2(new_n729), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n740), .B1(new_n687), .B2(new_n711), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n688), .B1(new_n687), .B2(new_n681), .ZN(new_n817));
  INV_X1    g631(.A(new_n680), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n655), .A2(new_n657), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n704), .B1(new_n445), .B2(new_n442), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n709), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n808), .A2(new_n821), .A3(KEYINPUT105), .A4(new_n580), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n815), .B(new_n816), .C1(new_n817), .C2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n690), .A2(KEYINPUT52), .A3(new_n815), .A4(new_n816), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n623), .A2(new_n673), .B1(new_n729), .B2(new_n736), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n703), .A2(new_n499), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n644), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n649), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n830), .A2(new_n831), .A3(new_n630), .A4(new_n629), .ZN(new_n832));
  AND4_X1   g646(.A1(new_n624), .A2(new_n828), .A3(new_n726), .A4(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n718), .A2(new_n721), .ZN(new_n834));
  INV_X1    g648(.A(new_n739), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n762), .A2(new_n766), .A3(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n672), .A2(new_n499), .A3(new_n678), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n446), .A2(new_n819), .A3(new_n747), .A4(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n326), .A2(new_n838), .A3(new_n630), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n775), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n772), .A2(new_n833), .A3(new_n834), .A4(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n812), .B1(new_n827), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n825), .A2(new_n844), .A3(new_n826), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n808), .A2(new_n759), .A3(new_n710), .A4(new_n381), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT42), .B1(new_n846), .B2(KEYINPUT109), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n760), .B1(new_n847), .B2(new_n769), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n833), .A2(new_n840), .A3(new_n834), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n740), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n712), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(new_n689), .B2(new_n683), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(KEYINPUT115), .A3(KEYINPUT52), .A4(new_n815), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n845), .A2(new_n850), .A3(new_n854), .A4(KEYINPUT53), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n842), .A2(new_n843), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT116), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT53), .B1(new_n827), .B2(new_n841), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n845), .A2(new_n850), .A3(new_n854), .A4(new_n812), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT54), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n842), .A2(new_n843), .A3(new_n855), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n857), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n686), .A2(new_n697), .ZN(new_n867));
  NOR4_X1   g681(.A1(new_n763), .A2(new_n381), .A3(new_n501), .A4(new_n716), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI211_X1 g683(.A(G952), .B(new_n386), .C1(new_n869), .C2(new_n644), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n734), .A2(new_n381), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n781), .A2(new_n502), .A3(new_n871), .A4(new_n783), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n724), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n763), .A2(new_n716), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n781), .A2(new_n502), .A3(new_n783), .A4(new_n875), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT118), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT48), .ZN(new_n878));
  INV_X1    g692(.A(new_n745), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n878), .B1(new_n877), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n874), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n633), .A2(new_n643), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n867), .A2(new_n868), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT119), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n867), .A2(new_n887), .A3(new_n868), .A4(new_n884), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n877), .A2(new_n835), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n784), .A2(new_n501), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n717), .A2(new_n705), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n699), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n890), .A2(new_n892), .A3(KEYINPUT50), .A4(new_n871), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT50), .ZN(new_n894));
  INV_X1    g708(.A(new_n892), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n894), .B1(new_n895), .B2(new_n872), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n889), .A2(KEYINPUT51), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n872), .A2(new_n777), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n716), .A2(new_n579), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n899), .B1(new_n807), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n882), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g716(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n877), .A2(new_n835), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n886), .A2(new_n888), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n904), .A2(new_n905), .A3(new_n897), .A4(KEYINPUT120), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n901), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT120), .B1(new_n889), .B2(new_n897), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n903), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n902), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT121), .ZN(new_n911));
  OAI22_X1  g725(.A1(new_n866), .A2(new_n911), .B1(G952), .B2(G953), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n716), .B(KEYINPUT49), .Z(new_n913));
  NAND4_X1  g727(.A1(new_n913), .A2(new_n382), .A3(new_n579), .A4(new_n581), .ZN(new_n914));
  OR3_X1    g728(.A1(new_n914), .A2(new_n699), .A3(new_n780), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n912), .B1(new_n698), .B2(new_n915), .ZN(G75));
  NAND2_X1  g730(.A1(new_n842), .A2(new_n855), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(G210), .A3(G902), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT56), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n597), .A2(new_n599), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(new_n604), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n921), .A2(KEYINPUT55), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(KEYINPUT55), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n919), .A2(KEYINPUT122), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n918), .A2(new_n919), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n925), .B1(new_n918), .B2(new_n919), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n386), .A2(G952), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(G51));
  NAND2_X1  g743(.A1(new_n788), .A2(new_n789), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT123), .ZN(new_n931));
  AOI211_X1 g745(.A(new_n315), .B(new_n931), .C1(new_n842), .C2(new_n855), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n572), .B(KEYINPUT57), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n843), .B1(new_n842), .B2(new_n855), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n933), .B1(new_n856), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n564), .A2(new_n570), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n932), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(KEYINPUT124), .B1(new_n938), .B2(new_n928), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT124), .ZN(new_n940));
  INV_X1    g754(.A(new_n928), .ZN(new_n941));
  AND4_X1   g755(.A1(KEYINPUT53), .A2(new_n845), .A3(new_n850), .A4(new_n854), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n825), .A2(new_n826), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT53), .B1(new_n850), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(KEYINPUT54), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n863), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n936), .B1(new_n946), .B2(new_n933), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n940), .B(new_n941), .C1(new_n947), .C2(new_n932), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n939), .A2(new_n948), .ZN(G54));
  AND4_X1   g763(.A1(KEYINPUT58), .A2(new_n917), .A3(G475), .A4(G902), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n941), .B1(new_n950), .B2(new_n439), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n439), .B2(new_n950), .ZN(G60));
  INV_X1    g766(.A(new_n946), .ZN(new_n953));
  XNOR2_X1  g767(.A(KEYINPUT125), .B(KEYINPUT59), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n447), .A2(new_n315), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n635), .A2(new_n636), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n941), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n866), .A2(new_n956), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n635), .A2(new_n636), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(G63));
  NAND2_X1  g775(.A1(G217), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT60), .Z(new_n963));
  NAND2_X1  g777(.A1(new_n917), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n369), .A2(new_n372), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n966), .B(new_n941), .C1(new_n666), .C2(new_n964), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT61), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(G66));
  NAND2_X1  g783(.A1(new_n833), .A2(new_n834), .ZN(new_n970));
  NAND2_X1  g784(.A1(G224), .A2(G953), .ZN(new_n971));
  OAI22_X1  g785(.A1(new_n970), .A2(G953), .B1(new_n505), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n920), .B1(G898), .B2(new_n386), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT126), .Z(new_n974));
  XNOR2_X1  g788(.A(new_n972), .B(new_n974), .ZN(G69));
  NAND2_X1  g789(.A1(new_n853), .A2(new_n707), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT62), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n693), .A2(new_n777), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n326), .A2(new_n978), .A3(new_n382), .A4(new_n830), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n797), .A2(new_n810), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n386), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n260), .A2(new_n261), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n238), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(new_n434), .Z(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT127), .Z(new_n985));
  NAND2_X1  g799(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n984), .B1(G900), .B2(G953), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n796), .A2(new_n729), .A3(new_n879), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n797), .A2(new_n775), .A3(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n989), .A2(new_n772), .A3(new_n810), .A4(new_n853), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n987), .B1(new_n990), .B2(G953), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n986), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n386), .B1(G227), .B2(G900), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n992), .B(new_n993), .ZN(G72));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT63), .Z(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n990), .B2(new_n970), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n928), .B1(new_n997), .B2(new_n282), .ZN(new_n998));
  INV_X1    g812(.A(new_n273), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n977), .A2(new_n970), .A3(new_n980), .ZN(new_n1000));
  INV_X1    g814(.A(new_n996), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n290), .B(new_n999), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n999), .A2(new_n280), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1001), .B1(new_n1004), .B2(new_n312), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1003), .B1(new_n861), .B2(new_n1005), .ZN(G57));
endmodule


