//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n202), .A3(new_n206), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G226gat), .A2(G233gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT26), .ZN(new_n218));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT64), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(G169gat), .A3(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT27), .B(G183gat), .ZN(new_n225));
  INV_X1    g024(.A(G190gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(KEYINPUT28), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n228));
  AOI21_X1  g027(.A(G190gat), .B1(new_n228), .B2(KEYINPUT27), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT27), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT28), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT68), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n227), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI211_X1 g033(.A(KEYINPUT68), .B(KEYINPUT28), .C1(new_n229), .C2(new_n231), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n216), .B(new_n224), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT24), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n216), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT66), .ZN(new_n239));
  OR2_X1    g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n216), .A2(new_n242), .A3(new_n237), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n239), .A2(new_n240), .A3(new_n241), .A4(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT23), .ZN(new_n246));
  INV_X1    g045(.A(G169gat), .ZN(new_n247));
  INV_X1    g046(.A(G176gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n245), .A2(new_n249), .B1(new_n220), .B2(new_n222), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n244), .A2(KEYINPUT25), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n238), .A2(new_n240), .A3(new_n241), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT25), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n251), .B1(new_n253), .B2(KEYINPUT65), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n245), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n252), .A2(new_n255), .A3(new_n223), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT25), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n256), .A2(KEYINPUT65), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n236), .B1(new_n254), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT29), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n215), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n256), .A2(new_n257), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT65), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n265), .A2(new_n258), .A3(new_n251), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n214), .B1(new_n266), .B2(new_n236), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n213), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n260), .A2(new_n215), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT29), .B1(new_n266), .B2(new_n236), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n269), .B(new_n212), .C1(new_n270), .C2(new_n215), .ZN(new_n271));
  XNOR2_X1  g070(.A(G8gat), .B(G36gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(G64gat), .B(G92gat), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n272), .B(new_n273), .Z(new_n274));
  NAND3_X1  g073(.A1(new_n268), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT30), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G225gat), .A2(G233gat), .ZN(new_n278));
  OR2_X1    g077(.A1(KEYINPUT73), .A2(G141gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(KEYINPUT73), .A2(G141gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(G148gat), .A3(new_n280), .ZN(new_n281));
  OR2_X1    g080(.A1(KEYINPUT74), .A2(G148gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(KEYINPUT74), .A2(G148gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(G141gat), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  OR3_X1    g084(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(G141gat), .A2(G148gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n290), .A2(KEYINPUT2), .ZN(new_n291));
  NAND2_X1  g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G155gat), .ZN(new_n294));
  INV_X1    g093(.A(G162gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n287), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n289), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT3), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT3), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n289), .A2(new_n300), .A3(new_n297), .ZN(new_n301));
  INV_X1    g100(.A(G120gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G113gat), .ZN(new_n303));
  INV_X1    g102(.A(G113gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G120gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT1), .ZN(new_n307));
  INV_X1    g106(.A(G134gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G127gat), .ZN(new_n309));
  INV_X1    g108(.A(G127gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G134gat), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n306), .A2(new_n307), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n309), .A2(new_n311), .A3(new_n307), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT69), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n316), .B1(new_n302), .B2(G113gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n304), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n303), .A3(new_n318), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n314), .A2(new_n315), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n315), .B1(new_n314), .B2(new_n319), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n313), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n299), .A2(new_n301), .A3(new_n322), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n322), .A2(KEYINPUT4), .A3(new_n298), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT4), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n314), .A2(new_n319), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT70), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n314), .A2(new_n319), .A3(new_n315), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n312), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n281), .A2(new_n284), .B1(new_n287), .B2(new_n286), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n296), .A2(new_n287), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n331), .B1(new_n292), .B2(new_n291), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n325), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n278), .B(new_n323), .C1(new_n324), .C2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT5), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n322), .A2(new_n298), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n333), .B(new_n313), .C1(new_n321), .C2(new_n320), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n278), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G1gat), .B(G29gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n343), .B(KEYINPUT0), .ZN(new_n344));
  XNOR2_X1  g143(.A(G57gat), .B(G85gat), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n344), .B(new_n345), .Z(new_n346));
  NAND2_X1  g145(.A1(new_n338), .A2(KEYINPUT4), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n329), .A2(new_n325), .A3(new_n333), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n349), .A2(new_n336), .A3(new_n278), .A4(new_n323), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n342), .A2(new_n346), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT6), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n346), .B1(new_n342), .B2(new_n350), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n342), .A2(new_n350), .ZN(new_n356));
  INV_X1    g155(.A(new_n346), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(KEYINPUT6), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n277), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  AND4_X1   g159(.A1(KEYINPUT30), .A2(new_n268), .A3(new_n271), .A4(new_n274), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n274), .B1(new_n268), .B2(new_n271), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT72), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n362), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT72), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n268), .A2(KEYINPUT30), .A3(new_n271), .A4(new_n274), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT75), .B1(new_n360), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n277), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n356), .A2(new_n357), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(new_n352), .A3(new_n351), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n370), .B1(new_n372), .B2(new_n358), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT75), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n373), .A2(new_n374), .A3(new_n367), .A4(new_n363), .ZN(new_n375));
  XNOR2_X1  g174(.A(G15gat), .B(G43gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(G71gat), .B(G99gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n236), .B(new_n329), .C1(new_n254), .C2(new_n259), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT71), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n266), .A2(KEYINPUT71), .A3(new_n329), .A4(new_n236), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n260), .A2(new_n322), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G227gat), .A2(G233gat), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT33), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n378), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n329), .B1(new_n266), .B2(new_n236), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n380), .B2(new_n379), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT34), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n391), .A2(new_n392), .A3(new_n385), .A4(new_n382), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n381), .A2(new_n383), .A3(new_n385), .A4(new_n382), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT34), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n389), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n387), .A2(KEYINPUT32), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT33), .B1(new_n384), .B2(new_n386), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n395), .B(new_n393), .C1(new_n400), .C2(new_n378), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n397), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n399), .B1(new_n397), .B2(new_n401), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G78gat), .B(G106gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(G22gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(KEYINPUT31), .B(G50gat), .Z(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT29), .B1(new_n210), .B2(new_n211), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n298), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(G228gat), .ZN(new_n412));
  INV_X1    g211(.A(G233gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(new_n299), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT77), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n330), .A2(new_n332), .A3(KEYINPUT3), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n417), .B1(new_n418), .B2(KEYINPUT29), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n301), .A2(KEYINPUT77), .A3(new_n261), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n420), .A3(new_n213), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n421), .A2(KEYINPUT78), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n301), .A2(new_n261), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n212), .B1(new_n424), .B2(new_n417), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n423), .B1(new_n425), .B2(new_n420), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n416), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT76), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n410), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n300), .B1(new_n410), .B2(new_n428), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n298), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n424), .A2(new_n213), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n414), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n409), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n421), .A2(KEYINPUT78), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n425), .A2(new_n423), .A3(new_n420), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n415), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n438), .A2(new_n433), .A3(new_n408), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n407), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n427), .A2(new_n434), .A3(new_n409), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n408), .B1(new_n438), .B2(new_n433), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n442), .A3(new_n406), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n369), .A2(new_n375), .A3(new_n404), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT35), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n404), .A2(KEYINPUT80), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT80), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n449), .B1(new_n402), .B2(new_n403), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n444), .A2(KEYINPUT35), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n361), .A2(new_n362), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n277), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n453), .B1(new_n358), .B2(new_n372), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n448), .A2(new_n450), .A3(new_n451), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n397), .A2(new_n401), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n398), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n397), .A2(new_n399), .A3(new_n401), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(KEYINPUT36), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT36), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n460), .B1(new_n402), .B2(new_n403), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT40), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n323), .B1(new_n324), .B2(new_n334), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT39), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(new_n464), .A3(new_n340), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n346), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT39), .B1(new_n339), .B2(new_n340), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n467), .B1(new_n340), .B2(new_n463), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n462), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n371), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n466), .A2(new_n468), .A3(new_n462), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n444), .B1(new_n453), .B2(new_n472), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n372), .A2(new_n358), .A3(new_n275), .ZN(new_n474));
  INV_X1    g273(.A(new_n274), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n475), .A2(KEYINPUT37), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n362), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT38), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n268), .A2(new_n271), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT37), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT79), .B(new_n475), .C1(new_n479), .C2(KEYINPUT37), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n477), .A2(new_n478), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n478), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n480), .B1(new_n362), .B2(new_n476), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n474), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n459), .A2(new_n461), .B1(new_n473), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n375), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n363), .A2(new_n367), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n374), .B1(new_n489), .B2(new_n373), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n444), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n447), .A2(new_n455), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G113gat), .B(G141gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(G169gat), .B(G197gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  XOR2_X1   g294(.A(KEYINPUT81), .B(KEYINPUT11), .Z(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(KEYINPUT12), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G43gat), .B(G50gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT15), .ZN(new_n501));
  NOR3_X1   g300(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(KEYINPUT84), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT82), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n503), .B1(KEYINPUT83), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n506), .A2(KEYINPUT83), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT85), .B(G36gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G29gat), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n501), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n502), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n500), .A2(KEYINPUT86), .A3(KEYINPUT15), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT15), .B1(new_n500), .B2(KEYINPUT86), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n511), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT17), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n518), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT17), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n507), .A2(new_n508), .B1(G29gat), .B2(new_n510), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n520), .B(new_n521), .C1(new_n522), .C2(new_n501), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  AND2_X1   g324(.A1(KEYINPUT87), .A2(G1gat), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT16), .B1(KEYINPUT87), .B2(G1gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n528), .B(KEYINPUT88), .C1(G1gat), .C2(new_n525), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(G8gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n530), .B1(new_n512), .B2(new_n518), .ZN(new_n533));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT89), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT18), .B1(new_n532), .B2(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n535), .B(KEYINPUT13), .Z(new_n539));
  NAND2_X1  g338(.A1(new_n509), .A2(new_n511), .ZN(new_n540));
  INV_X1    g339(.A(new_n501), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n531), .B1(new_n542), .B2(new_n520), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n512), .A2(new_n530), .A3(new_n518), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n539), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n530), .B1(new_n519), .B2(new_n523), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n533), .A2(KEYINPUT18), .A3(new_n535), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n499), .B1(new_n538), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT90), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n546), .A2(new_n547), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT18), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(new_n546), .B2(new_n536), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n551), .A2(new_n553), .A3(new_n545), .A4(new_n498), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n549), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  OAI211_X1 g354(.A(KEYINPUT90), .B(new_n499), .C1(new_n538), .C2(new_n548), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n492), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT95), .ZN(new_n559));
  XNOR2_X1  g358(.A(G183gat), .B(G211gat), .ZN(new_n560));
  OR2_X1    g359(.A1(G57gat), .A2(G64gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(G57gat), .A2(G64gat), .ZN(new_n562));
  AND2_X1   g361(.A1(G71gat), .A2(G78gat), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n561), .B(new_n562), .C1(new_n563), .C2(KEYINPUT9), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT91), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n564), .B1(new_n565), .B2(new_n563), .ZN(new_n566));
  NOR2_X1   g365(.A1(G71gat), .A2(G78gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n568), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n570), .B(new_n564), .C1(new_n565), .C2(new_n563), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(KEYINPUT21), .ZN(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n574), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n575), .A2(new_n310), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n310), .B1(new_n575), .B2(new_n576), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n560), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OR3_X1    g378(.A1(new_n577), .A2(new_n578), .A3(new_n560), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n530), .B1(KEYINPUT21), .B2(new_n572), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT92), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(new_n294), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT92), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n581), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(new_n584), .ZN(new_n589));
  AND4_X1   g388(.A1(new_n579), .A2(new_n580), .A3(new_n586), .A4(new_n589), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n579), .A2(new_n580), .B1(new_n586), .B2(new_n589), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(G190gat), .B(G218gat), .Z(new_n594));
  NAND2_X1  g393(.A1(G85gat), .A2(G92gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT7), .ZN(new_n596));
  XOR2_X1   g395(.A(G99gat), .B(G106gat), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G99gat), .A2(G106gat), .ZN(new_n599));
  INV_X1    g398(.A(G85gat), .ZN(new_n600));
  INV_X1    g399(.A(G92gat), .ZN(new_n601));
  AOI22_X1  g400(.A1(KEYINPUT8), .A2(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n596), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n598), .B1(new_n596), .B2(new_n602), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n605), .B1(new_n519), .B2(new_n523), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n605), .B1(new_n512), .B2(new_n518), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT41), .ZN(new_n608));
  NAND2_X1  g407(.A1(G232gat), .A2(G233gat), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n594), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NOR3_X1   g411(.A1(new_n606), .A2(new_n610), .A3(new_n594), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT94), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n609), .A2(new_n608), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n615), .B(KEYINPUT93), .Z(new_n616));
  XOR2_X1   g415(.A(G134gat), .B(G162gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  OAI22_X1  g417(.A1(new_n612), .A2(new_n613), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n613), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n618), .B(new_n614), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(new_n611), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n559), .B1(new_n593), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n623), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(new_n592), .A3(KEYINPUT95), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n605), .A2(new_n572), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT10), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n569), .B(new_n571), .C1(new_n603), .C2(new_n604), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n605), .A2(new_n572), .A3(KEYINPUT10), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G230gat), .A2(G233gat), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n633), .B1(new_n627), .B2(new_n629), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT96), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(G176gat), .B(G204gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n640), .B(new_n641), .Z(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n635), .A2(new_n638), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n642), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n633), .B(KEYINPUT97), .Z(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n630), .B2(new_n631), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n646), .B1(new_n648), .B2(new_n636), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n624), .A2(new_n626), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n558), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n372), .A2(new_n358), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT98), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(G1gat), .ZN(G1324gat));
  INV_X1    g457(.A(new_n453), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT99), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(G8gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(G8gat), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n663), .B1(new_n664), .B2(new_n660), .ZN(new_n665));
  MUX2_X1   g464(.A(new_n663), .B(new_n665), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g465(.A1(new_n461), .A2(new_n459), .ZN(new_n667));
  OAI21_X1  g466(.A(G15gat), .B1(new_n653), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n448), .A2(new_n450), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n669), .A2(G15gat), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n668), .B1(new_n653), .B2(new_n670), .ZN(G1326gat));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n444), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT100), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT43), .B(G22gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  NAND3_X1  g474(.A1(new_n593), .A2(new_n623), .A3(new_n651), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT101), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n558), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n656), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n678), .A2(G29gat), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT45), .Z(new_n681));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n557), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n555), .A2(KEYINPUT102), .A3(new_n556), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n650), .B(KEYINPUT103), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n593), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n473), .A2(new_n486), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n667), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n445), .B1(new_n369), .B2(new_n375), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n491), .A2(new_n487), .A3(KEYINPUT104), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n447), .A2(new_n455), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n447), .A2(KEYINPUT105), .A3(new_n455), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n694), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT106), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n694), .A2(new_n697), .A3(new_n701), .A4(new_n698), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n623), .A2(KEYINPUT107), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n619), .A2(new_n622), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(KEYINPUT44), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n700), .A2(new_n702), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT44), .B1(new_n492), .B2(new_n625), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n687), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n710), .A2(new_n656), .ZN(new_n711));
  INV_X1    g510(.A(G29gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n681), .B1(new_n711), .B2(new_n712), .ZN(G1328gat));
  NOR3_X1   g512(.A1(new_n678), .A2(new_n659), .A3(new_n510), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n710), .A2(new_n453), .ZN(new_n717));
  INV_X1    g516(.A(new_n510), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(G1329gat));
  INV_X1    g518(.A(new_n667), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n710), .A2(G43gat), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n678), .A2(new_n669), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(G43gat), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1330gat));
  NOR3_X1   g524(.A1(new_n678), .A2(G50gat), .A3(new_n445), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n444), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(G50gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g528(.A1(new_n700), .A2(new_n702), .ZN(new_n730));
  INV_X1    g529(.A(new_n685), .ZN(new_n731));
  INV_X1    g530(.A(new_n686), .ZN(new_n732));
  AND4_X1   g531(.A1(new_n624), .A2(new_n731), .A3(new_n626), .A4(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n730), .A2(new_n656), .A3(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT110), .B(G57gat), .Z(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1332gat));
  NAND3_X1  g535(.A1(new_n730), .A2(new_n453), .A3(new_n733), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT49), .B(G64gat), .Z(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(G1333gat));
  NAND3_X1  g539(.A1(new_n730), .A2(new_n720), .A3(new_n733), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G71gat), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n669), .A2(G71gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n730), .A2(new_n733), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT50), .Z(G1334gat));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n444), .A3(new_n733), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g547(.A1(new_n708), .A2(new_n709), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n731), .A2(new_n593), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n651), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT111), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n753));
  INV_X1    g552(.A(new_n751), .ZN(new_n754));
  AOI211_X1 g553(.A(new_n753), .B(new_n754), .C1(new_n708), .C2(new_n709), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n600), .B1(new_n756), .B2(new_n656), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n750), .A2(new_n625), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n699), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n761), .A2(new_n600), .A3(new_n650), .A4(new_n656), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT112), .B1(new_n757), .B2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n752), .A2(new_n755), .A3(new_n679), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n765), .B(new_n762), .C1(new_n766), .C2(new_n600), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n767), .ZN(G1336gat));
  AND2_X1   g567(.A1(new_n761), .A2(new_n732), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n659), .A2(G92gat), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n749), .A2(new_n751), .ZN(new_n773));
  OAI21_X1  g572(.A(G92gat), .B1(new_n773), .B2(new_n659), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT52), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n752), .A2(new_n755), .ZN(new_n776));
  OAI211_X1 g575(.A(KEYINPUT52), .B(G92gat), .C1(new_n776), .C2(new_n659), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n778), .B1(new_n769), .B2(new_n771), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n775), .B1(new_n777), .B2(new_n779), .ZN(G1337gat));
  OAI21_X1  g579(.A(G99gat), .B1(new_n776), .B2(new_n667), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n669), .A2(G99gat), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n761), .A2(new_n650), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(G1338gat));
  OAI21_X1  g583(.A(G106gat), .B1(new_n773), .B2(new_n445), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n445), .A2(G106gat), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n761), .A2(new_n732), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n785), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n788), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n756), .A2(new_n444), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n791), .B2(G106gat), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n789), .B1(new_n792), .B2(new_n786), .ZN(G1339gat));
  NAND3_X1  g592(.A1(new_n630), .A2(new_n631), .A3(new_n647), .ZN(new_n794));
  OAI211_X1 g593(.A(KEYINPUT54), .B(new_n794), .C1(new_n632), .C2(new_n634), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n642), .B1(new_n648), .B2(new_n796), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n795), .A2(KEYINPUT55), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT55), .B1(new_n795), .B2(new_n797), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n798), .A2(new_n799), .A3(new_n644), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n683), .B2(new_n684), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n535), .B1(new_n532), .B2(new_n533), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n543), .A2(new_n544), .A3(new_n539), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n497), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n650), .A2(new_n554), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n706), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n805), .A2(new_n554), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n703), .A2(new_n809), .A3(new_n705), .A4(new_n800), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n592), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n652), .A2(new_n731), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n444), .ZN(new_n814));
  INV_X1    g613(.A(new_n669), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n679), .A2(new_n453), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n817), .A2(new_n304), .A3(new_n557), .ZN(new_n818));
  INV_X1    g617(.A(new_n816), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n813), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n402), .A2(new_n444), .A3(new_n403), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n821), .A3(new_n685), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n818), .B1(new_n304), .B2(new_n822), .ZN(G1340gat));
  OAI21_X1  g622(.A(G120gat), .B1(new_n817), .B2(new_n686), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n820), .A2(new_n821), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n650), .A2(new_n302), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT114), .ZN(G1341gat));
  OAI21_X1  g627(.A(G127gat), .B1(new_n817), .B2(new_n593), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n592), .A2(new_n310), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n825), .B2(new_n830), .ZN(G1342gat));
  NOR3_X1   g630(.A1(new_n825), .A2(G134gat), .A3(new_n625), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n833), .A2(KEYINPUT56), .ZN(new_n834));
  OAI21_X1  g633(.A(G134gat), .B1(new_n817), .B2(new_n625), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(KEYINPUT56), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(G1343gat));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT58), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n445), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n555), .A2(new_n556), .A3(new_n800), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n806), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n625), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n623), .B1(new_n843), .B2(new_n806), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT115), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(new_n810), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n842), .B1(new_n850), .B2(new_n593), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n810), .B1(new_n848), .B2(KEYINPUT115), .ZN(new_n852));
  AOI211_X1 g651(.A(new_n846), .B(new_n623), .C1(new_n843), .C2(new_n806), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n842), .B(new_n593), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n652), .A2(new_n731), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n841), .B1(new_n851), .B2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(KEYINPUT117), .B(new_n841), .C1(new_n851), .C2(new_n856), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n840), .B1(new_n813), .B2(new_n445), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n819), .A2(new_n720), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n685), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n279), .A2(new_n280), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n720), .A2(new_n445), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n820), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n557), .A2(G141gat), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n839), .B1(new_n866), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n839), .ZN(new_n873));
  INV_X1    g672(.A(new_n557), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n862), .A2(new_n874), .A3(new_n863), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n873), .B1(new_n865), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n838), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n865), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT58), .B1(new_n869), .B2(new_n870), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n864), .A2(new_n865), .B1(new_n869), .B2(new_n870), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n880), .B(KEYINPUT118), .C1(new_n839), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n877), .A2(new_n882), .ZN(G1344gat));
  NAND2_X1  g682(.A1(new_n282), .A2(new_n283), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n868), .A2(new_n884), .A3(new_n651), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT119), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n862), .A2(new_n863), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n650), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n811), .A2(new_n812), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n841), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n809), .A2(new_n623), .A3(new_n800), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n592), .B1(new_n845), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n894), .B1(new_n557), .B2(new_n652), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n840), .B1(new_n895), .B2(new_n445), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g697(.A(KEYINPUT121), .B(new_n840), .C1(new_n895), .C2(new_n445), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n892), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n650), .B1(new_n863), .B2(KEYINPUT120), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n901), .B1(KEYINPUT120), .B2(new_n863), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n887), .B1(new_n903), .B2(G148gat), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n886), .B1(new_n890), .B2(new_n904), .ZN(G1345gat));
  NOR2_X1   g704(.A1(new_n868), .A2(new_n593), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n906), .A2(KEYINPUT122), .ZN(new_n907));
  AOI21_X1  g706(.A(G155gat), .B1(new_n906), .B2(KEYINPUT122), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n593), .A2(new_n294), .ZN(new_n909));
  AOI22_X1  g708(.A1(new_n907), .A2(new_n908), .B1(new_n889), .B2(new_n909), .ZN(G1346gat));
  AOI21_X1  g709(.A(G162gat), .B1(new_n869), .B2(new_n623), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n706), .A2(new_n295), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n889), .B2(new_n912), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n656), .A2(new_n659), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n814), .A2(new_n815), .A3(new_n914), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n915), .A2(new_n247), .A3(new_n557), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n891), .A2(new_n821), .A3(new_n914), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(G169gat), .B1(new_n918), .B2(new_n685), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n916), .A2(new_n919), .ZN(G1348gat));
  OAI21_X1  g719(.A(G176gat), .B1(new_n915), .B2(new_n686), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n918), .A2(new_n248), .A3(new_n650), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1349gat));
  OR2_X1    g722(.A1(new_n915), .A2(new_n593), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n592), .A2(new_n225), .ZN(new_n925));
  AOI22_X1  g724(.A1(new_n924), .A2(G183gat), .B1(new_n918), .B2(new_n925), .ZN(new_n926));
  XOR2_X1   g725(.A(KEYINPUT123), .B(KEYINPUT60), .Z(new_n927));
  XNOR2_X1  g726(.A(new_n926), .B(new_n927), .ZN(G1350gat));
  INV_X1    g727(.A(new_n706), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n918), .A2(new_n226), .A3(new_n929), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n915), .A2(new_n625), .ZN(new_n931));
  XNOR2_X1  g730(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n931), .A2(G190gat), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n931), .B2(G190gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(G1351gat));
  NAND2_X1  g734(.A1(new_n900), .A2(KEYINPUT125), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n914), .A2(new_n667), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n892), .A2(new_n898), .A3(new_n939), .A4(new_n899), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n936), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(G197gat), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n941), .A2(new_n942), .A3(new_n557), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n813), .A2(new_n445), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n938), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(G197gat), .B1(new_n946), .B2(new_n685), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n943), .A2(new_n947), .ZN(G1352gat));
  OAI21_X1  g747(.A(G204gat), .B1(new_n941), .B2(new_n686), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n651), .A2(G204gat), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n944), .A2(new_n938), .A3(new_n950), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT62), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT126), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n949), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1353gat));
  NOR2_X1   g756(.A1(new_n937), .A2(new_n593), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n204), .B1(new_n900), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT63), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n946), .A2(new_n204), .A3(new_n592), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1354gat));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n941), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(new_n623), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n941), .A2(new_n963), .ZN(new_n966));
  OAI21_X1  g765(.A(G218gat), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n946), .A2(new_n205), .A3(new_n929), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(G1355gat));
endmodule


