

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738;

  INV_X1 U372 ( .A(n479), .ZN(n354) );
  BUF_X1 U373 ( .A(G116), .Z(n353) );
  XNOR2_X2 U374 ( .A(n352), .B(n373), .ZN(n432) );
  XNOR2_X2 U375 ( .A(n372), .B(n371), .ZN(n352) );
  XNOR2_X1 U376 ( .A(n480), .B(n354), .ZN(n357) );
  NAND2_X1 U377 ( .A1(n478), .A2(n477), .ZN(n480) );
  OR2_X1 U378 ( .A1(n599), .A2(G902), .ZN(n437) );
  XNOR2_X1 U379 ( .A(n398), .B(n368), .ZN(n727) );
  XNOR2_X1 U380 ( .A(n661), .B(KEYINPUT6), .ZN(n490) );
  INV_X1 U381 ( .A(G953), .ZN(n728) );
  NOR2_X1 U382 ( .A1(n574), .A2(n642), .ZN(n553) );
  XNOR2_X1 U383 ( .A(n553), .B(KEYINPUT40), .ZN(n737) );
  AND2_X4 U384 ( .A1(n593), .A2(n592), .ZN(n622) );
  BUF_X1 U385 ( .A(n661), .Z(n355) );
  INV_X1 U386 ( .A(n566), .ZN(n657) );
  INV_X1 U387 ( .A(n488), .ZN(n566) );
  NOR2_X1 U388 ( .A1(n630), .A2(n649), .ZN(n512) );
  XNOR2_X1 U389 ( .A(G125), .B(G146), .ZN(n376) );
  XNOR2_X2 U390 ( .A(G119), .B(G116), .ZN(n372) );
  NOR2_X1 U391 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U392 ( .A(n570), .B(n569), .ZN(n571) );
  NOR2_X1 U393 ( .A1(n643), .A2(n675), .ZN(n556) );
  XNOR2_X1 U394 ( .A(n403), .B(G469), .ZN(n537) );
  XNOR2_X1 U395 ( .A(n432), .B(n375), .ZN(n719) );
  INV_X1 U396 ( .A(n376), .ZN(n404) );
  BUF_X1 U397 ( .A(n554), .Z(n356) );
  XNOR2_X2 U398 ( .A(n528), .B(n527), .ZN(n694) );
  OR2_X1 U399 ( .A1(n624), .A2(G902), .ZN(n403) );
  XNOR2_X1 U400 ( .A(n378), .B(n379), .ZN(n361) );
  XNOR2_X1 U401 ( .A(n366), .B(n365), .ZN(n572) );
  INV_X1 U402 ( .A(KEYINPUT46), .ZN(n365) );
  NOR2_X1 U403 ( .A1(n737), .A2(n736), .ZN(n366) );
  XNOR2_X1 U404 ( .A(n434), .B(n433), .ZN(n599) );
  XNOR2_X1 U405 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U406 ( .A(n727), .B(G146), .ZN(n434) );
  AND2_X1 U407 ( .A1(n363), .A2(n551), .ZN(n552) );
  INV_X1 U408 ( .A(n672), .ZN(n551) );
  INV_X1 U409 ( .A(KEYINPUT28), .ZN(n535) );
  XNOR2_X1 U410 ( .A(G122), .B(G143), .ZN(n445) );
  XNOR2_X1 U411 ( .A(n401), .B(n398), .ZN(n358) );
  XNOR2_X1 U412 ( .A(n719), .B(n360), .ZN(n359) );
  XNOR2_X1 U413 ( .A(n542), .B(n541), .ZN(n670) );
  AND2_X1 U414 ( .A1(n549), .A2(n550), .ZN(n363) );
  INV_X1 U415 ( .A(KEYINPUT89), .ZN(n395) );
  XNOR2_X1 U416 ( .A(n469), .B(n468), .ZN(n472) );
  INV_X1 U417 ( .A(n591), .ZN(n592) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n607) );
  XNOR2_X1 U419 ( .A(n377), .B(n361), .ZN(n360) );
  INV_X1 U420 ( .A(n692), .ZN(n585) );
  NAND2_X1 U421 ( .A1(n362), .A2(n582), .ZN(n692) );
  XNOR2_X1 U422 ( .A(n573), .B(KEYINPUT48), .ZN(n362) );
  NAND2_X1 U423 ( .A1(n692), .A2(KEYINPUT77), .ZN(n587) );
  NAND2_X1 U424 ( .A1(n363), .A2(n558), .ZN(n641) );
  XNOR2_X2 U425 ( .A(n364), .B(G143), .ZN(n463) );
  XNOR2_X2 U426 ( .A(G128), .B(KEYINPUT81), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n441), .B(n440), .ZN(n681) );
  BUF_X1 U428 ( .A(n694), .Z(n714) );
  XOR2_X1 U429 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n367) );
  XOR2_X1 U430 ( .A(n397), .B(n396), .Z(n368) );
  INV_X1 U431 ( .A(KEYINPUT68), .ZN(n569) );
  NOR2_X2 U432 ( .A1(n526), .A2(n525), .ZN(n528) );
  XNOR2_X1 U433 ( .A(n580), .B(n540), .ZN(n672) );
  XNOR2_X1 U434 ( .A(n419), .B(KEYINPUT25), .ZN(n420) );
  XNOR2_X1 U435 ( .A(n404), .B(KEYINPUT10), .ZN(n405) );
  NOR2_X1 U436 ( .A1(n672), .A2(n671), .ZN(n676) );
  INV_X1 U437 ( .A(KEYINPUT34), .ZN(n443) );
  XNOR2_X1 U438 ( .A(n405), .B(G140), .ZN(n726) );
  NAND2_X1 U439 ( .A1(n562), .A2(n561), .ZN(n577) );
  XOR2_X1 U440 ( .A(n472), .B(n471), .Z(n594) );
  INV_X1 U441 ( .A(KEYINPUT63), .ZN(n603) );
  XNOR2_X1 U442 ( .A(G107), .B(G104), .ZN(n369) );
  XNOR2_X1 U443 ( .A(n369), .B(G110), .ZN(n720) );
  XNOR2_X1 U444 ( .A(KEYINPUT64), .B(G101), .ZN(n429) );
  XNOR2_X1 U445 ( .A(n429), .B(KEYINPUT72), .ZN(n370) );
  XNOR2_X1 U446 ( .A(n720), .B(n370), .ZN(n401) );
  XNOR2_X2 U447 ( .A(G113), .B(KEYINPUT70), .ZN(n371) );
  XNOR2_X1 U448 ( .A(KEYINPUT71), .B(KEYINPUT3), .ZN(n373) );
  XNOR2_X1 U449 ( .A(KEYINPUT16), .B(G122), .ZN(n375) );
  XNOR2_X2 U450 ( .A(n463), .B(KEYINPUT4), .ZN(n398) );
  XOR2_X1 U451 ( .A(KEYINPUT18), .B(KEYINPUT79), .Z(n378) );
  XNOR2_X1 U452 ( .A(n404), .B(KEYINPUT17), .ZN(n377) );
  NAND2_X1 U453 ( .A1(n728), .A2(G224), .ZN(n379) );
  XNOR2_X1 U454 ( .A(KEYINPUT86), .B(KEYINPUT15), .ZN(n380) );
  XNOR2_X1 U455 ( .A(n380), .B(G902), .ZN(n591) );
  NAND2_X1 U456 ( .A1(n607), .A2(n591), .ZN(n383) );
  INV_X1 U457 ( .A(G237), .ZN(n381) );
  NAND2_X1 U458 ( .A1(n474), .A2(n381), .ZN(n384) );
  NAND2_X1 U459 ( .A1(n384), .A2(G210), .ZN(n382) );
  XNOR2_X2 U460 ( .A(n383), .B(n382), .ZN(n539) );
  NAND2_X1 U461 ( .A1(n384), .A2(G214), .ZN(n385) );
  XNOR2_X1 U462 ( .A(n385), .B(KEYINPUT87), .ZN(n671) );
  NOR2_X2 U463 ( .A1(n539), .A2(n671), .ZN(n563) );
  INV_X1 U464 ( .A(KEYINPUT78), .ZN(n386) );
  XOR2_X1 U465 ( .A(n386), .B(KEYINPUT19), .Z(n387) );
  XNOR2_X1 U466 ( .A(n563), .B(n387), .ZN(n554) );
  NAND2_X1 U467 ( .A1(G237), .A2(G234), .ZN(n388) );
  XNOR2_X1 U468 ( .A(n388), .B(KEYINPUT14), .ZN(n391) );
  NAND2_X1 U469 ( .A1(G902), .A2(n391), .ZN(n389) );
  XOR2_X1 U470 ( .A(KEYINPUT88), .B(n389), .Z(n390) );
  NAND2_X1 U471 ( .A1(G953), .A2(n390), .ZN(n529) );
  NOR2_X1 U472 ( .A1(n529), .A2(G898), .ZN(n392) );
  NAND2_X1 U473 ( .A1(G952), .A2(n391), .ZN(n688) );
  NOR2_X1 U474 ( .A1(n688), .A2(G953), .ZN(n531) );
  NOR2_X1 U475 ( .A1(n392), .A2(n531), .ZN(n393) );
  OR2_X2 U476 ( .A1(n554), .A2(n393), .ZN(n394) );
  XNOR2_X2 U477 ( .A(n394), .B(KEYINPUT0), .ZN(n509) );
  XNOR2_X1 U478 ( .A(n509), .B(n395), .ZN(n505) );
  INV_X1 U479 ( .A(n505), .ZN(n442) );
  XNOR2_X1 U480 ( .A(G137), .B(G134), .ZN(n397) );
  XNOR2_X1 U481 ( .A(G131), .B(KEYINPUT67), .ZN(n396) );
  NAND2_X1 U482 ( .A1(n728), .A2(G227), .ZN(n399) );
  XNOR2_X1 U483 ( .A(n399), .B(G140), .ZN(n400) );
  XNOR2_X1 U484 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U485 ( .A(n434), .B(n402), .ZN(n624) );
  XNOR2_X1 U486 ( .A(n537), .B(KEYINPUT1), .ZN(n488) );
  XOR2_X1 U487 ( .A(G137), .B(G119), .Z(n407) );
  XNOR2_X1 U488 ( .A(G128), .B(G110), .ZN(n406) );
  XNOR2_X1 U489 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U490 ( .A(n726), .B(n408), .ZN(n416) );
  XNOR2_X1 U491 ( .A(KEYINPUT91), .B(KEYINPUT24), .ZN(n409) );
  XNOR2_X1 U492 ( .A(n409), .B(KEYINPUT23), .ZN(n410) );
  XOR2_X1 U493 ( .A(KEYINPUT90), .B(n410), .Z(n414) );
  XOR2_X1 U494 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n412) );
  NAND2_X1 U495 ( .A1(G234), .A2(n728), .ZN(n411) );
  XNOR2_X1 U496 ( .A(n412), .B(n411), .ZN(n470) );
  NAND2_X1 U497 ( .A1(G221), .A2(n470), .ZN(n413) );
  XNOR2_X1 U498 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U499 ( .A(n416), .B(n415), .ZN(n707) );
  NOR2_X1 U500 ( .A1(n707), .A2(G902), .ZN(n421) );
  NAND2_X1 U501 ( .A1(n591), .A2(G234), .ZN(n418) );
  XNOR2_X1 U502 ( .A(KEYINPUT92), .B(KEYINPUT20), .ZN(n417) );
  XNOR2_X1 U503 ( .A(n418), .B(n417), .ZN(n422) );
  NAND2_X1 U504 ( .A1(n422), .A2(G217), .ZN(n419) );
  XNOR2_X2 U505 ( .A(n421), .B(n420), .ZN(n532) );
  INV_X1 U506 ( .A(n532), .ZN(n517) );
  NAND2_X1 U507 ( .A1(G221), .A2(n422), .ZN(n424) );
  INV_X1 U508 ( .A(KEYINPUT21), .ZN(n423) );
  XNOR2_X1 U509 ( .A(n424), .B(n423), .ZN(n659) );
  AND2_X1 U510 ( .A1(n532), .A2(n659), .ZN(n656) );
  NAND2_X1 U511 ( .A1(n488), .A2(n656), .ZN(n426) );
  INV_X1 U512 ( .A(KEYINPUT106), .ZN(n425) );
  XNOR2_X1 U513 ( .A(n426), .B(n425), .ZN(n438) );
  NOR2_X1 U514 ( .A1(G953), .A2(G237), .ZN(n451) );
  NAND2_X1 U515 ( .A1(n451), .A2(G210), .ZN(n428) );
  XNOR2_X1 U516 ( .A(KEYINPUT76), .B(KEYINPUT5), .ZN(n427) );
  XNOR2_X1 U517 ( .A(n428), .B(n427), .ZN(n430) );
  XNOR2_X1 U518 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U519 ( .A(n432), .B(n431), .ZN(n433) );
  INV_X1 U520 ( .A(KEYINPUT93), .ZN(n435) );
  XNOR2_X1 U521 ( .A(n435), .B(G472), .ZN(n436) );
  XNOR2_X2 U522 ( .A(n437), .B(n436), .ZN(n661) );
  INV_X1 U523 ( .A(n490), .ZN(n562) );
  NAND2_X1 U524 ( .A1(n438), .A2(n562), .ZN(n441) );
  XNOR2_X1 U525 ( .A(KEYINPUT107), .B(KEYINPUT33), .ZN(n439) );
  XNOR2_X1 U526 ( .A(n439), .B(KEYINPUT73), .ZN(n440) );
  NAND2_X1 U527 ( .A1(n442), .A2(n681), .ZN(n444) );
  XNOR2_X1 U528 ( .A(n444), .B(n443), .ZN(n478) );
  XOR2_X1 U529 ( .A(G104), .B(KEYINPUT97), .Z(n446) );
  XNOR2_X1 U530 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U531 ( .A(KEYINPUT96), .B(KEYINPUT98), .Z(n448) );
  XNOR2_X1 U532 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n447) );
  XNOR2_X1 U533 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U534 ( .A(n450), .B(n449), .ZN(n455) );
  XOR2_X1 U535 ( .A(G131), .B(G113), .Z(n453) );
  NAND2_X1 U536 ( .A1(n451), .A2(G214), .ZN(n452) );
  XNOR2_X1 U537 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U538 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U539 ( .A(n726), .B(n456), .ZN(n617) );
  NOR2_X1 U540 ( .A1(G902), .A2(n617), .ZN(n457) );
  XOR2_X1 U541 ( .A(G475), .B(n457), .Z(n459) );
  INV_X1 U542 ( .A(KEYINPUT13), .ZN(n458) );
  XNOR2_X1 U543 ( .A(n459), .B(n458), .ZN(n514) );
  XNOR2_X1 U544 ( .A(G478), .B(KEYINPUT103), .ZN(n476) );
  INV_X1 U545 ( .A(G902), .ZN(n474) );
  XNOR2_X1 U546 ( .A(KEYINPUT7), .B(KEYINPUT99), .ZN(n460) );
  XNOR2_X1 U547 ( .A(n367), .B(n460), .ZN(n462) );
  XOR2_X1 U548 ( .A(n353), .B(G107), .Z(n461) );
  XNOR2_X1 U549 ( .A(n462), .B(n461), .ZN(n469) );
  INV_X1 U550 ( .A(n463), .ZN(n467) );
  XOR2_X1 U551 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n465) );
  XNOR2_X1 U552 ( .A(G134), .B(G122), .ZN(n464) );
  XNOR2_X1 U553 ( .A(n465), .B(n464), .ZN(n466) );
  NAND2_X1 U554 ( .A1(G217), .A2(n470), .ZN(n471) );
  INV_X1 U555 ( .A(n594), .ZN(n473) );
  NAND2_X1 U556 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U557 ( .A(n476), .B(n475), .ZN(n513) );
  INV_X1 U558 ( .A(n513), .ZN(n484) );
  NAND2_X1 U559 ( .A1(n514), .A2(n484), .ZN(n557) );
  INV_X1 U560 ( .A(n557), .ZN(n477) );
  XNOR2_X1 U561 ( .A(KEYINPUT80), .B(KEYINPUT35), .ZN(n479) );
  XNOR2_X2 U562 ( .A(n480), .B(n479), .ZN(n615) );
  NOR2_X1 U563 ( .A1(KEYINPUT44), .A2(KEYINPUT65), .ZN(n481) );
  NAND2_X1 U564 ( .A1(n357), .A2(n481), .ZN(n483) );
  NAND2_X1 U565 ( .A1(n615), .A2(KEYINPUT65), .ZN(n482) );
  NAND2_X1 U566 ( .A1(n483), .A2(n482), .ZN(n497) );
  NOR2_X1 U567 ( .A1(n514), .A2(n484), .ZN(n673) );
  NAND2_X1 U568 ( .A1(n673), .A2(n659), .ZN(n485) );
  OR2_X1 U569 ( .A1(n509), .A2(n485), .ZN(n487) );
  XNOR2_X1 U570 ( .A(KEYINPUT74), .B(KEYINPUT22), .ZN(n486) );
  XNOR2_X1 U571 ( .A(n487), .B(n486), .ZN(n520) );
  NOR2_X1 U572 ( .A1(n566), .A2(n532), .ZN(n489) );
  XOR2_X1 U573 ( .A(KEYINPUT105), .B(n489), .Z(n491) );
  NAND2_X1 U574 ( .A1(n491), .A2(n490), .ZN(n492) );
  NOR2_X1 U575 ( .A1(n520), .A2(n492), .ZN(n493) );
  XNOR2_X1 U576 ( .A(n493), .B(KEYINPUT32), .ZN(n735) );
  OR2_X1 U577 ( .A1(n532), .A2(n355), .ZN(n494) );
  OR2_X1 U578 ( .A1(n657), .A2(n494), .ZN(n495) );
  NOR2_X1 U579 ( .A1(n520), .A2(n495), .ZN(n634) );
  NOR2_X1 U580 ( .A1(n735), .A2(n634), .ZN(n496) );
  NAND2_X1 U581 ( .A1(n497), .A2(n496), .ZN(n504) );
  INV_X1 U582 ( .A(KEYINPUT85), .ZN(n498) );
  NAND2_X1 U583 ( .A1(n615), .A2(n498), .ZN(n501) );
  OR2_X1 U584 ( .A1(n634), .A2(KEYINPUT65), .ZN(n499) );
  NOR2_X1 U585 ( .A1(n735), .A2(n499), .ZN(n500) );
  NAND2_X1 U586 ( .A1(n501), .A2(n500), .ZN(n502) );
  NAND2_X1 U587 ( .A1(n502), .A2(KEYINPUT44), .ZN(n503) );
  NAND2_X1 U588 ( .A1(n504), .A2(n503), .ZN(n526) );
  AND2_X1 U589 ( .A1(n656), .A2(n537), .ZN(n546) );
  INV_X1 U590 ( .A(n355), .ZN(n506) );
  NAND2_X1 U591 ( .A1(n546), .A2(n506), .ZN(n507) );
  NOR2_X1 U592 ( .A1(n505), .A2(n507), .ZN(n630) );
  AND2_X1 U593 ( .A1(n657), .A2(n656), .ZN(n508) );
  NAND2_X1 U594 ( .A1(n508), .A2(n355), .ZN(n665) );
  NOR2_X1 U595 ( .A1(n665), .A2(n509), .ZN(n511) );
  XOR2_X1 U596 ( .A(KEYINPUT94), .B(KEYINPUT31), .Z(n510) );
  XNOR2_X1 U597 ( .A(n511), .B(n510), .ZN(n649) );
  XOR2_X1 U598 ( .A(KEYINPUT95), .B(n512), .Z(n516) );
  AND2_X1 U599 ( .A1(n514), .A2(n513), .ZN(n645) );
  OR2_X1 U600 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X2 U601 ( .A(n515), .B(KEYINPUT104), .ZN(n635) );
  INV_X1 U602 ( .A(n635), .ZN(n648) );
  NOR2_X1 U603 ( .A1(n645), .A2(n648), .ZN(n675) );
  NOR2_X1 U604 ( .A1(n516), .A2(n675), .ZN(n521) );
  NOR2_X1 U605 ( .A1(n657), .A2(n517), .ZN(n518) );
  NAND2_X1 U606 ( .A1(n518), .A2(n490), .ZN(n519) );
  NOR2_X1 U607 ( .A1(n520), .A2(n519), .ZN(n605) );
  NOR2_X1 U608 ( .A1(n521), .A2(n605), .ZN(n524) );
  NAND2_X1 U609 ( .A1(n615), .A2(KEYINPUT44), .ZN(n522) );
  NAND2_X1 U610 ( .A1(n522), .A2(KEYINPUT85), .ZN(n523) );
  NAND2_X1 U611 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U612 ( .A(KEYINPUT84), .B(KEYINPUT45), .Z(n527) );
  NOR2_X1 U613 ( .A1(G900), .A2(n529), .ZN(n530) );
  NOR2_X1 U614 ( .A1(n531), .A2(n530), .ZN(n544) );
  NOR2_X1 U615 ( .A1(n544), .A2(n532), .ZN(n533) );
  NAND2_X1 U616 ( .A1(n533), .A2(n659), .ZN(n534) );
  XNOR2_X1 U617 ( .A(n534), .B(KEYINPUT69), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n560), .A2(n355), .ZN(n536) );
  XNOR2_X1 U619 ( .A(n536), .B(n535), .ZN(n538) );
  NAND2_X1 U620 ( .A1(n538), .A2(n537), .ZN(n555) );
  BUF_X1 U621 ( .A(n539), .Z(n580) );
  XNOR2_X1 U622 ( .A(KEYINPUT38), .B(KEYINPUT75), .ZN(n540) );
  NAND2_X1 U623 ( .A1(n676), .A2(n673), .ZN(n542) );
  XOR2_X1 U624 ( .A(KEYINPUT41), .B(KEYINPUT108), .Z(n541) );
  NOR2_X1 U625 ( .A1(n555), .A2(n670), .ZN(n543) );
  XNOR2_X1 U626 ( .A(n543), .B(KEYINPUT42), .ZN(n736) );
  INV_X1 U627 ( .A(n544), .ZN(n545) );
  AND2_X1 U628 ( .A1(n546), .A2(n545), .ZN(n550) );
  INV_X1 U629 ( .A(n671), .ZN(n547) );
  AND2_X1 U630 ( .A1(n661), .A2(n547), .ZN(n548) );
  XNOR2_X1 U631 ( .A(n548), .B(KEYINPUT30), .ZN(n549) );
  XNOR2_X1 U632 ( .A(n552), .B(KEYINPUT39), .ZN(n574) );
  INV_X1 U633 ( .A(n645), .ZN(n642) );
  OR2_X2 U634 ( .A1(n555), .A2(n356), .ZN(n643) );
  XNOR2_X1 U635 ( .A(n556), .B(KEYINPUT47), .ZN(n559) );
  NOR2_X1 U636 ( .A1(n580), .A2(n557), .ZN(n558) );
  AND2_X1 U637 ( .A1(n559), .A2(n641), .ZN(n568) );
  AND2_X1 U638 ( .A1(n560), .A2(n645), .ZN(n561) );
  XNOR2_X1 U639 ( .A(n577), .B(KEYINPUT109), .ZN(n564) );
  NAND2_X1 U640 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U641 ( .A(n565), .B(KEYINPUT36), .ZN(n567) );
  OR2_X2 U642 ( .A1(n567), .A2(n566), .ZN(n652) );
  AND2_X2 U643 ( .A1(n568), .A2(n652), .ZN(n570) );
  NOR2_X1 U644 ( .A1(n635), .A2(n574), .ZN(n575) );
  XNOR2_X1 U645 ( .A(n575), .B(KEYINPUT110), .ZN(n738) );
  OR2_X1 U646 ( .A1(n657), .A2(n671), .ZN(n576) );
  NOR2_X1 U647 ( .A1(n577), .A2(n576), .ZN(n579) );
  INV_X1 U648 ( .A(KEYINPUT43), .ZN(n578) );
  XNOR2_X1 U649 ( .A(n579), .B(n578), .ZN(n581) );
  AND2_X1 U650 ( .A1(n581), .A2(n580), .ZN(n606) );
  NOR2_X1 U651 ( .A1(n738), .A2(n606), .ZN(n582) );
  INV_X1 U652 ( .A(n692), .ZN(n697) );
  NAND2_X1 U653 ( .A1(n694), .A2(n697), .ZN(n583) );
  NAND2_X1 U654 ( .A1(n583), .A2(KEYINPUT2), .ZN(n590) );
  NOR2_X1 U655 ( .A1(KEYINPUT2), .A2(KEYINPUT77), .ZN(n584) );
  NAND2_X1 U656 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U658 ( .A1(n588), .A2(n694), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U660 ( .A1(n622), .A2(G478), .ZN(n595) );
  XNOR2_X1 U661 ( .A(n595), .B(n594), .ZN(n597) );
  INV_X1 U662 ( .A(G952), .ZN(n596) );
  AND2_X1 U663 ( .A1(n596), .A2(G953), .ZN(n709) );
  NOR2_X2 U664 ( .A1(n597), .A2(n709), .ZN(n598) );
  XNOR2_X1 U665 ( .A(n598), .B(KEYINPUT122), .ZN(G63) );
  NAND2_X1 U666 ( .A1(n622), .A2(G472), .ZN(n601) );
  XNOR2_X1 U667 ( .A(n599), .B(KEYINPUT62), .ZN(n600) );
  XNOR2_X1 U668 ( .A(n601), .B(n600), .ZN(n602) );
  NOR2_X2 U669 ( .A1(n602), .A2(n709), .ZN(n604) );
  XNOR2_X1 U670 ( .A(n604), .B(n603), .ZN(G57) );
  XOR2_X1 U671 ( .A(G101), .B(n605), .Z(G3) );
  XOR2_X1 U672 ( .A(G140), .B(n606), .Z(G42) );
  NAND2_X1 U673 ( .A1(n622), .A2(G210), .ZN(n611) );
  XNOR2_X1 U674 ( .A(KEYINPUT82), .B(KEYINPUT54), .ZN(n608) );
  XNOR2_X1 U675 ( .A(n608), .B(KEYINPUT55), .ZN(n609) );
  XNOR2_X1 U676 ( .A(n607), .B(n609), .ZN(n610) );
  XNOR2_X1 U677 ( .A(n611), .B(n610), .ZN(n612) );
  NOR2_X2 U678 ( .A1(n612), .A2(n709), .ZN(n614) );
  XOR2_X1 U679 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n613) );
  XNOR2_X1 U680 ( .A(n614), .B(n613), .ZN(G51) );
  XNOR2_X1 U681 ( .A(G122), .B(KEYINPUT127), .ZN(n616) );
  XNOR2_X1 U682 ( .A(n615), .B(n616), .ZN(G24) );
  NAND2_X1 U683 ( .A1(n622), .A2(G475), .ZN(n619) );
  XOR2_X1 U684 ( .A(KEYINPUT59), .B(n617), .Z(n618) );
  XNOR2_X1 U685 ( .A(n619), .B(n618), .ZN(n620) );
  NOR2_X2 U686 ( .A1(n620), .A2(n709), .ZN(n621) );
  XNOR2_X1 U687 ( .A(n621), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U688 ( .A1(n622), .A2(G469), .ZN(n626) );
  XOR2_X1 U689 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n623) );
  XNOR2_X1 U690 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U691 ( .A(n626), .B(n625), .ZN(n627) );
  NOR2_X1 U692 ( .A1(n627), .A2(n709), .ZN(G54) );
  XOR2_X1 U693 ( .A(G104), .B(KEYINPUT111), .Z(n629) );
  NAND2_X1 U694 ( .A1(n630), .A2(n645), .ZN(n628) );
  XNOR2_X1 U695 ( .A(n629), .B(n628), .ZN(G6) );
  XOR2_X1 U696 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n632) );
  NAND2_X1 U697 ( .A1(n630), .A2(n648), .ZN(n631) );
  XNOR2_X1 U698 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U699 ( .A(G107), .B(n633), .ZN(G9) );
  XOR2_X1 U700 ( .A(G110), .B(n634), .Z(G12) );
  NOR2_X1 U701 ( .A1(n643), .A2(n635), .ZN(n640) );
  XOR2_X1 U702 ( .A(KEYINPUT29), .B(KEYINPUT114), .Z(n637) );
  XNOR2_X1 U703 ( .A(G128), .B(KEYINPUT113), .ZN(n636) );
  XNOR2_X1 U704 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U705 ( .A(KEYINPUT112), .B(n638), .ZN(n639) );
  XNOR2_X1 U706 ( .A(n640), .B(n639), .ZN(G30) );
  XNOR2_X1 U707 ( .A(G143), .B(n641), .ZN(G45) );
  NOR2_X1 U708 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U709 ( .A(G146), .B(n644), .Z(G48) );
  XOR2_X1 U710 ( .A(G113), .B(KEYINPUT115), .Z(n647) );
  NAND2_X1 U711 ( .A1(n645), .A2(n649), .ZN(n646) );
  XNOR2_X1 U712 ( .A(n647), .B(n646), .ZN(G15) );
  NAND2_X1 U713 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U714 ( .A(n650), .B(KEYINPUT116), .ZN(n651) );
  XNOR2_X1 U715 ( .A(n353), .B(n651), .ZN(G18) );
  XOR2_X1 U716 ( .A(G125), .B(n652), .Z(n653) );
  XNOR2_X1 U717 ( .A(n653), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 U718 ( .A(n681), .ZN(n654) );
  NOR2_X1 U719 ( .A1(n654), .A2(n670), .ZN(n655) );
  NOR2_X1 U720 ( .A1(n655), .A2(G953), .ZN(n691) );
  XOR2_X1 U721 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n686) );
  NOR2_X1 U722 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U723 ( .A(KEYINPUT50), .B(n658), .Z(n664) );
  NOR2_X1 U724 ( .A1(n659), .A2(n532), .ZN(n660) );
  XOR2_X1 U725 ( .A(KEYINPUT49), .B(n660), .Z(n662) );
  NOR2_X1 U726 ( .A1(n662), .A2(n355), .ZN(n663) );
  NAND2_X1 U727 ( .A1(n664), .A2(n663), .ZN(n666) );
  NAND2_X1 U728 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U729 ( .A(n667), .B(KEYINPUT117), .Z(n668) );
  XNOR2_X1 U730 ( .A(KEYINPUT51), .B(n668), .ZN(n669) );
  NOR2_X1 U731 ( .A1(n670), .A2(n669), .ZN(n683) );
  NAND2_X1 U732 ( .A1(n672), .A2(n671), .ZN(n674) );
  NAND2_X1 U733 ( .A1(n674), .A2(n673), .ZN(n679) );
  INV_X1 U734 ( .A(n675), .ZN(n677) );
  NAND2_X1 U735 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U736 ( .A1(n679), .A2(n678), .ZN(n680) );
  AND2_X1 U737 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U738 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U739 ( .A(n684), .B(KEYINPUT52), .ZN(n685) );
  XNOR2_X1 U740 ( .A(n686), .B(n685), .ZN(n687) );
  NOR2_X1 U741 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U742 ( .A(KEYINPUT120), .B(n689), .Z(n690) );
  NAND2_X1 U743 ( .A1(n691), .A2(n690), .ZN(n704) );
  XNOR2_X1 U744 ( .A(KEYINPUT2), .B(KEYINPUT83), .ZN(n693) );
  NAND2_X1 U745 ( .A1(n693), .A2(n692), .ZN(n700) );
  NAND2_X1 U746 ( .A1(n714), .A2(KEYINPUT2), .ZN(n696) );
  INV_X1 U747 ( .A(KEYINPUT83), .ZN(n695) );
  NAND2_X1 U748 ( .A1(n696), .A2(n695), .ZN(n698) );
  NAND2_X1 U749 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U750 ( .A1(n700), .A2(n699), .ZN(n702) );
  NOR2_X1 U751 ( .A1(n714), .A2(KEYINPUT2), .ZN(n701) );
  NOR2_X1 U752 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U753 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U754 ( .A(KEYINPUT53), .B(n705), .ZN(G75) );
  NAND2_X1 U755 ( .A1(n622), .A2(G217), .ZN(n706) );
  XNOR2_X1 U756 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U757 ( .A1(n709), .A2(n708), .ZN(G66) );
  XOR2_X1 U758 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n711) );
  NAND2_X1 U759 ( .A1(G224), .A2(G953), .ZN(n710) );
  XNOR2_X1 U760 ( .A(n711), .B(n710), .ZN(n712) );
  NAND2_X1 U761 ( .A1(G898), .A2(n712), .ZN(n713) );
  XNOR2_X1 U762 ( .A(n713), .B(KEYINPUT124), .ZN(n717) );
  NAND2_X1 U763 ( .A1(n714), .A2(n728), .ZN(n715) );
  XOR2_X1 U764 ( .A(KEYINPUT125), .B(n715), .Z(n716) );
  NAND2_X1 U765 ( .A1(n717), .A2(n716), .ZN(n725) );
  XOR2_X1 U766 ( .A(G101), .B(KEYINPUT126), .Z(n718) );
  XNOR2_X1 U767 ( .A(n719), .B(n718), .ZN(n721) );
  XNOR2_X1 U768 ( .A(n721), .B(n720), .ZN(n723) );
  NOR2_X1 U769 ( .A1(n728), .A2(G898), .ZN(n722) );
  NOR2_X1 U770 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U771 ( .A(n725), .B(n724), .ZN(G69) );
  XNOR2_X1 U772 ( .A(n727), .B(n726), .ZN(n730) );
  XNOR2_X1 U773 ( .A(n697), .B(n730), .ZN(n729) );
  NAND2_X1 U774 ( .A1(n729), .A2(n728), .ZN(n734) );
  XOR2_X1 U775 ( .A(G227), .B(n730), .Z(n731) );
  NAND2_X1 U776 ( .A1(n731), .A2(G900), .ZN(n732) );
  NAND2_X1 U777 ( .A1(n732), .A2(G953), .ZN(n733) );
  NAND2_X1 U778 ( .A1(n734), .A2(n733), .ZN(G72) );
  XOR2_X1 U779 ( .A(G119), .B(n735), .Z(G21) );
  XOR2_X1 U780 ( .A(n736), .B(G137), .Z(G39) );
  XOR2_X1 U781 ( .A(G131), .B(n737), .Z(G33) );
  XOR2_X1 U782 ( .A(G134), .B(n738), .Z(G36) );
endmodule

