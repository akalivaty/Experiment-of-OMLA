//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n203), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT64), .B(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G58), .A2(G232), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n201), .ZN(new_n244));
  XOR2_X1   g0044(.A(KEYINPUT65), .B(G50), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n242), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G41), .ZN(new_n249));
  OAI211_X1 g0049(.A(G1), .B(G13), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT72), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n248), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G1698), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n251), .B1(new_n256), .B2(new_n231), .ZN(new_n257));
  AND2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(KEYINPUT72), .A3(G232), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1698), .B1(new_n253), .B2(new_n254), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n265), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n250), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT67), .A2(G41), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT67), .A2(G41), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G45), .ZN(new_n271));
  AOI21_X1  g0071(.A(G1), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n250), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n276), .B1(new_n220), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(KEYINPUT13), .B1(new_n267), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NOR3_X1   g0081(.A1(new_n267), .A2(KEYINPUT13), .A3(new_n279), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G169), .ZN(new_n284));
  OAI21_X1  g0084(.A(KEYINPUT14), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(G179), .ZN(new_n286));
  INV_X1    g0086(.A(new_n282), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n280), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT14), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(new_n289), .A3(G169), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n285), .A2(new_n286), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n215), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT68), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n293), .B(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n248), .A2(G20), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n296), .A2(G77), .B1(new_n297), .B2(G50), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(new_n207), .B2(new_n218), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT11), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT69), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT69), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n304), .A2(new_n206), .A3(G13), .A4(G20), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n293), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n207), .A2(G1), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G68), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n301), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  XOR2_X1   g0112(.A(KEYINPUT73), .B(KEYINPUT12), .Z(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(new_n306), .B2(new_n218), .ZN(new_n314));
  XOR2_X1   g0114(.A(new_n314), .B(KEYINPUT74), .Z(new_n315));
  NOR3_X1   g0115(.A1(new_n306), .A2(KEYINPUT12), .A3(G68), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n291), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G190), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n318), .B1(new_n288), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G200), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n283), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n306), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n295), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n329), .A2(G50), .A3(new_n310), .ZN(new_n330));
  OAI21_X1  g0130(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n331));
  INV_X1    g0131(.A(G150), .ZN(new_n332));
  INV_X1    g0132(.A(new_n297), .ZN(new_n333));
  INV_X1    g0133(.A(new_n296), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT8), .B(G58), .ZN(new_n335));
  OAI221_X1 g0135(.A(new_n331), .B1(new_n332), .B2(new_n333), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G50), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n336), .A2(new_n295), .B1(new_n337), .B2(new_n328), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n330), .A2(new_n338), .ZN(new_n339));
  XOR2_X1   g0139(.A(new_n339), .B(KEYINPUT9), .Z(new_n340));
  INV_X1    g0140(.A(G226), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n276), .B1(new_n341), .B2(new_n278), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n262), .A2(G223), .B1(G77), .B2(new_n260), .ZN(new_n343));
  INV_X1    g0143(.A(G222), .ZN(new_n344));
  INV_X1    g0144(.A(new_n265), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n342), .B1(new_n346), .B2(new_n273), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G190), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n323), .B2(new_n347), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n340), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n348), .B(KEYINPUT71), .C1(new_n323), .C2(new_n347), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT10), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n265), .A2(G232), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT70), .ZN(new_n356));
  INV_X1    g0156(.A(G107), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n256), .A2(new_n220), .B1(new_n357), .B2(new_n255), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(new_n250), .ZN(new_n360));
  INV_X1    g0160(.A(G244), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n276), .B1(new_n361), .B2(new_n278), .ZN(new_n362));
  OAI21_X1  g0162(.A(G200), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n362), .ZN(new_n364));
  OAI211_X1 g0164(.A(G190), .B(new_n364), .C1(new_n359), .C2(new_n250), .ZN(new_n365));
  INV_X1    g0165(.A(new_n335), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(new_n297), .B1(G20), .B2(G77), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT15), .B(G87), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n367), .B1(new_n334), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G77), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n369), .A2(new_n293), .B1(new_n370), .B2(new_n328), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n308), .A2(new_n370), .A3(new_n309), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n363), .A2(new_n365), .A3(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n284), .B1(new_n360), .B2(new_n362), .ZN(new_n377));
  INV_X1    g0177(.A(G179), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n378), .B(new_n364), .C1(new_n359), .C2(new_n250), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(new_n374), .A3(new_n379), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n352), .B(new_n351), .C1(new_n340), .C2(new_n349), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n347), .A2(new_n378), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n383), .B(new_n339), .C1(G169), .C2(new_n347), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n354), .A2(new_n381), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n335), .A2(new_n309), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n329), .A2(new_n386), .B1(new_n328), .B2(new_n335), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n253), .A2(new_n207), .A3(new_n254), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n253), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n254), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(KEYINPUT77), .A3(new_n391), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n391), .A2(KEYINPUT77), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n218), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT75), .ZN(new_n395));
  INV_X1    g0195(.A(G159), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n333), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(G58), .A2(G68), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n218), .B2(G58), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n395), .B(new_n398), .C1(new_n400), .C2(new_n207), .ZN(new_n401));
  AND2_X1   g0201(.A1(KEYINPUT64), .A2(G68), .ZN(new_n402));
  NOR2_X1   g0202(.A1(KEYINPUT64), .A2(G68), .ZN(new_n403));
  OAI21_X1  g0203(.A(G58), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n207), .B1(new_n404), .B2(new_n203), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT75), .B1(new_n405), .B2(new_n397), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n394), .A2(new_n401), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT16), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n293), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n390), .A2(new_n391), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G68), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT16), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n406), .A2(new_n401), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT76), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n406), .A2(new_n401), .A3(KEYINPUT76), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n413), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n387), .B1(new_n410), .B2(new_n418), .ZN(new_n419));
  MUX2_X1   g0219(.A(G223), .B(G226), .S(G1698), .Z(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(new_n255), .B1(G33), .B2(G87), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n276), .B1(new_n231), .B2(new_n278), .C1(new_n250), .C2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(new_n378), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(G169), .B2(new_n422), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n419), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n422), .A2(new_n323), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(G190), .B2(new_n422), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n387), .B(new_n429), .C1(new_n410), .C2(new_n418), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n387), .ZN(new_n433));
  INV_X1    g0233(.A(new_n413), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n406), .A2(new_n401), .A3(KEYINPUT76), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT76), .B1(new_n406), .B2(new_n401), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n307), .B1(new_n407), .B2(new_n408), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n433), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT18), .B1(new_n439), .B2(new_n424), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(KEYINPUT17), .A3(new_n429), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n427), .A2(new_n432), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n327), .A2(new_n385), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n392), .A2(G107), .A3(new_n393), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT79), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n333), .A2(new_n370), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  XNOR2_X1  g0248(.A(G97), .B(G107), .ZN(new_n449));
  NOR2_X1   g0249(.A1(KEYINPUT78), .A2(KEYINPUT6), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G97), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n450), .B1(KEYINPUT6), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n452), .B1(new_n449), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n448), .B1(new_n455), .B2(new_n207), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT79), .A4(G107), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n446), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n293), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n328), .A2(G97), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n293), .B(KEYINPUT68), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n206), .A2(G33), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(new_n306), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n461), .B1(new_n464), .B2(G97), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(G250), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G283), .ZN(new_n468));
  OAI211_X1 g0268(.A(G244), .B(new_n261), .C1(new_n258), .C2(new_n259), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT4), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n467), .B(new_n468), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT4), .B1(new_n265), .B2(G244), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n273), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT5), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n206), .B(G45), .C1(new_n474), .C2(G41), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n474), .B1(new_n268), .B2(new_n269), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n273), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g0278(.A(KEYINPUT67), .B(G41), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n475), .B1(new_n479), .B2(new_n474), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n478), .A2(G257), .B1(new_n480), .B2(new_n275), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G200), .ZN(new_n483));
  INV_X1    g0283(.A(new_n482), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G190), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n460), .A2(new_n466), .A3(new_n483), .A4(new_n485), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n473), .A2(new_n481), .A3(new_n378), .ZN(new_n487));
  AOI21_X1  g0287(.A(G169), .B1(new_n473), .B2(new_n481), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n456), .B1(new_n445), .B2(new_n444), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n307), .B1(new_n490), .B2(new_n458), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n489), .B1(new_n491), .B2(new_n465), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT82), .ZN(new_n494));
  INV_X1    g0294(.A(new_n368), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n306), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n462), .A2(G87), .A3(new_n306), .A4(new_n463), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT19), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n334), .B2(new_n453), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n255), .A2(new_n207), .A3(G68), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n207), .ZN(new_n504));
  OR2_X1    g0304(.A1(new_n504), .A2(KEYINPUT80), .ZN(new_n505));
  INV_X1    g0305(.A(G87), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(new_n453), .A3(new_n357), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT81), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT81), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n509), .A2(new_n506), .A3(new_n453), .A4(new_n357), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n508), .A2(new_n510), .B1(KEYINPUT80), .B2(new_n504), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n502), .B1(new_n505), .B2(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n497), .B(new_n498), .C1(new_n512), .C2(new_n307), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n206), .A2(new_n274), .A3(G45), .ZN(new_n515));
  INV_X1    g0315(.A(G250), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n271), .B2(G1), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n250), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(G238), .B(new_n261), .C1(new_n258), .C2(new_n259), .ZN(new_n520));
  OAI211_X1 g0320(.A(G244), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n521));
  INV_X1    g0321(.A(G116), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n520), .B(new_n521), .C1(new_n248), .C2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n519), .B1(new_n523), .B2(new_n273), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n524), .A2(new_n323), .ZN(new_n525));
  AOI211_X1 g0325(.A(new_n321), .B(new_n519), .C1(new_n523), .C2(new_n273), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n524), .A2(G169), .ZN(new_n528));
  AOI211_X1 g0328(.A(G179), .B(new_n519), .C1(new_n523), .C2(new_n273), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n462), .A2(new_n306), .A3(new_n495), .A4(new_n463), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n531), .B(new_n497), .C1(new_n512), .C2(new_n307), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n514), .A2(new_n527), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n493), .A2(new_n494), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n493), .A2(new_n533), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT82), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n328), .A2(new_n522), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n306), .A2(new_n307), .A3(G116), .A4(new_n463), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n468), .B(new_n207), .C1(G33), .C2(new_n453), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n522), .A2(G20), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n293), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT20), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n541), .A2(new_n542), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n537), .B(new_n538), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(G264), .B(G1698), .C1(new_n258), .C2(new_n259), .ZN(new_n546));
  OAI211_X1 g0346(.A(G257), .B(new_n261), .C1(new_n258), .C2(new_n259), .ZN(new_n547));
  INV_X1    g0347(.A(G303), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n546), .B(new_n547), .C1(new_n548), .C2(new_n255), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n273), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n478), .A2(G270), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n480), .A2(new_n275), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n545), .A2(new_n553), .A3(G169), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT21), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n553), .A2(new_n378), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n545), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n545), .A2(new_n553), .A3(KEYINPUT21), .A4(G169), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n255), .A2(G257), .A3(G1698), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G294), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n562), .B(new_n563), .C1(new_n345), .C2(new_n516), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n273), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n478), .A2(G264), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n552), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n284), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n565), .A2(new_n378), .A3(new_n552), .A4(new_n566), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OR3_X1    g0370(.A1(new_n306), .A2(KEYINPUT25), .A3(G107), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT25), .B1(new_n306), .B2(G107), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(new_n464), .C2(new_n357), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT85), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n329), .A2(G107), .A3(new_n463), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n576), .A2(KEYINPUT85), .A3(new_n571), .A4(new_n572), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT23), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(new_n357), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n357), .A3(G20), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n581), .A2(KEYINPUT84), .B1(new_n582), .B2(G20), .ZN(new_n583));
  AOI211_X1 g0383(.A(new_n580), .B(new_n583), .C1(KEYINPUT84), .C2(new_n581), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n255), .A2(new_n207), .A3(G87), .ZN(new_n585));
  XNOR2_X1  g0385(.A(new_n585), .B(KEYINPUT22), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT24), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n584), .A2(new_n586), .A3(KEYINPUT24), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(new_n293), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n570), .B1(new_n578), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n565), .A2(new_n566), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(G190), .A3(new_n552), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n567), .A2(G200), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n578), .A2(new_n591), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n553), .A2(G200), .ZN(new_n598));
  INV_X1    g0398(.A(new_n545), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n598), .B(new_n599), .C1(new_n321), .C2(new_n553), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT83), .ZN(new_n601));
  OR2_X1    g0401(.A1(new_n553), .A2(new_n321), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT83), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n602), .A2(new_n603), .A3(new_n599), .A4(new_n598), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  AND4_X1   g0405(.A1(new_n561), .A2(new_n593), .A3(new_n597), .A4(new_n605), .ZN(new_n606));
  AND4_X1   g0406(.A1(new_n443), .A2(new_n534), .A3(new_n536), .A4(new_n606), .ZN(G372));
  INV_X1    g0407(.A(new_n384), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n326), .A2(new_n432), .A3(new_n441), .ZN(new_n609));
  INV_X1    g0409(.A(new_n380), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n291), .B2(new_n319), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n440), .B(new_n427), .C1(new_n609), .C2(new_n611), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n354), .A2(new_n382), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n608), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT86), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n560), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n556), .A2(new_n558), .A3(KEYINPUT86), .A4(new_n559), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n592), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n597), .A2(new_n486), .A3(new_n492), .A4(new_n533), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n530), .A2(new_n532), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT87), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n532), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n524), .A2(new_n378), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(G169), .B2(new_n524), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n524), .A2(G190), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n323), .B2(new_n524), .ZN(new_n628));
  OAI22_X1  g0428(.A1(new_n624), .A2(new_n626), .B1(new_n628), .B2(new_n513), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT26), .B1(new_n492), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n460), .A2(new_n466), .ZN(new_n631));
  XOR2_X1   g0431(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n632));
  NAND4_X1  g0432(.A1(new_n533), .A2(new_n631), .A3(new_n489), .A4(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n623), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  OR2_X1    g0434(.A1(new_n620), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n443), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n614), .A2(new_n636), .ZN(G369));
  NAND3_X1  g0437(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G213), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n641), .B(KEYINPUT89), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G343), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n592), .A2(new_n643), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n578), .A2(new_n591), .A3(new_n595), .A4(new_n596), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n643), .B1(new_n578), .B2(new_n591), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n593), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n560), .A2(new_n643), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n644), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT90), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI211_X1 g0452(.A(KEYINPUT90), .B(new_n644), .C1(new_n648), .C2(new_n649), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n605), .B(new_n561), .C1(new_n599), .C2(new_n643), .ZN(new_n655));
  INV_X1    g0455(.A(new_n643), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n616), .A2(new_n545), .A3(new_n617), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(G330), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n647), .A2(new_n644), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n654), .A2(new_n662), .ZN(G399));
  INV_X1    g0463(.A(new_n210), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(new_n479), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n508), .A2(new_n522), .A3(new_n510), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n665), .A2(new_n206), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n667), .B1(new_n214), .B2(new_n665), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n668), .B(KEYINPUT28), .Z(new_n669));
  INV_X1    g0469(.A(G330), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n536), .A2(new_n606), .A3(new_n534), .A4(new_n643), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n557), .A2(new_n594), .A3(new_n484), .A4(new_n524), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT30), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n524), .A2(G179), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n567), .A2(new_n675), .A3(new_n482), .A4(new_n553), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n672), .A2(new_n673), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n678), .A2(KEYINPUT31), .A3(new_n656), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT31), .B1(new_n678), .B2(new_n656), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n670), .B1(new_n671), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n643), .B1(new_n620), .B2(new_n634), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT91), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT29), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT91), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n686), .B(new_n643), .C1(new_n620), .C2(new_n634), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n632), .B1(new_n492), .B2(new_n629), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n533), .A2(new_n631), .A3(KEYINPUT26), .A4(new_n489), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT92), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n492), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(KEYINPUT92), .A3(KEYINPUT26), .A4(new_n533), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n692), .A2(KEYINPUT93), .A3(new_n623), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n593), .A2(new_n561), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(new_n493), .A3(new_n533), .A4(new_n597), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n621), .B(KEYINPUT87), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT26), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n492), .A2(new_n629), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n699), .B1(new_n701), .B2(KEYINPUT92), .ZN(new_n702));
  AOI21_X1  g0502(.A(KEYINPUT93), .B1(new_n702), .B2(new_n692), .ZN(new_n703));
  OAI211_X1 g0503(.A(KEYINPUT29), .B(new_n643), .C1(new_n698), .C2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n682), .B1(new_n688), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n669), .B1(new_n705), .B2(G1), .ZN(G364));
  NAND2_X1  g0506(.A1(new_n207), .A2(G13), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n206), .B1(new_n708), .B2(G45), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n665), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n658), .B2(G330), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(G330), .B2(new_n658), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n664), .A2(new_n260), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G355), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(G116), .B2(new_n210), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n246), .A2(new_n271), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n664), .A2(new_n255), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n271), .B2(new_n214), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n716), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G13), .A2(G33), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n215), .B1(G20), .B2(new_n284), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n711), .B1(new_n721), .B2(new_n727), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n321), .A2(G179), .A3(G200), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n207), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n207), .A2(new_n378), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G190), .A2(G200), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n731), .A2(G294), .B1(new_n735), .B2(G311), .ZN(new_n736));
  INV_X1    g0536(.A(G326), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n732), .A2(G200), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n321), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n736), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT94), .Z(new_n742));
  NOR2_X1   g0542(.A1(new_n207), .A2(G179), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n733), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G329), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n732), .A2(G190), .A3(new_n323), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n255), .B1(new_n748), .B2(G322), .ZN(new_n749));
  INV_X1    g0549(.A(G283), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n743), .A2(new_n321), .A3(G200), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n743), .A2(G190), .A3(G200), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n750), .A2(new_n751), .B1(new_n752), .B2(new_n548), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n738), .A2(G190), .ZN(new_n754));
  INV_X1    g0554(.A(G317), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n755), .A2(KEYINPUT33), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(KEYINPUT33), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n753), .B1(new_n754), .B2(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n742), .A2(new_n746), .A3(new_n749), .A4(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT32), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n744), .A2(new_n396), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n740), .A2(new_n337), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(G68), .B2(new_n754), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n255), .B1(new_n734), .B2(new_n370), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(G58), .B2(new_n748), .ZN(new_n766));
  INV_X1    g0566(.A(new_n752), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n731), .A2(G97), .B1(new_n767), .B2(G87), .ZN(new_n768));
  INV_X1    g0568(.A(new_n751), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n761), .A2(new_n762), .B1(new_n769), .B2(G107), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n764), .A2(new_n766), .A3(new_n768), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n760), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n728), .B1(new_n772), .B2(new_n725), .ZN(new_n773));
  INV_X1    g0573(.A(new_n724), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n773), .B1(new_n658), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n713), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(G396));
  INV_X1    g0577(.A(G132), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n255), .B1(new_n744), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(G68), .B2(new_n769), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n731), .A2(G58), .B1(new_n767), .B2(G50), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n748), .A2(G143), .B1(new_n735), .B2(G159), .ZN(new_n782));
  INV_X1    g0582(.A(G137), .ZN(new_n783));
  INV_X1    g0583(.A(new_n754), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n782), .B1(new_n740), .B2(new_n783), .C1(new_n332), .C2(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT96), .B(KEYINPUT34), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n780), .B(new_n781), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n754), .A2(KEYINPUT95), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n754), .A2(KEYINPUT95), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n750), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n731), .A2(G97), .B1(new_n767), .B2(G107), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n739), .A2(G303), .B1(new_n769), .B2(G87), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n255), .B1(new_n748), .B2(G294), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G116), .A2(new_n735), .B1(new_n745), .B2(G311), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n793), .A2(new_n794), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n787), .A2(new_n788), .B1(new_n792), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n725), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n725), .A2(new_n722), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n799), .B(new_n711), .C1(G77), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n380), .A2(new_n656), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n376), .B1(new_n375), .B2(new_n643), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(new_n804), .B2(new_n380), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n802), .B1(new_n806), .B2(new_n722), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n684), .A2(new_n687), .A3(new_n806), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n805), .B(new_n643), .C1(new_n620), .C2(new_n634), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n682), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n711), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n808), .A2(new_n682), .A3(new_n809), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n807), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(G384));
  NAND2_X1  g0614(.A1(new_n416), .A2(new_n417), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n462), .B1(new_n815), .B2(new_n434), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n412), .B1(new_n435), .B2(new_n436), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n408), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n433), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n642), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n442), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT97), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n442), .A2(KEYINPUT97), .A3(new_n821), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n430), .B1(new_n819), .B2(new_n424), .ZN(new_n827));
  OAI21_X1  g0627(.A(KEYINPUT37), .B1(new_n827), .B2(new_n821), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n419), .A2(new_n425), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n419), .A2(new_n642), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT37), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n829), .A2(new_n830), .A3(new_n831), .A4(new_n430), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(KEYINPUT38), .B1(new_n826), .B2(new_n833), .ZN(new_n834));
  AND3_X1   g0634(.A1(new_n442), .A2(KEYINPUT97), .A3(new_n821), .ZN(new_n835));
  AOI21_X1  g0635(.A(KEYINPUT97), .B1(new_n442), .B2(new_n821), .ZN(new_n836));
  OAI211_X1 g0636(.A(KEYINPUT38), .B(new_n833), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(KEYINPUT98), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT38), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT98), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n842), .A2(new_n843), .A3(new_n837), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n671), .A2(new_n681), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n319), .A2(new_n656), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n320), .A2(new_n326), .A3(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n319), .B(new_n656), .C1(new_n291), .C2(new_n325), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n846), .A2(new_n850), .A3(new_n805), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT40), .B1(new_n845), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n430), .B1(new_n439), .B2(new_n424), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n439), .A2(new_n820), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT37), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n856), .A2(new_n832), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n442), .A2(new_n855), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n841), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n837), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT40), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n851), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n853), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n443), .A2(new_n846), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n865), .A2(new_n866), .A3(new_n670), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n842), .A2(KEYINPUT39), .A3(new_n837), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT39), .B1(new_n837), .B2(new_n859), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n291), .A2(new_n319), .A3(new_n643), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n803), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n809), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n845), .A2(new_n850), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n427), .A2(new_n440), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n820), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n873), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n688), .A2(new_n704), .A3(new_n443), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n614), .ZN(new_n881));
  XOR2_X1   g0681(.A(new_n879), .B(new_n881), .Z(new_n882));
  OAI22_X1  g0682(.A1(new_n867), .A2(new_n882), .B1(new_n206), .B2(new_n708), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n882), .B2(new_n867), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT35), .ZN(new_n885));
  OAI211_X1 g0685(.A(G116), .B(new_n216), .C1(new_n455), .C2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(new_n885), .B2(new_n455), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT36), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n214), .A2(G77), .A3(new_n404), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n337), .A2(G68), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n206), .B(G13), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  OR3_X1    g0691(.A1(new_n884), .A2(new_n888), .A3(new_n891), .ZN(G367));
  OAI221_X1 g0692(.A(new_n726), .B1(new_n210), .B2(new_n368), .C1(new_n719), .C2(new_n237), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n893), .A2(new_n711), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n514), .A2(new_n643), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n699), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n629), .B2(new_n895), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n739), .A2(G311), .B1(new_n769), .B2(G97), .ZN(new_n898));
  INV_X1    g0698(.A(G294), .ZN(new_n899));
  OAI221_X1 g0699(.A(new_n898), .B1(new_n357), .B2(new_n730), .C1(new_n791), .C2(new_n899), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n767), .A2(KEYINPUT46), .A3(G116), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT46), .B1(new_n767), .B2(G116), .ZN(new_n902));
  AOI22_X1  g0702(.A1(G283), .A2(new_n735), .B1(new_n745), .B2(G317), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n903), .B(new_n260), .C1(new_n548), .C2(new_n747), .ZN(new_n904));
  NOR4_X1   g0704(.A1(new_n900), .A2(new_n901), .A3(new_n902), .A4(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT106), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n791), .A2(new_n396), .ZN(new_n907));
  AOI22_X1  g0707(.A1(G68), .A2(new_n731), .B1(new_n739), .B2(G143), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n260), .B1(new_n735), .B2(G50), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n748), .A2(G150), .B1(new_n745), .B2(G137), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n767), .A2(G58), .B1(new_n769), .B2(G77), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n908), .A2(new_n909), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n906), .B1(new_n907), .B2(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n913), .B(KEYINPUT47), .Z(new_n914));
  INV_X1    g0714(.A(new_n725), .ZN(new_n915));
  OAI221_X1 g0715(.A(new_n894), .B1(new_n774), .B2(new_n897), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n631), .A2(new_n656), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n493), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n693), .A2(new_n656), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT45), .B1(new_n654), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT45), .ZN(new_n922));
  INV_X1    g0722(.A(new_n920), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n922), .B(new_n923), .C1(new_n652), .C2(new_n653), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT44), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n654), .B2(new_n920), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n927), .A2(KEYINPUT102), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n652), .A2(KEYINPUT44), .A3(new_n653), .A4(new_n923), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n927), .A2(KEYINPUT102), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n925), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT103), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n931), .A2(new_n932), .A3(new_n662), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n660), .A2(new_n649), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT104), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n660), .A2(new_n649), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n660), .A2(new_n935), .A3(new_n649), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n659), .A2(KEYINPUT105), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n705), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n933), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n930), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n921), .A2(new_n924), .B1(new_n927), .B2(KEYINPUT102), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n661), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n925), .A2(new_n928), .A3(new_n662), .A4(new_n930), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n950), .A2(new_n951), .B1(new_n931), .B2(new_n932), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n705), .B1(new_n947), .B2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n665), .B(KEYINPUT41), .Z(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n710), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n934), .A2(new_n920), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(KEYINPUT101), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT42), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n957), .A2(KEYINPUT101), .ZN(new_n961));
  OR3_X1    g0761(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n920), .B(KEYINPUT100), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n492), .B1(new_n963), .B2(new_n593), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n643), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n960), .B1(new_n959), .B2(new_n961), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n962), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n897), .A2(KEYINPUT99), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n897), .A2(KEYINPUT99), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(KEYINPUT43), .B2(new_n897), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n967), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n967), .B2(new_n971), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n662), .A2(new_n963), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n975), .B(new_n976), .Z(new_n977));
  OAI21_X1  g0777(.A(new_n916), .B1(new_n956), .B2(new_n977), .ZN(G387));
  AOI22_X1  g0778(.A1(new_n714), .A2(new_n666), .B1(new_n357), .B2(new_n664), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n234), .A2(G45), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT107), .ZN(new_n981));
  XOR2_X1   g0781(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n366), .B2(new_n337), .ZN(new_n983));
  AOI211_X1 g0783(.A(G45), .B(new_n983), .C1(G68), .C2(G77), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n666), .A2(KEYINPUT108), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n366), .A2(new_n982), .A3(new_n337), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n666), .A2(KEYINPUT108), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n718), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n979), .B1(new_n981), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n711), .B1(new_n991), .B2(new_n727), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n747), .A2(new_n755), .B1(new_n734), .B2(new_n548), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G322), .B2(new_n739), .ZN(new_n994));
  INV_X1    g0794(.A(G311), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n994), .B1(new_n791), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT48), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n997), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n730), .A2(new_n750), .B1(new_n752), .B2(new_n899), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT110), .Z(new_n1001));
  NAND3_X1  g0801(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT49), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n260), .B1(new_n744), .B2(new_n737), .C1(new_n522), .C2(new_n751), .ZN(new_n1006));
  OR3_X1    g0806(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n734), .A2(new_n202), .B1(new_n744), .B2(new_n332), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n260), .B(new_n1008), .C1(G50), .C2(new_n748), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n767), .A2(G77), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n495), .A2(new_n731), .B1(new_n754), .B2(new_n366), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n739), .A2(G159), .B1(new_n769), .B2(G97), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n915), .B1(new_n1007), .B2(new_n1013), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n992), .B(new_n1014), .C1(new_n660), .C2(new_n724), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n944), .B2(new_n710), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n944), .A2(new_n705), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n945), .A2(new_n665), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(G393));
  AND2_X1   g0819(.A1(new_n950), .A2(new_n951), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n710), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n242), .A2(new_n719), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n726), .B1(new_n453), .B2(new_n210), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n711), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n255), .B1(new_n734), .B2(new_n335), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n731), .A2(G77), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n506), .B2(new_n751), .C1(new_n219), .C2(new_n752), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1025), .B(new_n1027), .C1(G143), .C2(new_n745), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n740), .A2(new_n332), .B1(new_n396), .B2(new_n747), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT51), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1028), .B(new_n1030), .C1(new_n337), .C2(new_n791), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT111), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n740), .A2(new_n755), .B1(new_n995), .B2(new_n747), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT52), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n791), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(G303), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n260), .B1(new_n734), .B2(new_n899), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G322), .B2(new_n745), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n357), .A2(new_n751), .B1(new_n752), .B2(new_n750), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G116), .B2(new_n731), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1035), .A2(new_n1037), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1033), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1024), .B1(new_n1044), .B2(new_n725), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n963), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1045), .B1(new_n1046), .B2(new_n774), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n665), .B1(new_n1020), .B2(new_n946), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n947), .A2(new_n952), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1021), .B(new_n1047), .C1(new_n1048), .C2(new_n1049), .ZN(G390));
  AOI21_X1  g0850(.A(new_n872), .B1(new_n875), .B2(new_n850), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n868), .B2(new_n869), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n860), .A2(new_n871), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n848), .A2(new_n849), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n804), .A2(new_n380), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n643), .B(new_n1056), .C1(new_n698), .C2(new_n703), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1055), .B1(new_n1057), .B2(new_n874), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n682), .A2(new_n805), .A3(new_n850), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1053), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n846), .A2(G330), .A3(new_n805), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1062), .A2(new_n1055), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n842), .A2(KEYINPUT39), .A3(new_n837), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT39), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n860), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1051), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1063), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1061), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n682), .A2(new_n443), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n880), .A2(new_n614), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n850), .B1(new_n682), .B2(new_n805), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n875), .B1(new_n1063), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1062), .A2(new_n1055), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1075), .A2(new_n874), .A3(new_n1057), .A4(new_n1060), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1072), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1070), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1061), .A2(new_n1069), .A3(new_n1077), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(new_n665), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1061), .A2(new_n1069), .A3(new_n710), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n711), .B1(new_n366), .B2(new_n801), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(KEYINPUT54), .B(G143), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n731), .A2(G159), .B1(new_n735), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n791), .B2(new_n783), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT112), .Z(new_n1088));
  NAND2_X1  g0888(.A1(new_n767), .A2(G150), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT53), .ZN(new_n1090));
  INV_X1    g0890(.A(G125), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n255), .B1(new_n744), .B2(new_n1091), .C1(new_n747), .C2(new_n778), .ZN(new_n1092));
  INV_X1    g0892(.A(G128), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n740), .A2(new_n1093), .B1(new_n751), .B2(new_n337), .ZN(new_n1094));
  OR3_X1    g0894(.A1(new_n1090), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n751), .A2(new_n202), .B1(new_n744), .B2(new_n899), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT113), .Z(new_n1097));
  OAI221_X1 g0897(.A(new_n260), .B1(new_n734), .B2(new_n453), .C1(new_n522), .C2(new_n747), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1026), .B1(new_n506), .B2(new_n752), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(G283), .C2(new_n739), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n357), .B2(new_n791), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n1088), .A2(new_n1095), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1083), .B1(new_n1102), .B2(new_n725), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n870), .B2(new_n723), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1081), .A2(new_n1082), .A3(new_n1104), .ZN(G378));
  INV_X1    g0905(.A(KEYINPUT117), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n670), .B1(new_n862), .B2(new_n860), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1106), .B1(new_n853), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n851), .B1(new_n839), .B2(new_n844), .ZN(new_n1110));
  OAI211_X1 g0910(.A(KEYINPUT117), .B(new_n1107), .C1(new_n1110), .C2(KEYINPUT40), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n613), .A2(new_n384), .ZN(new_n1114));
  XOR2_X1   g0914(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n1115));
  OR2_X1    g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n339), .A2(new_n642), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1117), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1113), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1121), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(new_n1112), .A3(new_n1119), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1109), .A2(new_n1111), .A3(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n853), .A2(new_n1108), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1128), .A2(KEYINPUT117), .A3(new_n1125), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n879), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1072), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1080), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT118), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1080), .A2(KEYINPUT118), .A3(new_n1132), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n879), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1127), .A2(new_n1138), .A3(new_n1129), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1131), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT57), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1131), .A2(new_n1137), .A3(KEYINPUT57), .A4(new_n1139), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n665), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1131), .A2(new_n710), .A3(new_n1139), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n800), .A2(new_n337), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n711), .A2(new_n1146), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n784), .A2(new_n778), .B1(new_n740), .B2(new_n1091), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n748), .A2(G128), .B1(new_n735), .B2(G137), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n752), .B2(new_n1084), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1148), .B(new_n1150), .C1(G150), .C2(new_n731), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n769), .A2(G159), .ZN(new_n1155));
  AOI211_X1 g0955(.A(G33), .B(G41), .C1(new_n745), .C2(G124), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n740), .A2(new_n522), .B1(new_n751), .B2(new_n201), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G97), .B2(new_n754), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n255), .B(new_n479), .C1(new_n745), .C2(G283), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n748), .A2(G107), .B1(new_n735), .B2(new_n495), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n731), .A2(G68), .B1(new_n767), .B2(G77), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT114), .B(KEYINPUT58), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n337), .B1(G33), .B2(G41), .C1(new_n255), .C2(new_n479), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1157), .A2(new_n1165), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1147), .B1(new_n1168), .B2(new_n725), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n1126), .B2(new_n723), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1145), .A2(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1144), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(G375));
  NAND2_X1  g0973(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n710), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n711), .B1(G68), .B2(new_n801), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n740), .A2(new_n899), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n260), .B1(new_n734), .B2(new_n357), .C1(new_n750), .C2(new_n747), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n730), .A2(new_n368), .B1(new_n751), .B2(new_n370), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n522), .B2(new_n791), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n752), .A2(new_n453), .B1(new_n744), .B2(new_n548), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT119), .Z(new_n1183));
  OAI22_X1  g0983(.A1(new_n734), .A2(new_n332), .B1(new_n744), .B2(new_n1093), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n260), .B(new_n1184), .C1(G137), .C2(new_n748), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n739), .A2(G132), .B1(new_n769), .B2(G58), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n731), .A2(G50), .B1(new_n767), .B2(G159), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n791), .A2(new_n1084), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n1181), .A2(new_n1183), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1176), .B1(new_n1190), .B2(new_n725), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n850), .B2(new_n723), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1175), .A2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1077), .A2(new_n954), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1174), .A2(new_n1132), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1193), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(G381));
  NOR2_X1   g0998(.A1(G393), .A2(G396), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(KEYINPUT120), .B1(new_n1200), .B2(G384), .ZN(new_n1201));
  INV_X1    g1001(.A(G390), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1201), .A2(new_n1202), .A3(new_n1197), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1200), .A2(KEYINPUT120), .A3(G384), .ZN(new_n1204));
  NOR4_X1   g1004(.A1(new_n1203), .A2(G387), .A3(G378), .A4(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n1172), .ZN(G407));
  INV_X1    g1006(.A(G378), .ZN(new_n1207));
  INV_X1    g1007(.A(G213), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(G343), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1172), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT121), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1211), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1012(.A(KEYINPUT61), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1144), .A2(G378), .A3(new_n1171), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1145), .B(new_n1170), .C1(new_n1140), .C2(new_n954), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n1207), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1209), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1078), .A2(new_n1195), .A3(KEYINPUT60), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1218), .A2(new_n665), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1195), .B1(KEYINPUT60), .B2(new_n1078), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1193), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n813), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(G384), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1209), .A2(G2897), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1226), .B(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1213), .B1(new_n1217), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(KEYINPUT124), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT124), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1232), .B(new_n1213), .C1(new_n1217), .C2(new_n1229), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1226), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1217), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT62), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT62), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1217), .A2(new_n1237), .A3(new_n1234), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1231), .A2(new_n1233), .A3(new_n1236), .A4(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(G393), .B(new_n776), .ZN(new_n1240));
  OAI211_X1 g1040(.A(G390), .B(new_n916), .C1(new_n956), .C2(new_n977), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT122), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1240), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(G387), .A2(new_n1202), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1241), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1245), .A2(new_n1243), .A3(new_n1241), .A4(new_n1240), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1239), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1230), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1249), .B1(new_n1235), .B2(new_n1252), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1217), .A2(new_n1234), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT123), .B1(new_n1254), .B2(KEYINPUT63), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT123), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1235), .A2(new_n1256), .A3(new_n1252), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1251), .B(new_n1253), .C1(new_n1255), .C2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1250), .A2(new_n1258), .ZN(G405));
  INV_X1    g1059(.A(KEYINPUT126), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1247), .A2(new_n1260), .A3(new_n1248), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT127), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1261), .B(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1214), .A2(KEYINPUT125), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(G375), .A2(new_n1207), .A3(new_n1234), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1226), .B1(new_n1172), .B2(G378), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1265), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1249), .A2(KEYINPUT126), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1266), .A2(new_n1265), .A3(new_n1267), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1263), .A2(new_n1269), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1261), .B(KEYINPUT127), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1270), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1273), .B1(new_n1274), .B2(new_n1268), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1275), .ZN(G402));
endmodule


