

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(n689), .A2(n691), .ZN(n582) );
  INV_X1 U549 ( .A(n634), .ZN(n654) );
  XNOR2_X2 U550 ( .A(KEYINPUT17), .B(KEYINPUT69), .ZN(n513) );
  NOR2_X2 U551 ( .A1(G2104), .A2(G2105), .ZN(n512) );
  OR2_X1 U552 ( .A1(n622), .A2(n621), .ZN(n625) );
  XNOR2_X1 U553 ( .A(KEYINPUT67), .B(KEYINPUT23), .ZN(n522) );
  AND2_X2 U554 ( .A1(n517), .A2(G2104), .ZN(n868) );
  NOR2_X1 U555 ( .A1(n529), .A2(n528), .ZN(G160) );
  INV_X1 U556 ( .A(KEYINPUT28), .ZN(n629) );
  NOR2_X1 U557 ( .A1(n647), .A2(n646), .ZN(n648) );
  INV_X1 U558 ( .A(n983), .ZN(n673) );
  AND2_X1 U559 ( .A1(n660), .A2(n659), .ZN(n649) );
  NAND2_X1 U560 ( .A1(n654), .A2(G8), .ZN(n588) );
  INV_X1 U561 ( .A(KEYINPUT66), .ZN(n580) );
  NOR2_X1 U562 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U563 ( .A1(G651), .A2(n541), .ZN(n790) );
  XNOR2_X1 U564 ( .A(n523), .B(n522), .ZN(n525) );
  NOR2_X1 U565 ( .A1(n521), .A2(n520), .ZN(G164) );
  XNOR2_X2 U566 ( .A(n513), .B(n512), .ZN(n869) );
  NAND2_X1 U567 ( .A1(n869), .A2(G138), .ZN(n515) );
  INV_X1 U568 ( .A(G2105), .ZN(n517) );
  NAND2_X1 U569 ( .A1(G102), .A2(n868), .ZN(n514) );
  NAND2_X1 U570 ( .A1(n515), .A2(n514), .ZN(n521) );
  NAND2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  XOR2_X1 U572 ( .A(KEYINPUT68), .B(n516), .Z(n698) );
  NAND2_X1 U573 ( .A1(G114), .A2(n698), .ZN(n519) );
  NOR2_X2 U574 ( .A1(G2104), .A2(n517), .ZN(n873) );
  NAND2_X1 U575 ( .A1(n873), .A2(G126), .ZN(n518) );
  NAND2_X1 U576 ( .A1(n519), .A2(n518), .ZN(n520) );
  NAND2_X1 U577 ( .A1(G101), .A2(n868), .ZN(n523) );
  NAND2_X1 U578 ( .A1(G113), .A2(n698), .ZN(n524) );
  NAND2_X1 U579 ( .A1(n525), .A2(n524), .ZN(n529) );
  NAND2_X1 U580 ( .A1(G137), .A2(n869), .ZN(n527) );
  NAND2_X1 U581 ( .A1(G125), .A2(n873), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U583 ( .A(KEYINPUT2), .B(KEYINPUT86), .Z(n531) );
  XOR2_X1 U584 ( .A(G543), .B(KEYINPUT0), .Z(n541) );
  INV_X1 U585 ( .A(G651), .ZN(n536) );
  NOR2_X1 U586 ( .A1(n541), .A2(n536), .ZN(n783) );
  NAND2_X1 U587 ( .A1(G73), .A2(n783), .ZN(n530) );
  XNOR2_X1 U588 ( .A(n531), .B(n530), .ZN(n535) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n782) );
  NAND2_X1 U590 ( .A1(G86), .A2(n782), .ZN(n533) );
  NAND2_X1 U591 ( .A1(G48), .A2(n790), .ZN(n532) );
  NAND2_X1 U592 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U593 ( .A1(n535), .A2(n534), .ZN(n540) );
  NOR2_X1 U594 ( .A1(G543), .A2(n536), .ZN(n537) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n537), .Z(n538) );
  XNOR2_X1 U596 ( .A(KEYINPUT70), .B(n538), .ZN(n787) );
  NAND2_X1 U597 ( .A1(G61), .A2(n787), .ZN(n539) );
  NAND2_X1 U598 ( .A1(n540), .A2(n539), .ZN(G305) );
  NAND2_X1 U599 ( .A1(G49), .A2(n790), .ZN(n543) );
  NAND2_X1 U600 ( .A1(G87), .A2(n541), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U602 ( .A1(n787), .A2(n544), .ZN(n547) );
  NAND2_X1 U603 ( .A1(G74), .A2(G651), .ZN(n545) );
  XOR2_X1 U604 ( .A(KEYINPUT85), .B(n545), .Z(n546) );
  NAND2_X1 U605 ( .A1(n547), .A2(n546), .ZN(G288) );
  NAND2_X1 U606 ( .A1(G90), .A2(n782), .ZN(n549) );
  NAND2_X1 U607 ( .A1(G77), .A2(n783), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U609 ( .A(n550), .B(KEYINPUT9), .ZN(n552) );
  NAND2_X1 U610 ( .A1(G52), .A2(n790), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n555) );
  NAND2_X1 U612 ( .A1(G64), .A2(n787), .ZN(n553) );
  XNOR2_X1 U613 ( .A(KEYINPUT71), .B(n553), .ZN(n554) );
  NOR2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U615 ( .A(KEYINPUT72), .B(n556), .ZN(G171) );
  NAND2_X1 U616 ( .A1(G51), .A2(n790), .ZN(n558) );
  NAND2_X1 U617 ( .A1(G63), .A2(n787), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U619 ( .A(KEYINPUT6), .B(n559), .ZN(n566) );
  NAND2_X1 U620 ( .A1(n782), .A2(G89), .ZN(n560) );
  XNOR2_X1 U621 ( .A(n560), .B(KEYINPUT4), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G76), .A2(n783), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U624 ( .A(KEYINPUT78), .B(n563), .Z(n564) );
  XNOR2_X1 U625 ( .A(KEYINPUT5), .B(n564), .ZN(n565) );
  NOR2_X1 U626 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U627 ( .A(KEYINPUT7), .B(n567), .Z(G168) );
  NAND2_X1 U628 ( .A1(G88), .A2(n782), .ZN(n569) );
  NAND2_X1 U629 ( .A1(G75), .A2(n783), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U631 ( .A1(G50), .A2(n790), .ZN(n571) );
  NAND2_X1 U632 ( .A1(G62), .A2(n787), .ZN(n570) );
  NAND2_X1 U633 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U634 ( .A1(n573), .A2(n572), .ZN(G166) );
  XNOR2_X1 U635 ( .A(KEYINPUT91), .B(G166), .ZN(G303) );
  XOR2_X1 U636 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U637 ( .A1(G85), .A2(n782), .ZN(n575) );
  NAND2_X1 U638 ( .A1(G72), .A2(n783), .ZN(n574) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U640 ( .A1(G47), .A2(n790), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G60), .A2(n787), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  OR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(G290) );
  NOR2_X1 U644 ( .A1(G164), .A2(G1384), .ZN(n581) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n689) );
  NAND2_X1 U646 ( .A1(G160), .A2(G40), .ZN(n691) );
  XNOR2_X2 U647 ( .A(KEYINPUT64), .B(n582), .ZN(n634) );
  NOR2_X1 U648 ( .A1(G1981), .A2(G305), .ZN(n583) );
  XOR2_X1 U649 ( .A(n583), .B(KEYINPUT24), .Z(n584) );
  NOR2_X1 U650 ( .A1(n588), .A2(n584), .ZN(n681) );
  XOR2_X1 U651 ( .A(G1981), .B(G305), .Z(n990) );
  NOR2_X1 U652 ( .A1(G288), .A2(G1976), .ZN(n585) );
  XNOR2_X1 U653 ( .A(n585), .B(KEYINPUT100), .ZN(n670) );
  INV_X1 U654 ( .A(n670), .ZN(n984) );
  NOR2_X1 U655 ( .A1(n588), .A2(n984), .ZN(n586) );
  NAND2_X1 U656 ( .A1(KEYINPUT33), .A2(n586), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n990), .A2(n587), .ZN(n679) );
  OR2_X1 U658 ( .A1(n588), .A2(G1966), .ZN(n642) );
  INV_X1 U659 ( .A(n642), .ZN(n650) );
  NAND2_X1 U660 ( .A1(G53), .A2(n790), .ZN(n590) );
  NAND2_X1 U661 ( .A1(G65), .A2(n787), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U663 ( .A1(G91), .A2(n782), .ZN(n592) );
  NAND2_X1 U664 ( .A1(G78), .A2(n783), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n798) );
  NAND2_X1 U667 ( .A1(G2072), .A2(n634), .ZN(n595) );
  XNOR2_X1 U668 ( .A(n595), .B(KEYINPUT27), .ZN(n597) );
  INV_X1 U669 ( .A(G1956), .ZN(n932) );
  NOR2_X1 U670 ( .A1(n634), .A2(n932), .ZN(n596) );
  NOR2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n628) );
  NAND2_X1 U672 ( .A1(n798), .A2(n628), .ZN(n627) );
  NAND2_X1 U673 ( .A1(n782), .A2(G81), .ZN(n598) );
  XNOR2_X1 U674 ( .A(n598), .B(KEYINPUT12), .ZN(n600) );
  NAND2_X1 U675 ( .A1(G68), .A2(n783), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U677 ( .A(n601), .B(KEYINPUT13), .ZN(n603) );
  NAND2_X1 U678 ( .A1(G43), .A2(n790), .ZN(n602) );
  NAND2_X1 U679 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n787), .A2(G56), .ZN(n604) );
  XOR2_X1 U681 ( .A(KEYINPUT14), .B(n604), .Z(n605) );
  NOR2_X1 U682 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U683 ( .A(KEYINPUT77), .B(n607), .ZN(n993) );
  NAND2_X1 U684 ( .A1(n634), .A2(G1996), .ZN(n608) );
  XNOR2_X1 U685 ( .A(n608), .B(KEYINPUT26), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n654), .A2(G1341), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U688 ( .A1(n993), .A2(n611), .ZN(n622) );
  NAND2_X1 U689 ( .A1(G54), .A2(n790), .ZN(n613) );
  NAND2_X1 U690 ( .A1(G66), .A2(n787), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U692 ( .A1(G92), .A2(n782), .ZN(n615) );
  NAND2_X1 U693 ( .A1(G79), .A2(n783), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U696 ( .A(n618), .B(KEYINPUT15), .ZN(n994) );
  NAND2_X1 U697 ( .A1(G2067), .A2(n634), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n654), .A2(G1348), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n623) );
  NOR2_X1 U700 ( .A1(n994), .A2(n623), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n994), .A2(n623), .ZN(n624) );
  NAND2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n632) );
  NOR2_X1 U704 ( .A1(n798), .A2(n628), .ZN(n630) );
  XNOR2_X1 U705 ( .A(n630), .B(n629), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U707 ( .A(n633), .B(KEYINPUT29), .ZN(n638) );
  INV_X1 U708 ( .A(G1961), .ZN(n925) );
  NOR2_X1 U709 ( .A1(n634), .A2(n925), .ZN(n636) );
  XNOR2_X1 U710 ( .A(G2078), .B(KEYINPUT25), .ZN(n902) );
  NOR2_X1 U711 ( .A1(n654), .A2(n902), .ZN(n635) );
  NOR2_X1 U712 ( .A1(n636), .A2(n635), .ZN(n645) );
  AND2_X1 U713 ( .A1(n645), .A2(G171), .ZN(n637) );
  NOR2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U715 ( .A(n639), .B(KEYINPUT99), .ZN(n660) );
  INV_X1 U716 ( .A(G8), .ZN(n640) );
  NOR2_X1 U717 ( .A1(n654), .A2(G2084), .ZN(n651) );
  NOR2_X1 U718 ( .A1(n640), .A2(n651), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U720 ( .A(KEYINPUT30), .B(n643), .ZN(n644) );
  NOR2_X1 U721 ( .A1(G168), .A2(n644), .ZN(n647) );
  NOR2_X1 U722 ( .A1(n645), .A2(G171), .ZN(n646) );
  XOR2_X1 U723 ( .A(KEYINPUT31), .B(n648), .Z(n659) );
  NOR2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n653) );
  NAND2_X1 U725 ( .A1(G8), .A2(n651), .ZN(n652) );
  NAND2_X1 U726 ( .A1(n653), .A2(n652), .ZN(n668) );
  NOR2_X1 U727 ( .A1(n654), .A2(G2090), .ZN(n656) );
  NOR2_X1 U728 ( .A1(G1971), .A2(n588), .ZN(n655) );
  NOR2_X1 U729 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U730 ( .A1(n657), .A2(G303), .ZN(n658) );
  OR2_X1 U731 ( .A1(n640), .A2(n658), .ZN(n662) );
  AND2_X1 U732 ( .A1(n659), .A2(n662), .ZN(n661) );
  NAND2_X1 U733 ( .A1(n661), .A2(n660), .ZN(n665) );
  INV_X1 U734 ( .A(n662), .ZN(n663) );
  OR2_X1 U735 ( .A1(n663), .A2(G286), .ZN(n664) );
  NAND2_X1 U736 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U737 ( .A(n666), .B(KEYINPUT32), .ZN(n667) );
  NAND2_X1 U738 ( .A1(n668), .A2(n667), .ZN(n684) );
  NOR2_X1 U739 ( .A1(G1971), .A2(G303), .ZN(n669) );
  XOR2_X1 U740 ( .A(KEYINPUT101), .B(n669), .Z(n671) );
  NOR2_X1 U741 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U742 ( .A1(n684), .A2(n672), .ZN(n675) );
  NAND2_X1 U743 ( .A1(G1976), .A2(G288), .ZN(n983) );
  NOR2_X1 U744 ( .A1(n588), .A2(n673), .ZN(n674) );
  NAND2_X1 U745 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U746 ( .A(n676), .B(KEYINPUT65), .ZN(n677) );
  NOR2_X1 U747 ( .A1(n677), .A2(KEYINPUT33), .ZN(n678) );
  NOR2_X1 U748 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U749 ( .A1(n681), .A2(n680), .ZN(n688) );
  NOR2_X1 U750 ( .A1(G2090), .A2(G303), .ZN(n682) );
  NAND2_X1 U751 ( .A1(G8), .A2(n682), .ZN(n683) );
  XNOR2_X1 U752 ( .A(n683), .B(KEYINPUT102), .ZN(n685) );
  NAND2_X1 U753 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U754 ( .A1(n588), .A2(n686), .ZN(n687) );
  NAND2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n693) );
  INV_X1 U756 ( .A(n689), .ZN(n690) );
  NOR2_X1 U757 ( .A1(n691), .A2(n690), .ZN(n741) );
  XNOR2_X1 U758 ( .A(G1986), .B(G290), .ZN(n982) );
  NAND2_X1 U759 ( .A1(n741), .A2(n982), .ZN(n692) );
  NAND2_X1 U760 ( .A1(n693), .A2(n692), .ZN(n726) );
  XNOR2_X1 U761 ( .A(KEYINPUT37), .B(G2067), .ZN(n738) );
  XNOR2_X1 U762 ( .A(KEYINPUT34), .B(KEYINPUT92), .ZN(n697) );
  NAND2_X1 U763 ( .A1(G104), .A2(n868), .ZN(n695) );
  NAND2_X1 U764 ( .A1(G140), .A2(n869), .ZN(n694) );
  NAND2_X1 U765 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U766 ( .A(n697), .B(n696), .ZN(n705) );
  XNOR2_X1 U767 ( .A(KEYINPUT94), .B(KEYINPUT35), .ZN(n703) );
  NAND2_X1 U768 ( .A1(n873), .A2(G128), .ZN(n701) );
  BUF_X1 U769 ( .A(n698), .Z(n876) );
  NAND2_X1 U770 ( .A1(G116), .A2(n876), .ZN(n699) );
  XOR2_X1 U771 ( .A(KEYINPUT93), .B(n699), .Z(n700) );
  NAND2_X1 U772 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U773 ( .A(n703), .B(n702), .Z(n704) );
  NOR2_X1 U774 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U775 ( .A(n706), .B(KEYINPUT36), .Z(n707) );
  XNOR2_X1 U776 ( .A(KEYINPUT95), .B(n707), .ZN(n892) );
  NOR2_X1 U777 ( .A1(n738), .A2(n892), .ZN(n965) );
  NAND2_X1 U778 ( .A1(n741), .A2(n965), .ZN(n736) );
  NAND2_X1 U779 ( .A1(G141), .A2(n869), .ZN(n709) );
  NAND2_X1 U780 ( .A1(G117), .A2(n876), .ZN(n708) );
  NAND2_X1 U781 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U782 ( .A1(n868), .A2(G105), .ZN(n710) );
  XOR2_X1 U783 ( .A(KEYINPUT38), .B(n710), .Z(n711) );
  NOR2_X1 U784 ( .A1(n712), .A2(n711), .ZN(n714) );
  NAND2_X1 U785 ( .A1(n873), .A2(G129), .ZN(n713) );
  NAND2_X1 U786 ( .A1(n714), .A2(n713), .ZN(n882) );
  NAND2_X1 U787 ( .A1(G1996), .A2(n882), .ZN(n715) );
  XNOR2_X1 U788 ( .A(n715), .B(KEYINPUT97), .ZN(n723) );
  NAND2_X1 U789 ( .A1(G95), .A2(n868), .ZN(n717) );
  NAND2_X1 U790 ( .A1(G131), .A2(n869), .ZN(n716) );
  NAND2_X1 U791 ( .A1(n717), .A2(n716), .ZN(n721) );
  NAND2_X1 U792 ( .A1(n873), .A2(G119), .ZN(n719) );
  NAND2_X1 U793 ( .A1(G107), .A2(n876), .ZN(n718) );
  NAND2_X1 U794 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U795 ( .A1(n721), .A2(n720), .ZN(n887) );
  XOR2_X1 U796 ( .A(KEYINPUT96), .B(G1991), .Z(n911) );
  NOR2_X1 U797 ( .A1(n887), .A2(n911), .ZN(n722) );
  NOR2_X1 U798 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U799 ( .A(KEYINPUT98), .B(n724), .Z(n961) );
  NAND2_X1 U800 ( .A1(n741), .A2(n961), .ZN(n728) );
  NAND2_X1 U801 ( .A1(n736), .A2(n728), .ZN(n725) );
  XNOR2_X1 U802 ( .A(n727), .B(KEYINPUT103), .ZN(n743) );
  NOR2_X1 U803 ( .A1(G1996), .A2(n882), .ZN(n957) );
  INV_X1 U804 ( .A(n728), .ZN(n732) );
  NOR2_X1 U805 ( .A1(G1986), .A2(G290), .ZN(n730) );
  NAND2_X1 U806 ( .A1(n911), .A2(n887), .ZN(n729) );
  XOR2_X1 U807 ( .A(KEYINPUT104), .B(n729), .Z(n955) );
  NOR2_X1 U808 ( .A1(n730), .A2(n955), .ZN(n731) );
  NOR2_X1 U809 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U810 ( .A(KEYINPUT105), .B(n733), .Z(n734) );
  NOR2_X1 U811 ( .A1(n957), .A2(n734), .ZN(n735) );
  XNOR2_X1 U812 ( .A(n735), .B(KEYINPUT39), .ZN(n737) );
  NAND2_X1 U813 ( .A1(n737), .A2(n736), .ZN(n739) );
  NAND2_X1 U814 ( .A1(n738), .A2(n892), .ZN(n974) );
  NAND2_X1 U815 ( .A1(n739), .A2(n974), .ZN(n740) );
  NAND2_X1 U816 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U817 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U818 ( .A(n744), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U819 ( .A(G2443), .B(G2446), .Z(n746) );
  XNOR2_X1 U820 ( .A(G2427), .B(G2451), .ZN(n745) );
  XNOR2_X1 U821 ( .A(n746), .B(n745), .ZN(n752) );
  XOR2_X1 U822 ( .A(G2430), .B(G2454), .Z(n748) );
  XNOR2_X1 U823 ( .A(G1341), .B(G1348), .ZN(n747) );
  XNOR2_X1 U824 ( .A(n748), .B(n747), .ZN(n750) );
  XOR2_X1 U825 ( .A(G2435), .B(G2438), .Z(n749) );
  XNOR2_X1 U826 ( .A(n750), .B(n749), .ZN(n751) );
  XOR2_X1 U827 ( .A(n752), .B(n751), .Z(n753) );
  AND2_X1 U828 ( .A1(G14), .A2(n753), .ZN(G401) );
  AND2_X1 U829 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U830 ( .A(G57), .ZN(G237) );
  INV_X1 U831 ( .A(n798), .ZN(G299) );
  XOR2_X1 U832 ( .A(KEYINPUT10), .B(KEYINPUT75), .Z(n755) );
  NAND2_X1 U833 ( .A1(G7), .A2(G661), .ZN(n754) );
  XNOR2_X1 U834 ( .A(n755), .B(n754), .ZN(G223) );
  XOR2_X1 U835 ( .A(KEYINPUT76), .B(KEYINPUT11), .Z(n757) );
  INV_X1 U836 ( .A(G223), .ZN(n824) );
  NAND2_X1 U837 ( .A1(G567), .A2(n824), .ZN(n756) );
  XNOR2_X1 U838 ( .A(n757), .B(n756), .ZN(G234) );
  INV_X1 U839 ( .A(G860), .ZN(n762) );
  OR2_X1 U840 ( .A1(n993), .A2(n762), .ZN(G153) );
  INV_X1 U841 ( .A(G171), .ZN(G301) );
  NAND2_X1 U842 ( .A1(G301), .A2(G868), .ZN(n759) );
  INV_X1 U843 ( .A(G868), .ZN(n805) );
  NAND2_X1 U844 ( .A1(n994), .A2(n805), .ZN(n758) );
  NAND2_X1 U845 ( .A1(n759), .A2(n758), .ZN(G284) );
  NOR2_X1 U846 ( .A1(G286), .A2(n805), .ZN(n761) );
  NOR2_X1 U847 ( .A1(G868), .A2(G299), .ZN(n760) );
  NOR2_X1 U848 ( .A1(n761), .A2(n760), .ZN(G297) );
  NAND2_X1 U849 ( .A1(n762), .A2(G559), .ZN(n763) );
  INV_X1 U850 ( .A(n994), .ZN(n779) );
  NAND2_X1 U851 ( .A1(n763), .A2(n779), .ZN(n764) );
  XNOR2_X1 U852 ( .A(n764), .B(KEYINPUT16), .ZN(n765) );
  XOR2_X1 U853 ( .A(KEYINPUT79), .B(n765), .Z(G148) );
  NOR2_X1 U854 ( .A1(n994), .A2(n805), .ZN(n766) );
  XOR2_X1 U855 ( .A(KEYINPUT80), .B(n766), .Z(n767) );
  NOR2_X1 U856 ( .A1(G559), .A2(n767), .ZN(n769) );
  NOR2_X1 U857 ( .A1(G868), .A2(n993), .ZN(n768) );
  NOR2_X1 U858 ( .A1(n769), .A2(n768), .ZN(G282) );
  NAND2_X1 U859 ( .A1(G135), .A2(n869), .ZN(n771) );
  NAND2_X1 U860 ( .A1(G111), .A2(n876), .ZN(n770) );
  NAND2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n873), .A2(G123), .ZN(n772) );
  XOR2_X1 U863 ( .A(KEYINPUT18), .B(n772), .Z(n773) );
  NOR2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n868), .A2(G99), .ZN(n775) );
  NAND2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n952) );
  XOR2_X1 U867 ( .A(n952), .B(G2096), .Z(n778) );
  XNOR2_X1 U868 ( .A(G2100), .B(KEYINPUT81), .ZN(n777) );
  NAND2_X1 U869 ( .A1(n778), .A2(n777), .ZN(G156) );
  NAND2_X1 U870 ( .A1(G559), .A2(n779), .ZN(n780) );
  XNOR2_X1 U871 ( .A(n780), .B(KEYINPUT82), .ZN(n803) );
  XNOR2_X1 U872 ( .A(n803), .B(n993), .ZN(n781) );
  NOR2_X1 U873 ( .A1(n781), .A2(G860), .ZN(n794) );
  NAND2_X1 U874 ( .A1(G93), .A2(n782), .ZN(n785) );
  NAND2_X1 U875 ( .A1(G80), .A2(n783), .ZN(n784) );
  NAND2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U877 ( .A(n786), .B(KEYINPUT83), .ZN(n789) );
  NAND2_X1 U878 ( .A1(G67), .A2(n787), .ZN(n788) );
  NAND2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n793) );
  NAND2_X1 U880 ( .A1(n790), .A2(G55), .ZN(n791) );
  XOR2_X1 U881 ( .A(KEYINPUT84), .B(n791), .Z(n792) );
  OR2_X1 U882 ( .A1(n793), .A2(n792), .ZN(n806) );
  XOR2_X1 U883 ( .A(n794), .B(n806), .Z(G145) );
  XOR2_X1 U884 ( .A(KEYINPUT19), .B(n806), .Z(n796) );
  XNOR2_X1 U885 ( .A(G288), .B(KEYINPUT87), .ZN(n795) );
  XNOR2_X1 U886 ( .A(n796), .B(n795), .ZN(n797) );
  XNOR2_X1 U887 ( .A(G166), .B(n797), .ZN(n800) );
  XNOR2_X1 U888 ( .A(n993), .B(n798), .ZN(n799) );
  XNOR2_X1 U889 ( .A(n800), .B(n799), .ZN(n801) );
  XOR2_X1 U890 ( .A(n801), .B(G290), .Z(n802) );
  XNOR2_X1 U891 ( .A(G305), .B(n802), .ZN(n830) );
  XNOR2_X1 U892 ( .A(n803), .B(n830), .ZN(n804) );
  NOR2_X1 U893 ( .A1(n805), .A2(n804), .ZN(n808) );
  NOR2_X1 U894 ( .A1(G868), .A2(n806), .ZN(n807) );
  NOR2_X1 U895 ( .A1(n808), .A2(n807), .ZN(G295) );
  NAND2_X1 U896 ( .A1(G2078), .A2(G2084), .ZN(n809) );
  XOR2_X1 U897 ( .A(KEYINPUT20), .B(n809), .Z(n810) );
  NAND2_X1 U898 ( .A1(G2090), .A2(n810), .ZN(n811) );
  XNOR2_X1 U899 ( .A(KEYINPUT21), .B(n811), .ZN(n812) );
  NAND2_X1 U900 ( .A1(n812), .A2(G2072), .ZN(n813) );
  XNOR2_X1 U901 ( .A(KEYINPUT88), .B(n813), .ZN(G158) );
  XOR2_X1 U902 ( .A(KEYINPUT74), .B(G82), .Z(G220) );
  XNOR2_X1 U903 ( .A(KEYINPUT73), .B(G132), .ZN(G219) );
  XNOR2_X1 U904 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U905 ( .A1(G220), .A2(G219), .ZN(n815) );
  XNOR2_X1 U906 ( .A(KEYINPUT22), .B(KEYINPUT89), .ZN(n814) );
  XNOR2_X1 U907 ( .A(n815), .B(n814), .ZN(n816) );
  NOR2_X1 U908 ( .A1(n816), .A2(G218), .ZN(n817) );
  NAND2_X1 U909 ( .A1(G96), .A2(n817), .ZN(n828) );
  NAND2_X1 U910 ( .A1(n828), .A2(G2106), .ZN(n822) );
  NAND2_X1 U911 ( .A1(G120), .A2(G69), .ZN(n818) );
  NOR2_X1 U912 ( .A1(G237), .A2(n818), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n819), .A2(G108), .ZN(n820) );
  XNOR2_X1 U914 ( .A(n820), .B(KEYINPUT90), .ZN(n829) );
  NAND2_X1 U915 ( .A1(n829), .A2(G567), .ZN(n821) );
  NAND2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n901) );
  NAND2_X1 U917 ( .A1(G483), .A2(G661), .ZN(n823) );
  NOR2_X1 U918 ( .A1(n901), .A2(n823), .ZN(n827) );
  NAND2_X1 U919 ( .A1(n827), .A2(G36), .ZN(G176) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n824), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n825) );
  NAND2_X1 U922 ( .A1(G661), .A2(n825), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U924 ( .A1(n827), .A2(n826), .ZN(G188) );
  XOR2_X1 U925 ( .A(G69), .B(KEYINPUT106), .Z(G235) );
  INV_X1 U927 ( .A(G120), .ZN(G236) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  NOR2_X1 U929 ( .A1(n829), .A2(n828), .ZN(G325) );
  INV_X1 U930 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U931 ( .A(G286), .B(n994), .ZN(n831) );
  XNOR2_X1 U932 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U933 ( .A(n832), .B(G171), .ZN(n833) );
  NOR2_X1 U934 ( .A1(G37), .A2(n833), .ZN(G397) );
  XOR2_X1 U935 ( .A(KEYINPUT41), .B(G1976), .Z(n835) );
  XNOR2_X1 U936 ( .A(G1986), .B(G1971), .ZN(n834) );
  XNOR2_X1 U937 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U938 ( .A(n836), .B(KEYINPUT108), .Z(n838) );
  XNOR2_X1 U939 ( .A(G1996), .B(G1991), .ZN(n837) );
  XNOR2_X1 U940 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U941 ( .A(G1981), .B(G1956), .Z(n840) );
  XNOR2_X1 U942 ( .A(G1966), .B(G1961), .ZN(n839) );
  XNOR2_X1 U943 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U944 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U945 ( .A(KEYINPUT107), .B(G2474), .ZN(n843) );
  XNOR2_X1 U946 ( .A(n844), .B(n843), .ZN(G229) );
  XOR2_X1 U947 ( .A(G2100), .B(G2096), .Z(n846) );
  XNOR2_X1 U948 ( .A(KEYINPUT42), .B(G2678), .ZN(n845) );
  XNOR2_X1 U949 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U950 ( .A(KEYINPUT43), .B(G2090), .Z(n848) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2072), .ZN(n847) );
  XNOR2_X1 U952 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U953 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U954 ( .A(G2078), .B(G2084), .ZN(n851) );
  XNOR2_X1 U955 ( .A(n852), .B(n851), .ZN(G227) );
  NAND2_X1 U956 ( .A1(G124), .A2(n873), .ZN(n853) );
  XNOR2_X1 U957 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U958 ( .A1(G112), .A2(n876), .ZN(n854) );
  NAND2_X1 U959 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U960 ( .A1(G100), .A2(n868), .ZN(n857) );
  NAND2_X1 U961 ( .A1(G136), .A2(n869), .ZN(n856) );
  NAND2_X1 U962 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U963 ( .A1(n859), .A2(n858), .ZN(G162) );
  NAND2_X1 U964 ( .A1(G103), .A2(n868), .ZN(n861) );
  NAND2_X1 U965 ( .A1(G139), .A2(n869), .ZN(n860) );
  NAND2_X1 U966 ( .A1(n861), .A2(n860), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n873), .A2(G127), .ZN(n863) );
  NAND2_X1 U968 ( .A1(G115), .A2(n876), .ZN(n862) );
  NAND2_X1 U969 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U970 ( .A(KEYINPUT111), .B(n864), .ZN(n865) );
  XNOR2_X1 U971 ( .A(KEYINPUT47), .B(n865), .ZN(n866) );
  NOR2_X1 U972 ( .A1(n867), .A2(n866), .ZN(n967) );
  XNOR2_X1 U973 ( .A(G160), .B(n967), .ZN(n891) );
  NAND2_X1 U974 ( .A1(G106), .A2(n868), .ZN(n871) );
  NAND2_X1 U975 ( .A1(G142), .A2(n869), .ZN(n870) );
  NAND2_X1 U976 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U977 ( .A(n872), .B(KEYINPUT45), .ZN(n875) );
  NAND2_X1 U978 ( .A1(G130), .A2(n873), .ZN(n874) );
  NAND2_X1 U979 ( .A1(n875), .A2(n874), .ZN(n879) );
  NAND2_X1 U980 ( .A1(G118), .A2(n876), .ZN(n877) );
  XNOR2_X1 U981 ( .A(KEYINPUT109), .B(n877), .ZN(n878) );
  NOR2_X1 U982 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U983 ( .A(G162), .B(n880), .Z(n881) );
  XNOR2_X1 U984 ( .A(n952), .B(n881), .ZN(n886) );
  XNOR2_X1 U985 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n882), .B(KEYINPUT110), .ZN(n883) );
  XNOR2_X1 U987 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U988 ( .A(n886), .B(n885), .Z(n889) );
  XNOR2_X1 U989 ( .A(G164), .B(n887), .ZN(n888) );
  XNOR2_X1 U990 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n891), .B(n890), .ZN(n893) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U993 ( .A1(G37), .A2(n894), .ZN(G395) );
  NOR2_X1 U994 ( .A1(G229), .A2(G227), .ZN(n895) );
  XNOR2_X1 U995 ( .A(KEYINPUT49), .B(n895), .ZN(n896) );
  NOR2_X1 U996 ( .A1(G397), .A2(n896), .ZN(n900) );
  NOR2_X1 U997 ( .A1(n901), .A2(G401), .ZN(n897) );
  XOR2_X1 U998 ( .A(KEYINPUT112), .B(n897), .Z(n898) );
  NOR2_X1 U999 ( .A1(G395), .A2(n898), .ZN(n899) );
  NAND2_X1 U1000 ( .A1(n900), .A2(n899), .ZN(G225) );
  INV_X1 U1001 ( .A(G225), .ZN(G308) );
  INV_X1 U1002 ( .A(n901), .ZN(G319) );
  INV_X1 U1003 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1004 ( .A(G29), .B(KEYINPUT120), .Z(n924) );
  XNOR2_X1 U1005 ( .A(G27), .B(n902), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(G2067), .B(G26), .ZN(n904) );
  XNOR2_X1 U1007 ( .A(G33), .B(G2072), .ZN(n903) );
  NOR2_X1 U1008 ( .A1(n904), .A2(n903), .ZN(n905) );
  NAND2_X1 U1009 ( .A1(n906), .A2(n905), .ZN(n908) );
  XNOR2_X1 U1010 ( .A(G32), .B(G1996), .ZN(n907) );
  NOR2_X1 U1011 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1012 ( .A(KEYINPUT118), .B(n909), .ZN(n910) );
  NAND2_X1 U1013 ( .A1(n910), .A2(G28), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(KEYINPUT117), .B(n911), .ZN(n912) );
  XNOR2_X1 U1015 ( .A(G25), .B(n912), .ZN(n913) );
  NOR2_X1 U1016 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1017 ( .A(n915), .B(KEYINPUT53), .ZN(n916) );
  XNOR2_X1 U1018 ( .A(n916), .B(KEYINPUT119), .ZN(n919) );
  XOR2_X1 U1019 ( .A(G2084), .B(G34), .Z(n917) );
  XNOR2_X1 U1020 ( .A(KEYINPUT54), .B(n917), .ZN(n918) );
  NAND2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(G35), .B(G2090), .ZN(n920) );
  NOR2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1024 ( .A(n922), .B(KEYINPUT55), .ZN(n923) );
  NAND2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n1012) );
  XNOR2_X1 U1026 ( .A(G5), .B(n925), .ZN(n944) );
  XNOR2_X1 U1027 ( .A(G1986), .B(G24), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(G1971), .B(G22), .ZN(n927) );
  XNOR2_X1 U1029 ( .A(G1976), .B(G23), .ZN(n926) );
  NOR2_X1 U1030 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1031 ( .A(KEYINPUT125), .B(n928), .ZN(n929) );
  NOR2_X1 U1032 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1033 ( .A(KEYINPUT58), .B(n931), .Z(n942) );
  XNOR2_X1 U1034 ( .A(G20), .B(n932), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(G1341), .B(G19), .ZN(n934) );
  XNOR2_X1 U1036 ( .A(G1981), .B(G6), .ZN(n933) );
  NOR2_X1 U1037 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n939) );
  XOR2_X1 U1039 ( .A(KEYINPUT59), .B(G1348), .Z(n937) );
  XNOR2_X1 U1040 ( .A(G4), .B(n937), .ZN(n938) );
  NOR2_X1 U1041 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1042 ( .A(KEYINPUT60), .B(n940), .Z(n941) );
  NOR2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n947) );
  XNOR2_X1 U1045 ( .A(G21), .B(G1966), .ZN(n945) );
  XNOR2_X1 U1046 ( .A(KEYINPUT124), .B(n945), .ZN(n946) );
  NOR2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1048 ( .A(KEYINPUT61), .B(n948), .Z(n949) );
  NOR2_X1 U1049 ( .A1(G16), .A2(n949), .ZN(n950) );
  XOR2_X1 U1050 ( .A(KEYINPUT126), .B(n950), .Z(n951) );
  NAND2_X1 U1051 ( .A1(G11), .A2(n951), .ZN(n1010) );
  INV_X1 U1052 ( .A(KEYINPUT55), .ZN(n979) );
  XOR2_X1 U1053 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n977) );
  XNOR2_X1 U1054 ( .A(G160), .B(G2084), .ZN(n953) );
  NAND2_X1 U1055 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1056 ( .A1(n955), .A2(n954), .ZN(n963) );
  XOR2_X1 U1057 ( .A(G2090), .B(G162), .Z(n956) );
  NOR2_X1 U1058 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1059 ( .A(KEYINPUT113), .B(n958), .Z(n959) );
  XNOR2_X1 U1060 ( .A(n959), .B(KEYINPUT51), .ZN(n960) );
  NOR2_X1 U1061 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1062 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1064 ( .A(KEYINPUT114), .B(n966), .Z(n973) );
  XOR2_X1 U1065 ( .A(n967), .B(KEYINPUT115), .Z(n968) );
  XOR2_X1 U1066 ( .A(G2072), .B(n968), .Z(n970) );
  XOR2_X1 U1067 ( .A(G164), .B(G2078), .Z(n969) );
  NOR2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1069 ( .A(KEYINPUT50), .B(n971), .Z(n972) );
  NOR2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1072 ( .A(n977), .B(n976), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n980), .A2(G29), .ZN(n1008) );
  XNOR2_X1 U1075 ( .A(G16), .B(KEYINPUT56), .ZN(n1006) );
  XNOR2_X1 U1076 ( .A(G1956), .B(G299), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(G1971), .B(G303), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(KEYINPUT122), .B(n985), .ZN(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n1003) );
  XNOR2_X1 U1083 ( .A(G1966), .B(G168), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(n992), .B(KEYINPUT57), .ZN(n1001) );
  XNOR2_X1 U1086 ( .A(n993), .B(G1341), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(n994), .B(G1348), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(G301), .B(G1961), .ZN(n995) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1090 ( .A(KEYINPUT121), .B(n997), .ZN(n998) );
  NOR2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(KEYINPUT123), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(n1013), .B(KEYINPUT62), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(KEYINPUT127), .B(n1014), .ZN(G311) );
  INV_X1 U1101 ( .A(G311), .ZN(G150) );
endmodule

