

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(G651), .A2(n639), .ZN(n659) );
  XOR2_X1 U556 ( .A(n724), .B(KEYINPUT93), .Z(n786) );
  NOR2_X1 U557 ( .A1(n769), .A2(n728), .ZN(n729) );
  INV_X1 U558 ( .A(KEYINPUT31), .ZN(n737) );
  XNOR2_X1 U559 ( .A(n738), .B(n737), .ZN(n767) );
  NAND2_X1 U560 ( .A1(n767), .A2(n766), .ZN(n772) );
  INV_X1 U561 ( .A(KEYINPUT96), .ZN(n794) );
  XNOR2_X1 U562 ( .A(n795), .B(n794), .ZN(n796) );
  NAND2_X1 U563 ( .A1(n773), .A2(G8), .ZN(n724) );
  NOR2_X1 U564 ( .A1(G164), .A2(G1384), .ZN(n721) );
  NOR2_X1 U565 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U566 ( .A1(n552), .A2(n551), .ZN(G160) );
  XNOR2_X1 U567 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n522) );
  NOR2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  XNOR2_X2 U569 ( .A(n522), .B(n521), .ZN(n875) );
  NAND2_X1 U570 ( .A1(G138), .A2(n875), .ZN(n524) );
  INV_X1 U571 ( .A(G2104), .ZN(n525) );
  NOR2_X4 U572 ( .A1(G2105), .A2(n525), .ZN(n883) );
  NAND2_X1 U573 ( .A1(G102), .A2(n883), .ZN(n523) );
  NAND2_X1 U574 ( .A1(n524), .A2(n523), .ZN(n529) );
  AND2_X1 U575 ( .A1(n525), .A2(G2105), .ZN(n877) );
  NAND2_X1 U576 ( .A1(G126), .A2(n877), .ZN(n527) );
  AND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n878) );
  NAND2_X1 U578 ( .A1(G114), .A2(n878), .ZN(n526) );
  NAND2_X1 U579 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U580 ( .A1(n529), .A2(n528), .ZN(G164) );
  INV_X1 U581 ( .A(G651), .ZN(n537) );
  NOR2_X1 U582 ( .A1(G543), .A2(n537), .ZN(n531) );
  XNOR2_X1 U583 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n530) );
  XNOR2_X1 U584 ( .A(n531), .B(n530), .ZN(n650) );
  NAND2_X1 U585 ( .A1(G63), .A2(n650), .ZN(n533) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n639) );
  NAND2_X1 U587 ( .A1(G51), .A2(n659), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U589 ( .A(KEYINPUT6), .B(n534), .ZN(n543) );
  NOR2_X1 U590 ( .A1(G543), .A2(G651), .ZN(n535) );
  XNOR2_X1 U591 ( .A(n535), .B(KEYINPUT64), .ZN(n651) );
  NAND2_X1 U592 ( .A1(G89), .A2(n651), .ZN(n536) );
  XNOR2_X1 U593 ( .A(n536), .B(KEYINPUT4), .ZN(n539) );
  NOR2_X1 U594 ( .A1(n639), .A2(n537), .ZN(n654) );
  NAND2_X1 U595 ( .A1(G76), .A2(n654), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U597 ( .A(KEYINPUT74), .B(n540), .Z(n541) );
  XNOR2_X1 U598 ( .A(KEYINPUT5), .B(n541), .ZN(n542) );
  NOR2_X1 U599 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U600 ( .A(KEYINPUT7), .B(n544), .Z(G168) );
  XNOR2_X1 U601 ( .A(G168), .B(KEYINPUT8), .ZN(n545) );
  XNOR2_X1 U602 ( .A(n545), .B(KEYINPUT75), .ZN(G286) );
  NAND2_X1 U603 ( .A1(n877), .A2(G125), .ZN(n548) );
  NAND2_X1 U604 ( .A1(G101), .A2(n883), .ZN(n546) );
  XOR2_X1 U605 ( .A(KEYINPUT23), .B(n546), .Z(n547) );
  NAND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n552) );
  NAND2_X1 U607 ( .A1(G137), .A2(n875), .ZN(n550) );
  NAND2_X1 U608 ( .A1(G113), .A2(n878), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U610 ( .A(G2451), .B(G2427), .ZN(n562) );
  XOR2_X1 U611 ( .A(G2430), .B(G2443), .Z(n554) );
  XNOR2_X1 U612 ( .A(KEYINPUT101), .B(G2438), .ZN(n553) );
  XNOR2_X1 U613 ( .A(n554), .B(n553), .ZN(n558) );
  XOR2_X1 U614 ( .A(G2435), .B(G2454), .Z(n556) );
  XNOR2_X1 U615 ( .A(G1341), .B(G1348), .ZN(n555) );
  XNOR2_X1 U616 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U617 ( .A(n558), .B(n557), .Z(n560) );
  XNOR2_X1 U618 ( .A(G2446), .B(KEYINPUT102), .ZN(n559) );
  XNOR2_X1 U619 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U620 ( .A(n562), .B(n561), .ZN(n563) );
  AND2_X1 U621 ( .A1(n563), .A2(G14), .ZN(G401) );
  NAND2_X1 U622 ( .A1(G64), .A2(n650), .ZN(n565) );
  NAND2_X1 U623 ( .A1(G52), .A2(n659), .ZN(n564) );
  NAND2_X1 U624 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U625 ( .A(KEYINPUT69), .B(n566), .Z(n571) );
  NAND2_X1 U626 ( .A1(n654), .A2(G77), .ZN(n568) );
  NAND2_X1 U627 ( .A1(G90), .A2(n651), .ZN(n567) );
  NAND2_X1 U628 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U629 ( .A(KEYINPUT9), .B(n569), .Z(n570) );
  NOR2_X1 U630 ( .A1(n571), .A2(n570), .ZN(G171) );
  AND2_X1 U631 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U632 ( .A(G57), .ZN(G237) );
  INV_X1 U633 ( .A(G132), .ZN(G219) );
  INV_X1 U634 ( .A(G82), .ZN(G220) );
  NAND2_X1 U635 ( .A1(G62), .A2(n650), .ZN(n573) );
  NAND2_X1 U636 ( .A1(G50), .A2(n659), .ZN(n572) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT80), .B(n574), .Z(n578) );
  NAND2_X1 U639 ( .A1(n651), .A2(G88), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n654), .A2(G75), .ZN(n575) );
  AND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(G303) );
  NAND2_X1 U643 ( .A1(G7), .A2(G661), .ZN(n579) );
  XOR2_X1 U644 ( .A(n579), .B(KEYINPUT10), .Z(n912) );
  NAND2_X1 U645 ( .A1(n912), .A2(G567), .ZN(n580) );
  XOR2_X1 U646 ( .A(KEYINPUT11), .B(n580), .Z(G234) );
  NAND2_X1 U647 ( .A1(G56), .A2(n650), .ZN(n581) );
  XOR2_X1 U648 ( .A(KEYINPUT14), .B(n581), .Z(n587) );
  NAND2_X1 U649 ( .A1(G81), .A2(n651), .ZN(n582) );
  XNOR2_X1 U650 ( .A(n582), .B(KEYINPUT12), .ZN(n584) );
  NAND2_X1 U651 ( .A1(G68), .A2(n654), .ZN(n583) );
  NAND2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U653 ( .A(KEYINPUT13), .B(n585), .Z(n586) );
  NOR2_X1 U654 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U655 ( .A1(n659), .A2(G43), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n975) );
  INV_X1 U657 ( .A(G860), .ZN(n611) );
  OR2_X1 U658 ( .A1(n975), .A2(n611), .ZN(G153) );
  INV_X1 U659 ( .A(G171), .ZN(G301) );
  NAND2_X1 U660 ( .A1(G868), .A2(G301), .ZN(n600) );
  NAND2_X1 U661 ( .A1(G66), .A2(n650), .ZN(n590) );
  XNOR2_X1 U662 ( .A(n590), .B(KEYINPUT72), .ZN(n597) );
  NAND2_X1 U663 ( .A1(n654), .A2(G79), .ZN(n592) );
  NAND2_X1 U664 ( .A1(G92), .A2(n651), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U666 ( .A1(G54), .A2(n659), .ZN(n593) );
  XNOR2_X1 U667 ( .A(KEYINPUT73), .B(n593), .ZN(n594) );
  NOR2_X1 U668 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U669 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U670 ( .A(KEYINPUT15), .B(n598), .ZN(n970) );
  INV_X1 U671 ( .A(n970), .ZN(n756) );
  INV_X1 U672 ( .A(G868), .ZN(n671) );
  NAND2_X1 U673 ( .A1(n756), .A2(n671), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(G284) );
  NAND2_X1 U675 ( .A1(n654), .A2(G78), .ZN(n602) );
  NAND2_X1 U676 ( .A1(G91), .A2(n651), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U678 ( .A(KEYINPUT70), .B(n603), .ZN(n606) );
  NAND2_X1 U679 ( .A1(G65), .A2(n650), .ZN(n604) );
  XNOR2_X1 U680 ( .A(KEYINPUT71), .B(n604), .ZN(n605) );
  NOR2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n659), .A2(G53), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n608), .A2(n607), .ZN(G299) );
  NOR2_X1 U684 ( .A1(G286), .A2(n671), .ZN(n610) );
  NOR2_X1 U685 ( .A1(G868), .A2(G299), .ZN(n609) );
  NOR2_X1 U686 ( .A1(n610), .A2(n609), .ZN(G297) );
  NAND2_X1 U687 ( .A1(n611), .A2(G559), .ZN(n612) );
  NAND2_X1 U688 ( .A1(n612), .A2(n970), .ZN(n613) );
  XNOR2_X1 U689 ( .A(n613), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U690 ( .A1(G868), .A2(n975), .ZN(n616) );
  NAND2_X1 U691 ( .A1(G868), .A2(n970), .ZN(n614) );
  NOR2_X1 U692 ( .A1(G559), .A2(n614), .ZN(n615) );
  NOR2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U694 ( .A(KEYINPUT76), .B(n617), .ZN(G282) );
  NAND2_X1 U695 ( .A1(G123), .A2(n877), .ZN(n618) );
  XOR2_X1 U696 ( .A(KEYINPUT77), .B(n618), .Z(n619) );
  XNOR2_X1 U697 ( .A(n619), .B(KEYINPUT18), .ZN(n621) );
  NAND2_X1 U698 ( .A1(G99), .A2(n883), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G135), .A2(n875), .ZN(n623) );
  NAND2_X1 U701 ( .A1(G111), .A2(n878), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n919) );
  XNOR2_X1 U704 ( .A(G2096), .B(n919), .ZN(n626) );
  INV_X1 U705 ( .A(G2100), .ZN(n838) );
  NAND2_X1 U706 ( .A1(n626), .A2(n838), .ZN(G156) );
  NAND2_X1 U707 ( .A1(G559), .A2(n970), .ZN(n627) );
  XNOR2_X1 U708 ( .A(n627), .B(n975), .ZN(n669) );
  NOR2_X1 U709 ( .A1(G860), .A2(n669), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n650), .A2(G67), .ZN(n629) );
  NAND2_X1 U711 ( .A1(G93), .A2(n651), .ZN(n628) );
  NAND2_X1 U712 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U713 ( .A1(G80), .A2(n654), .ZN(n631) );
  NAND2_X1 U714 ( .A1(G55), .A2(n659), .ZN(n630) );
  NAND2_X1 U715 ( .A1(n631), .A2(n630), .ZN(n632) );
  OR2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n672) );
  XOR2_X1 U717 ( .A(n672), .B(KEYINPUT78), .Z(n634) );
  XNOR2_X1 U718 ( .A(n635), .B(n634), .ZN(G145) );
  NAND2_X1 U719 ( .A1(G49), .A2(n659), .ZN(n637) );
  NAND2_X1 U720 ( .A1(G74), .A2(G651), .ZN(n636) );
  NAND2_X1 U721 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U722 ( .A1(n650), .A2(n638), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n639), .A2(G87), .ZN(n640) );
  NAND2_X1 U724 ( .A1(n641), .A2(n640), .ZN(G288) );
  NAND2_X1 U725 ( .A1(n650), .A2(G60), .ZN(n648) );
  NAND2_X1 U726 ( .A1(G72), .A2(n654), .ZN(n643) );
  NAND2_X1 U727 ( .A1(G47), .A2(n659), .ZN(n642) );
  NAND2_X1 U728 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U729 ( .A1(n651), .A2(G85), .ZN(n644) );
  XOR2_X1 U730 ( .A(KEYINPUT66), .B(n644), .Z(n645) );
  NOR2_X1 U731 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U732 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U733 ( .A(n649), .B(KEYINPUT68), .ZN(G290) );
  NAND2_X1 U734 ( .A1(n650), .A2(G61), .ZN(n653) );
  NAND2_X1 U735 ( .A1(G86), .A2(n651), .ZN(n652) );
  NAND2_X1 U736 ( .A1(n653), .A2(n652), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n654), .A2(G73), .ZN(n655) );
  XOR2_X1 U738 ( .A(KEYINPUT2), .B(n655), .Z(n656) );
  NOR2_X1 U739 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U740 ( .A(KEYINPUT79), .B(n658), .Z(n661) );
  NAND2_X1 U741 ( .A1(n659), .A2(G48), .ZN(n660) );
  NAND2_X1 U742 ( .A1(n661), .A2(n660), .ZN(G305) );
  XNOR2_X1 U743 ( .A(KEYINPUT82), .B(KEYINPUT19), .ZN(n663) );
  XNOR2_X1 U744 ( .A(G288), .B(KEYINPUT81), .ZN(n662) );
  XNOR2_X1 U745 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U746 ( .A(n664), .B(n672), .ZN(n666) );
  XOR2_X1 U747 ( .A(G290), .B(G299), .Z(n665) );
  XNOR2_X1 U748 ( .A(n666), .B(n665), .ZN(n667) );
  XOR2_X1 U749 ( .A(G303), .B(n667), .Z(n668) );
  XNOR2_X1 U750 ( .A(n668), .B(G305), .ZN(n899) );
  XNOR2_X1 U751 ( .A(n669), .B(n899), .ZN(n670) );
  NAND2_X1 U752 ( .A1(n670), .A2(G868), .ZN(n674) );
  NAND2_X1 U753 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U754 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U757 ( .A1(G2090), .A2(n676), .ZN(n678) );
  XOR2_X1 U758 ( .A(KEYINPUT83), .B(KEYINPUT21), .Z(n677) );
  XNOR2_X1 U759 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U760 ( .A1(G2072), .A2(n679), .ZN(G158) );
  XNOR2_X1 U761 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U762 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U763 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U764 ( .A1(G218), .A2(n681), .ZN(n682) );
  XNOR2_X1 U765 ( .A(KEYINPUT84), .B(n682), .ZN(n683) );
  NAND2_X1 U766 ( .A1(n683), .A2(G96), .ZN(n831) );
  NAND2_X1 U767 ( .A1(n831), .A2(G2106), .ZN(n687) );
  NAND2_X1 U768 ( .A1(G108), .A2(G120), .ZN(n684) );
  NOR2_X1 U769 ( .A1(G237), .A2(n684), .ZN(n685) );
  NAND2_X1 U770 ( .A1(G69), .A2(n685), .ZN(n832) );
  NAND2_X1 U771 ( .A1(n832), .A2(G567), .ZN(n686) );
  NAND2_X1 U772 ( .A1(n687), .A2(n686), .ZN(n911) );
  NAND2_X1 U773 ( .A1(G661), .A2(G483), .ZN(n688) );
  NOR2_X1 U774 ( .A1(n911), .A2(n688), .ZN(n830) );
  NAND2_X1 U775 ( .A1(G36), .A2(n830), .ZN(n689) );
  XOR2_X1 U776 ( .A(KEYINPUT85), .B(n689), .Z(G176) );
  XOR2_X1 U777 ( .A(G1986), .B(G290), .Z(n974) );
  NAND2_X1 U778 ( .A1(G160), .A2(G40), .ZN(n722) );
  NOR2_X1 U779 ( .A1(n721), .A2(n722), .ZN(n823) );
  INV_X1 U780 ( .A(n823), .ZN(n709) );
  OR2_X1 U781 ( .A1(n974), .A2(n709), .ZN(n811) );
  XNOR2_X1 U782 ( .A(KEYINPUT88), .B(G1991), .ZN(n949) );
  NAND2_X1 U783 ( .A1(G119), .A2(n877), .ZN(n691) );
  NAND2_X1 U784 ( .A1(G107), .A2(n878), .ZN(n690) );
  NAND2_X1 U785 ( .A1(n691), .A2(n690), .ZN(n696) );
  NAND2_X1 U786 ( .A1(G131), .A2(n875), .ZN(n693) );
  NAND2_X1 U787 ( .A1(G95), .A2(n883), .ZN(n692) );
  NAND2_X1 U788 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U789 ( .A(KEYINPUT87), .B(n694), .Z(n695) );
  OR2_X1 U790 ( .A1(n696), .A2(n695), .ZN(n871) );
  AND2_X1 U791 ( .A1(n949), .A2(n871), .ZN(n697) );
  XNOR2_X1 U792 ( .A(n697), .B(KEYINPUT89), .ZN(n707) );
  NAND2_X1 U793 ( .A1(G105), .A2(n883), .ZN(n698) );
  XNOR2_X1 U794 ( .A(n698), .B(KEYINPUT38), .ZN(n705) );
  NAND2_X1 U795 ( .A1(G141), .A2(n875), .ZN(n700) );
  NAND2_X1 U796 ( .A1(G129), .A2(n877), .ZN(n699) );
  NAND2_X1 U797 ( .A1(n700), .A2(n699), .ZN(n703) );
  NAND2_X1 U798 ( .A1(n878), .A2(G117), .ZN(n701) );
  XOR2_X1 U799 ( .A(KEYINPUT90), .B(n701), .Z(n702) );
  NOR2_X1 U800 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U801 ( .A1(n705), .A2(n704), .ZN(n893) );
  NAND2_X1 U802 ( .A1(G1996), .A2(n893), .ZN(n706) );
  NAND2_X1 U803 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U804 ( .A(KEYINPUT91), .B(n708), .ZN(n930) );
  NOR2_X1 U805 ( .A1(n930), .A2(n709), .ZN(n815) );
  XOR2_X1 U806 ( .A(KEYINPUT92), .B(n815), .Z(n720) );
  XNOR2_X1 U807 ( .A(G2067), .B(KEYINPUT37), .ZN(n710) );
  XNOR2_X1 U808 ( .A(n710), .B(KEYINPUT86), .ZN(n812) );
  NAND2_X1 U809 ( .A1(G140), .A2(n875), .ZN(n712) );
  NAND2_X1 U810 ( .A1(G104), .A2(n883), .ZN(n711) );
  NAND2_X1 U811 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U812 ( .A(KEYINPUT34), .B(n713), .ZN(n718) );
  NAND2_X1 U813 ( .A1(G128), .A2(n877), .ZN(n715) );
  NAND2_X1 U814 ( .A1(G116), .A2(n878), .ZN(n714) );
  NAND2_X1 U815 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U816 ( .A(KEYINPUT35), .B(n716), .Z(n717) );
  NOR2_X1 U817 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U818 ( .A(KEYINPUT36), .B(n719), .ZN(n896) );
  NOR2_X1 U819 ( .A1(n812), .A2(n896), .ZN(n925) );
  NAND2_X1 U820 ( .A1(n823), .A2(n925), .ZN(n819) );
  NAND2_X1 U821 ( .A1(n720), .A2(n819), .ZN(n809) );
  OR2_X1 U822 ( .A1(G1981), .A2(G305), .ZN(n790) );
  XOR2_X1 U823 ( .A(KEYINPUT24), .B(n790), .Z(n725) );
  INV_X1 U824 ( .A(n721), .ZN(n723) );
  NOR2_X4 U825 ( .A1(n723), .A2(n722), .ZN(n750) );
  INV_X1 U826 ( .A(n750), .ZN(n773) );
  INV_X1 U827 ( .A(n786), .ZN(n799) );
  NAND2_X1 U828 ( .A1(n725), .A2(n799), .ZN(n788) );
  NOR2_X1 U829 ( .A1(G2090), .A2(G303), .ZN(n726) );
  NAND2_X1 U830 ( .A1(G8), .A2(n726), .ZN(n727) );
  XNOR2_X1 U831 ( .A(n727), .B(KEYINPUT98), .ZN(n784) );
  NOR2_X1 U832 ( .A1(G2084), .A2(n773), .ZN(n728) );
  NAND2_X1 U833 ( .A1(G8), .A2(n728), .ZN(n771) );
  NOR2_X1 U834 ( .A1(G1966), .A2(n786), .ZN(n769) );
  NAND2_X1 U835 ( .A1(n729), .A2(G8), .ZN(n730) );
  XNOR2_X1 U836 ( .A(KEYINPUT30), .B(n730), .ZN(n731) );
  NOR2_X1 U837 ( .A1(G168), .A2(n731), .ZN(n736) );
  XNOR2_X1 U838 ( .A(G2078), .B(KEYINPUT25), .ZN(n943) );
  NAND2_X1 U839 ( .A1(n750), .A2(n943), .ZN(n732) );
  XNOR2_X1 U840 ( .A(n732), .B(KEYINPUT94), .ZN(n734) );
  OR2_X1 U841 ( .A1(G1961), .A2(n750), .ZN(n733) );
  NAND2_X1 U842 ( .A1(n734), .A2(n733), .ZN(n739) );
  NOR2_X1 U843 ( .A1(G171), .A2(n739), .ZN(n735) );
  NOR2_X1 U844 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U845 ( .A1(n739), .A2(G171), .ZN(n765) );
  INV_X1 U846 ( .A(G299), .ZN(n745) );
  NAND2_X1 U847 ( .A1(n750), .A2(G2072), .ZN(n740) );
  XNOR2_X1 U848 ( .A(n740), .B(KEYINPUT27), .ZN(n742) );
  INV_X1 U849 ( .A(G1956), .ZN(n845) );
  NOR2_X1 U850 ( .A1(n845), .A2(n750), .ZN(n741) );
  NOR2_X1 U851 ( .A1(n742), .A2(n741), .ZN(n744) );
  NOR2_X1 U852 ( .A1(n745), .A2(n744), .ZN(n743) );
  XOR2_X1 U853 ( .A(n743), .B(KEYINPUT28), .Z(n762) );
  NAND2_X1 U854 ( .A1(n745), .A2(n744), .ZN(n760) );
  AND2_X1 U855 ( .A1(n750), .A2(G1996), .ZN(n746) );
  XOR2_X1 U856 ( .A(n746), .B(KEYINPUT26), .Z(n748) );
  NAND2_X1 U857 ( .A1(n773), .A2(G1341), .ZN(n747) );
  NAND2_X1 U858 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U859 ( .A1(n975), .A2(n749), .ZN(n754) );
  NAND2_X1 U860 ( .A1(G1348), .A2(n773), .ZN(n752) );
  NAND2_X1 U861 ( .A1(G2067), .A2(n750), .ZN(n751) );
  NAND2_X1 U862 ( .A1(n752), .A2(n751), .ZN(n755) );
  NOR2_X1 U863 ( .A1(n756), .A2(n755), .ZN(n753) );
  OR2_X1 U864 ( .A1(n754), .A2(n753), .ZN(n758) );
  NAND2_X1 U865 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U866 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U867 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U868 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U869 ( .A(KEYINPUT29), .B(n763), .Z(n764) );
  NAND2_X1 U870 ( .A1(n765), .A2(n764), .ZN(n766) );
  INV_X1 U871 ( .A(n772), .ZN(n768) );
  NOR2_X1 U872 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U873 ( .A1(n771), .A2(n770), .ZN(n783) );
  XOR2_X1 U874 ( .A(KEYINPUT32), .B(KEYINPUT95), .Z(n781) );
  NAND2_X1 U875 ( .A1(n772), .A2(G286), .ZN(n778) );
  NOR2_X1 U876 ( .A1(G1971), .A2(n786), .ZN(n775) );
  NOR2_X1 U877 ( .A1(G2090), .A2(n773), .ZN(n774) );
  NOR2_X1 U878 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U879 ( .A1(n776), .A2(G303), .ZN(n777) );
  NAND2_X1 U880 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U881 ( .A1(n779), .A2(G8), .ZN(n780) );
  XNOR2_X1 U882 ( .A(n781), .B(n780), .ZN(n782) );
  NAND2_X1 U883 ( .A1(n783), .A2(n782), .ZN(n792) );
  NAND2_X1 U884 ( .A1(n784), .A2(n792), .ZN(n785) );
  NAND2_X1 U885 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U886 ( .A1(n788), .A2(n787), .ZN(n807) );
  NAND2_X1 U887 ( .A1(G1981), .A2(G305), .ZN(n789) );
  NAND2_X1 U888 ( .A1(n790), .A2(n789), .ZN(n984) );
  NOR2_X1 U889 ( .A1(G1976), .A2(G288), .ZN(n798) );
  NOR2_X1 U890 ( .A1(G1971), .A2(G303), .ZN(n791) );
  NOR2_X1 U891 ( .A1(n798), .A2(n791), .ZN(n973) );
  NAND2_X1 U892 ( .A1(n792), .A2(n973), .ZN(n793) );
  NAND2_X1 U893 ( .A1(G1976), .A2(G288), .ZN(n969) );
  NAND2_X1 U894 ( .A1(n793), .A2(n969), .ZN(n795) );
  NAND2_X1 U895 ( .A1(n796), .A2(n799), .ZN(n797) );
  INV_X1 U896 ( .A(KEYINPUT33), .ZN(n801) );
  NAND2_X1 U897 ( .A1(n797), .A2(n801), .ZN(n804) );
  NAND2_X1 U898 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U899 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U900 ( .A(n802), .B(KEYINPUT97), .ZN(n803) );
  NAND2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U902 ( .A1(n984), .A2(n805), .ZN(n806) );
  NOR2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n826) );
  NAND2_X1 U905 ( .A1(n812), .A2(n896), .ZN(n917) );
  NOR2_X1 U906 ( .A1(G1996), .A2(n893), .ZN(n932) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U908 ( .A1(n949), .A2(n871), .ZN(n920) );
  NOR2_X1 U909 ( .A1(n813), .A2(n920), .ZN(n814) );
  NOR2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U911 ( .A(KEYINPUT99), .B(n816), .Z(n817) );
  NOR2_X1 U912 ( .A1(n932), .A2(n817), .ZN(n818) );
  XNOR2_X1 U913 ( .A(n818), .B(KEYINPUT39), .ZN(n820) );
  NAND2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n917), .A2(n821), .ZN(n822) );
  XNOR2_X1 U916 ( .A(KEYINPUT100), .B(n822), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U919 ( .A(n827), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n912), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U922 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n830), .A2(n829), .ZN(G188) );
  XNOR2_X1 U925 ( .A(G120), .B(KEYINPUT103), .ZN(G236) );
  INV_X1 U927 ( .A(G108), .ZN(G238) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  NOR2_X1 U929 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U930 ( .A(G325), .ZN(G261) );
  XOR2_X1 U931 ( .A(G2096), .B(KEYINPUT43), .Z(n834) );
  XNOR2_X1 U932 ( .A(G2072), .B(KEYINPUT104), .ZN(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U934 ( .A(n835), .B(G2678), .Z(n837) );
  XNOR2_X1 U935 ( .A(G2067), .B(G2090), .ZN(n836) );
  XNOR2_X1 U936 ( .A(n837), .B(n836), .ZN(n842) );
  XNOR2_X1 U937 ( .A(KEYINPUT42), .B(n838), .ZN(n840) );
  XNOR2_X1 U938 ( .A(G2078), .B(G2084), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(G227) );
  XOR2_X1 U941 ( .A(G1976), .B(G1971), .Z(n844) );
  XNOR2_X1 U942 ( .A(G1991), .B(G1961), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n849) );
  XNOR2_X1 U944 ( .A(G1981), .B(n845), .ZN(n847) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1966), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U947 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U948 ( .A(G2474), .B(KEYINPUT41), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U950 ( .A(KEYINPUT105), .B(n852), .ZN(n853) );
  XOR2_X1 U951 ( .A(n853), .B(G1996), .Z(G229) );
  NAND2_X1 U952 ( .A1(G100), .A2(n883), .ZN(n855) );
  NAND2_X1 U953 ( .A1(G112), .A2(n878), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n855), .A2(n854), .ZN(n863) );
  XOR2_X1 U955 ( .A(KEYINPUT44), .B(KEYINPUT106), .Z(n857) );
  NAND2_X1 U956 ( .A1(G124), .A2(n877), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n860) );
  NAND2_X1 U958 ( .A1(n875), .A2(G136), .ZN(n858) );
  XNOR2_X1 U959 ( .A(KEYINPUT107), .B(n858), .ZN(n859) );
  NOR2_X1 U960 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U961 ( .A(KEYINPUT108), .B(n861), .Z(n862) );
  NOR2_X1 U962 ( .A1(n863), .A2(n862), .ZN(G162) );
  NAND2_X1 U963 ( .A1(G130), .A2(n877), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G118), .A2(n878), .ZN(n864) );
  NAND2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n870) );
  NAND2_X1 U966 ( .A1(G142), .A2(n875), .ZN(n867) );
  NAND2_X1 U967 ( .A1(G106), .A2(n883), .ZN(n866) );
  NAND2_X1 U968 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U969 ( .A(n868), .B(KEYINPUT45), .Z(n869) );
  NOR2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n872) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n892) );
  XOR2_X1 U972 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n874) );
  XNOR2_X1 U973 ( .A(G164), .B(KEYINPUT111), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(n888) );
  NAND2_X1 U975 ( .A1(n875), .A2(G139), .ZN(n876) );
  XNOR2_X1 U976 ( .A(KEYINPUT109), .B(n876), .ZN(n887) );
  NAND2_X1 U977 ( .A1(G127), .A2(n877), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G115), .A2(n878), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U980 ( .A(n881), .B(KEYINPUT110), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n882), .B(KEYINPUT47), .ZN(n885) );
  NAND2_X1 U982 ( .A1(n883), .A2(G103), .ZN(n884) );
  NAND2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n886) );
  NOR2_X1 U984 ( .A1(n887), .A2(n886), .ZN(n913) );
  XOR2_X1 U985 ( .A(n888), .B(n913), .Z(n890) );
  XNOR2_X1 U986 ( .A(G160), .B(n919), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n892), .B(n891), .ZN(n895) );
  XNOR2_X1 U989 ( .A(n893), .B(G162), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n895), .B(n894), .ZN(n897) );
  XOR2_X1 U991 ( .A(n897), .B(n896), .Z(n898) );
  NOR2_X1 U992 ( .A1(G37), .A2(n898), .ZN(G395) );
  XNOR2_X1 U993 ( .A(G286), .B(n975), .ZN(n900) );
  XNOR2_X1 U994 ( .A(n900), .B(n899), .ZN(n902) );
  XOR2_X1 U995 ( .A(n970), .B(G171), .Z(n901) );
  XNOR2_X1 U996 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U997 ( .A1(G37), .A2(n903), .ZN(G397) );
  NOR2_X1 U998 ( .A1(G227), .A2(G229), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n904), .B(KEYINPUT49), .ZN(n907) );
  NOR2_X1 U1000 ( .A1(G395), .A2(G397), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n905), .B(KEYINPUT113), .ZN(n906) );
  NOR2_X1 U1002 ( .A1(n907), .A2(n906), .ZN(n910) );
  NOR2_X1 U1003 ( .A1(G401), .A2(n911), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n908), .B(KEYINPUT112), .ZN(n909) );
  NAND2_X1 U1005 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(G303), .ZN(G166) );
  INV_X1 U1008 ( .A(n911), .ZN(G319) );
  INV_X1 U1009 ( .A(G69), .ZN(G235) );
  INV_X1 U1010 ( .A(n912), .ZN(G223) );
  XOR2_X1 U1011 ( .A(G2072), .B(n913), .Z(n915) );
  XOR2_X1 U1012 ( .A(G164), .B(G2078), .Z(n914) );
  NOR2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(n916), .B(KEYINPUT50), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(n928) );
  XNOR2_X1 U1016 ( .A(G160), .B(G2084), .ZN(n922) );
  NOR2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(KEYINPUT114), .B(n923), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1021 ( .A(KEYINPUT115), .B(n926), .ZN(n927) );
  NOR2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1023 ( .A1(n930), .A2(n929), .ZN(n936) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1025 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1026 ( .A(KEYINPUT51), .B(n933), .Z(n934) );
  XOR2_X1 U1027 ( .A(KEYINPUT116), .B(n934), .Z(n935) );
  NOR2_X1 U1028 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1029 ( .A(KEYINPUT52), .B(n937), .ZN(n938) );
  INV_X1 U1030 ( .A(KEYINPUT55), .ZN(n961) );
  NAND2_X1 U1031 ( .A1(n938), .A2(n961), .ZN(n939) );
  NAND2_X1 U1032 ( .A1(n939), .A2(G29), .ZN(n1022) );
  XNOR2_X1 U1033 ( .A(G29), .B(KEYINPUT121), .ZN(n964) );
  XNOR2_X1 U1034 ( .A(G2067), .B(G26), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(G33), .B(G2072), .ZN(n940) );
  NOR2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n948) );
  XOR2_X1 U1037 ( .A(G32), .B(G1996), .Z(n942) );
  NAND2_X1 U1038 ( .A1(n942), .A2(G28), .ZN(n946) );
  XOR2_X1 U1039 ( .A(G27), .B(n943), .Z(n944) );
  XNOR2_X1 U1040 ( .A(KEYINPUT118), .B(n944), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(G25), .B(n949), .ZN(n950) );
  NOR2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1045 ( .A(KEYINPUT53), .B(n952), .Z(n956) );
  XNOR2_X1 U1046 ( .A(KEYINPUT54), .B(G34), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(n953), .B(KEYINPUT119), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(G2084), .B(n954), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n959) );
  XOR2_X1 U1050 ( .A(KEYINPUT117), .B(G2090), .Z(n957) );
  XNOR2_X1 U1051 ( .A(G35), .B(n957), .ZN(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1053 ( .A(n961), .B(n960), .Z(n962) );
  XNOR2_X1 U1054 ( .A(n962), .B(KEYINPUT120), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1056 ( .A1(n965), .A2(G11), .ZN(n1020) );
  INV_X1 U1057 ( .A(G16), .ZN(n1016) );
  XOR2_X1 U1058 ( .A(n1016), .B(KEYINPUT56), .Z(n990) );
  XOR2_X1 U1059 ( .A(G299), .B(G1956), .Z(n967) );
  XOR2_X1 U1060 ( .A(G301), .B(G1961), .Z(n966) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n981) );
  NAND2_X1 U1062 ( .A1(G1971), .A2(G303), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n972) );
  XOR2_X1 U1064 ( .A(G1348), .B(n970), .Z(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n979) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n977) );
  XNOR2_X1 U1067 ( .A(G1341), .B(n975), .ZN(n976) );
  NOR2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1071 ( .A(KEYINPUT123), .B(n982), .Z(n988) );
  XOR2_X1 U1072 ( .A(G168), .B(G1966), .Z(n983) );
  NOR2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1074 ( .A(KEYINPUT57), .B(n985), .Z(n986) );
  XNOR2_X1 U1075 ( .A(KEYINPUT122), .B(n986), .ZN(n987) );
  NAND2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n990), .A2(n989), .ZN(n1018) );
  XNOR2_X1 U1078 ( .A(G1961), .B(KEYINPUT124), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(n991), .B(G5), .ZN(n1002) );
  XNOR2_X1 U1080 ( .A(KEYINPUT59), .B(G1348), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(n992), .B(G4), .ZN(n998) );
  XOR2_X1 U1082 ( .A(G1341), .B(G19), .Z(n994) );
  XOR2_X1 U1083 ( .A(G1956), .B(G20), .Z(n993) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(G6), .B(G1981), .ZN(n995) );
  NOR2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1088 ( .A(n999), .B(KEYINPUT60), .Z(n1000) );
  XNOR2_X1 U1089 ( .A(KEYINPUT125), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XOR2_X1 U1091 ( .A(G1966), .B(KEYINPUT126), .Z(n1003) );
  XNOR2_X1 U1092 ( .A(G21), .B(n1003), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1013) );
  XNOR2_X1 U1094 ( .A(G1986), .B(G24), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G23), .B(G1976), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(G1971), .B(KEYINPUT127), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(n1008), .B(G22), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1023), .ZN(G150) );
  INV_X1 U1108 ( .A(G150), .ZN(G311) );
endmodule

