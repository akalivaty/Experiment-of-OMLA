//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n561,
    new_n562, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n590, new_n591, new_n594, new_n596, new_n597, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1140, new_n1141;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(G137), .ZN(new_n467));
  NAND2_X1  g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(G160));
  OR2_X1    g045(.A1(G100), .A2(G2105), .ZN(new_n471));
  OAI211_X1 g046(.A(new_n471), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT64), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT3), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(new_n462), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n478), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n473), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT65), .ZN(G162));
  NAND3_X1  g059(.A1(new_n462), .A2(G102), .A3(G2104), .ZN(new_n485));
  AND2_X1   g060(.A1(G114), .A2(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(new_n463), .B2(G126), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n485), .B1(new_n487), .B2(new_n462), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n475), .A2(new_n477), .A3(G138), .A4(new_n462), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n463), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n488), .A2(new_n493), .ZN(G164));
  NAND2_X1  g069(.A1(G75), .A2(G543), .ZN(new_n495));
  NAND2_X1  g070(.A1(KEYINPUT66), .A2(KEYINPUT5), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G543), .ZN(new_n497));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(KEYINPUT66), .A3(KEYINPUT5), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G62), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n495), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G651), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT67), .B(G88), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n506), .A2(new_n498), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n503), .B(new_n509), .C1(new_n510), .C2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  AND2_X1   g089(.A1(new_n497), .A2(new_n499), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n511), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n511), .A2(new_n518), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G51), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT69), .B(KEYINPUT7), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT70), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n526), .B(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n507), .A2(G89), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n528), .A2(KEYINPUT71), .A3(new_n529), .ZN(new_n533));
  AOI211_X1 g108(.A(new_n517), .B(new_n524), .C1(new_n532), .C2(new_n533), .ZN(G168));
  AOI22_X1  g109(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  INV_X1    g113(.A(new_n507), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n520), .A2(new_n521), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI221_X1 g116(.A(new_n537), .B1(new_n538), .B2(new_n539), .C1(new_n540), .C2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(new_n507), .A2(G81), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n545), .B2(new_n536), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n546), .B1(new_n522), .B2(G43), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(new_n507), .A2(G91), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  NOR3_X1   g131(.A1(new_n512), .A2(KEYINPUT9), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n511), .B2(G53), .ZN(new_n559));
  OAI221_X1 g134(.A(new_n554), .B1(new_n555), .B2(new_n536), .C1(new_n557), .C2(new_n559), .ZN(G299));
  INV_X1    g135(.A(new_n533), .ZN(new_n561));
  AOI21_X1  g136(.A(KEYINPUT71), .B1(new_n528), .B2(new_n529), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n516), .B(new_n523), .C1(new_n561), .C2(new_n562), .ZN(G286));
  NAND2_X1  g138(.A1(new_n507), .A2(G87), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n565));
  INV_X1    g140(.A(G49), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n564), .B(new_n565), .C1(new_n566), .C2(new_n512), .ZN(G288));
  NAND2_X1  g142(.A1(new_n511), .A2(G48), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT72), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n568), .B(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(new_n536), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n507), .A2(G86), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(G305));
  AOI22_X1  g149(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n536), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT73), .Z(new_n577));
  NAND2_X1  g152(.A1(new_n507), .A2(G85), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n522), .A2(G47), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G290));
  NAND2_X1  g155(.A1(G301), .A2(G868), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n522), .A2(G54), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n507), .A2(G92), .ZN(new_n583));
  XOR2_X1   g158(.A(new_n583), .B(KEYINPUT10), .Z(new_n584));
  AOI22_X1  g159(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n582), .B(new_n584), .C1(new_n536), .C2(new_n585), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT74), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n581), .B1(new_n587), .B2(G868), .ZN(G284));
  XNOR2_X1  g163(.A(G284), .B(KEYINPUT75), .ZN(G321));
  INV_X1    g164(.A(G868), .ZN(new_n590));
  NAND2_X1  g165(.A1(G299), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n591), .B1(G168), .B2(new_n590), .ZN(G297));
  OAI21_X1  g167(.A(new_n591), .B1(G168), .B2(new_n590), .ZN(G280));
  INV_X1    g168(.A(G559), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n587), .B1(new_n594), .B2(G860), .ZN(G148));
  NAND2_X1  g170(.A1(new_n587), .A2(new_n594), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G868), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g173(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g174(.A1(new_n479), .A2(G123), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n481), .A2(G135), .ZN(new_n601));
  NOR2_X1   g176(.A1(G99), .A2(G2105), .ZN(new_n602));
  OAI21_X1  g177(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n600), .B(new_n601), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(G2096), .Z(new_n605));
  XOR2_X1   g180(.A(KEYINPUT76), .B(KEYINPUT12), .Z(new_n606));
  NOR3_X1   g181(.A1(new_n476), .A2(new_n474), .A3(G2105), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g183(.A(KEYINPUT13), .B(G2100), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n605), .A2(new_n610), .ZN(G156));
  XNOR2_X1  g186(.A(G2451), .B(G2454), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT16), .ZN(new_n613));
  XOR2_X1   g188(.A(G2443), .B(G2446), .Z(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(G1341), .B(G1348), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(G2427), .B(G2438), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2430), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT15), .B(G2435), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(KEYINPUT14), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n617), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G14), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT77), .Z(G401));
  XOR2_X1   g200(.A(G2067), .B(G2678), .Z(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G2084), .B(G2090), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AND2_X1   g204(.A1(new_n629), .A2(KEYINPUT17), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n627), .A2(new_n628), .ZN(new_n631));
  AOI21_X1  g206(.A(KEYINPUT18), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2072), .B(G2078), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n629), .A2(KEYINPUT18), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n632), .B2(new_n633), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2100), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT78), .B(G2096), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(G227));
  XNOR2_X1  g214(.A(G1971), .B(G1976), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT19), .ZN(new_n641));
  XOR2_X1   g216(.A(G1956), .B(G2474), .Z(new_n642));
  XOR2_X1   g217(.A(G1961), .B(G1966), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT79), .B(KEYINPUT20), .Z(new_n646));
  INV_X1    g221(.A(new_n641), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n642), .A2(new_n643), .ZN(new_n648));
  AOI22_X1  g223(.A1(new_n645), .A2(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n650), .A2(new_n641), .A3(new_n644), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n649), .B(new_n651), .C1(new_n645), .C2(new_n646), .ZN(new_n652));
  XOR2_X1   g227(.A(G1991), .B(G1996), .Z(new_n653));
  XNOR2_X1  g228(.A(G1981), .B(G1986), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT80), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n656), .B(new_n658), .ZN(G229));
  NAND2_X1  g234(.A1(KEYINPUT24), .A2(G34), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(KEYINPUT24), .A2(G34), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n661), .A2(new_n662), .A3(G29), .ZN(new_n663));
  INV_X1    g238(.A(G160), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n663), .B1(new_n664), .B2(G29), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n666), .A2(G2084), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT27), .B(G1996), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT86), .ZN(new_n669));
  OR2_X1    g244(.A1(G29), .A2(G32), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n479), .A2(G129), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n481), .A2(G141), .ZN(new_n672));
  NAND3_X1  g247(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT26), .Z(new_n674));
  NAND3_X1  g249(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT85), .ZN(new_n676));
  NAND4_X1  g251(.A1(new_n671), .A2(new_n672), .A3(new_n674), .A4(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(G29), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n670), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(G5), .A2(G16), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(G171), .B2(G16), .ZN(new_n681));
  OAI221_X1 g256(.A(new_n667), .B1(new_n669), .B2(new_n679), .C1(new_n681), .C2(G1961), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT89), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G4), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(new_n587), .B2(new_n685), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n687), .A2(G1348), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G162), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G29), .ZN(new_n691));
  INV_X1    g266(.A(G35), .ZN(new_n692));
  OAI21_X1  g267(.A(KEYINPUT91), .B1(new_n692), .B2(G29), .ZN(new_n693));
  OR3_X1    g268(.A1(new_n692), .A2(KEYINPUT91), .A3(G29), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(KEYINPUT29), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT29), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n691), .A2(new_n697), .A3(new_n693), .A4(new_n694), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n699), .A2(G2090), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n687), .A2(G1348), .ZN(new_n701));
  OR2_X1    g276(.A1(G29), .A2(G33), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT25), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n481), .A2(G139), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n704), .B(new_n705), .C1(new_n462), .C2(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n702), .B1(new_n707), .B2(new_n678), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(G2072), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT84), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n685), .A2(G19), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n547), .B2(new_n685), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n711), .B1(G1341), .B2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G27), .ZN(new_n715));
  OAI21_X1  g290(.A(KEYINPUT90), .B1(new_n715), .B2(G29), .ZN(new_n716));
  OR3_X1    g291(.A1(new_n715), .A2(KEYINPUT90), .A3(G29), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n716), .B(new_n717), .C1(G164), .C2(new_n678), .ZN(new_n718));
  INV_X1    g293(.A(G2078), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n709), .A2(G2072), .B1(new_n669), .B2(new_n679), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n666), .A2(G2084), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n713), .A2(G1341), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n678), .A2(G26), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n479), .A2(G128), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n481), .A2(G140), .ZN(new_n727));
  OR2_X1    g302(.A1(G104), .A2(G2105), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n728), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n725), .B1(new_n731), .B2(new_n678), .ZN(new_n732));
  MUX2_X1   g307(.A(new_n725), .B(new_n732), .S(KEYINPUT28), .Z(new_n733));
  AND2_X1   g308(.A1(new_n733), .A2(G2067), .ZN(new_n734));
  NOR4_X1   g309(.A1(new_n714), .A2(new_n723), .A3(new_n724), .A4(new_n734), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n689), .A2(new_n700), .A3(new_n701), .A4(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT23), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n685), .A2(G20), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n737), .B(new_n738), .C1(G299), .C2(G16), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n737), .B2(new_n738), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT93), .B(G1956), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT92), .ZN(new_n743));
  AND3_X1   g318(.A1(new_n699), .A2(new_n743), .A3(G2090), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n743), .B1(new_n699), .B2(G2090), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT94), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g323(.A(KEYINPUT94), .B(new_n742), .C1(new_n744), .C2(new_n745), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n736), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n733), .A2(G2067), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT31), .B(G11), .ZN(new_n752));
  INV_X1    g327(.A(G28), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n753), .B2(KEYINPUT30), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(KEYINPUT30), .B2(new_n753), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n604), .B2(new_n678), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n681), .B2(G1961), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT87), .ZN(new_n758));
  NAND3_X1  g333(.A1(G168), .A2(new_n758), .A3(G16), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(G16), .B2(G21), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G286), .B2(new_n685), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(G1966), .ZN(new_n763));
  INV_X1    g338(.A(G1966), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n759), .B2(new_n761), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n752), .B(new_n757), .C1(new_n763), .C2(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT88), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n750), .A2(new_n751), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(KEYINPUT95), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT95), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n750), .A2(new_n770), .A3(new_n751), .A4(new_n767), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n685), .A2(G23), .ZN(new_n772));
  INV_X1    g347(.A(G288), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n685), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT33), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1976), .ZN(new_n776));
  MUX2_X1   g351(.A(G6), .B(G305), .S(G16), .Z(new_n777));
  XOR2_X1   g352(.A(KEYINPUT32), .B(G1981), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n685), .A2(G22), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G166), .B2(new_n685), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT83), .B(G1971), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n776), .A2(new_n779), .A3(new_n783), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT34), .Z(new_n785));
  NOR2_X1   g360(.A1(G16), .A2(G24), .ZN(new_n786));
  XOR2_X1   g361(.A(G290), .B(KEYINPUT82), .Z(new_n787));
  AOI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(G16), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(G1986), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n479), .A2(G119), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n481), .A2(G131), .ZN(new_n791));
  NOR2_X1   g366(.A1(G95), .A2(G2105), .ZN(new_n792));
  OAI21_X1  g367(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n790), .B(new_n791), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  MUX2_X1   g369(.A(G25), .B(new_n794), .S(G29), .Z(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT35), .B(G1991), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT81), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n795), .B(new_n797), .Z(new_n798));
  NAND3_X1  g373(.A1(new_n785), .A2(new_n789), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(KEYINPUT36), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n799), .A2(KEYINPUT36), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n769), .A2(new_n771), .B1(new_n800), .B2(new_n801), .ZN(G311));
  NAND2_X1  g377(.A1(new_n769), .A2(new_n771), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n800), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(G150));
  NAND2_X1  g380(.A1(new_n507), .A2(G93), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(new_n536), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n522), .B2(G55), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(G860), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT96), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT37), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n587), .A2(G559), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT38), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n547), .B(new_n809), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT39), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n815), .B(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n813), .B1(new_n818), .B2(G860), .ZN(G145));
  XNOR2_X1  g394(.A(G164), .B(new_n608), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n479), .A2(G130), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n481), .A2(G142), .ZN(new_n823));
  OR2_X1    g398(.A1(G106), .A2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n824), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n794), .B(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(new_n677), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n707), .B(new_n730), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n827), .A2(new_n677), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n830), .B1(new_n828), .B2(new_n831), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n821), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n828), .A2(new_n831), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(new_n829), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n836), .A2(new_n820), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT97), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n834), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G162), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n834), .A2(new_n838), .A3(new_n839), .A4(new_n690), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n604), .B(G160), .Z(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G37), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n841), .A2(new_n844), .A3(new_n842), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n846), .A2(KEYINPUT98), .A3(new_n847), .A4(new_n848), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g429(.A1(new_n810), .A2(new_n590), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n773), .B(G303), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(G305), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(G290), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT99), .ZN(new_n859));
  MUX2_X1   g434(.A(new_n858), .B(new_n859), .S(KEYINPUT42), .Z(new_n860));
  INV_X1    g435(.A(new_n816), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n596), .B(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n586), .A2(G299), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n586), .A2(G299), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n865), .A2(KEYINPUT41), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT41), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(new_n863), .B2(new_n864), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n867), .B1(new_n871), .B2(new_n862), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n860), .B(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n855), .B1(new_n873), .B2(new_n590), .ZN(G295));
  OAI21_X1  g449(.A(new_n855), .B1(new_n873), .B2(new_n590), .ZN(G331));
  INV_X1    g450(.A(new_n859), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n868), .A2(KEYINPUT103), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n868), .A2(KEYINPUT103), .A3(new_n870), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n879));
  NAND3_X1  g454(.A1(G286), .A2(new_n879), .A3(G301), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n524), .B1(new_n532), .B2(new_n533), .ZN(new_n881));
  NAND2_X1  g456(.A1(G171), .A2(KEYINPUT100), .ZN(new_n882));
  NAND2_X1  g457(.A1(G301), .A2(new_n879), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n516), .A4(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n861), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n880), .A2(new_n884), .A3(new_n861), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT102), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n880), .A2(new_n884), .A3(new_n890), .A4(new_n861), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  AOI211_X1 g467(.A(new_n877), .B(new_n878), .C1(new_n887), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n880), .A2(new_n884), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n816), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n888), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT104), .B1(new_n896), .B2(new_n865), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n895), .A2(new_n898), .A3(new_n866), .A4(new_n888), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n876), .B1(new_n893), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n895), .A2(new_n886), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n885), .A2(KEYINPUT101), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n892), .A2(new_n902), .A3(new_n866), .A4(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n896), .B1(new_n868), .B2(new_n870), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n859), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n906), .A2(new_n847), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n901), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n847), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n859), .B1(new_n905), .B2(new_n904), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT43), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n904), .A2(new_n905), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n876), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n917), .A2(new_n908), .A3(new_n847), .A4(new_n906), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n914), .B1(new_n918), .B2(KEYINPUT105), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n877), .B1(new_n887), .B2(new_n892), .ZN(new_n920));
  INV_X1    g495(.A(new_n878), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n900), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n859), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT43), .B1(new_n924), .B2(new_n910), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n907), .A2(new_n926), .A3(new_n908), .A4(new_n917), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n919), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n915), .A2(new_n928), .ZN(G397));
  INV_X1    g504(.A(G1384), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(new_n488), .B2(new_n493), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XOR2_X1   g508(.A(KEYINPUT106), .B(G40), .Z(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(G160), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n730), .B(G2067), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(KEYINPUT108), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(G1996), .A3(new_n677), .ZN(new_n941));
  INV_X1    g516(.A(new_n937), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n942), .A2(G1996), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT107), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n940), .B(new_n941), .C1(new_n944), .C2(new_n677), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n794), .B(new_n797), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n945), .B1(new_n937), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(G290), .A2(G1986), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n937), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT48), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n937), .B1(new_n677), .B2(new_n938), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n944), .A2(KEYINPUT46), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n944), .A2(KEYINPUT46), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n955), .B(KEYINPUT47), .Z(new_n956));
  OR2_X1    g531(.A1(new_n794), .A2(new_n797), .ZN(new_n957));
  OAI22_X1  g532(.A1(new_n945), .A2(new_n957), .B1(G2067), .B2(new_n730), .ZN(new_n958));
  AOI211_X1 g533(.A(new_n951), .B(new_n956), .C1(new_n937), .C2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n931), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n936), .B1(new_n960), .B2(KEYINPUT45), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n931), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g538(.A(KEYINPUT109), .B(new_n930), .C1(new_n488), .C2(new_n493), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n961), .B1(new_n965), .B2(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n764), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n936), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n931), .A2(KEYINPUT50), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT114), .B(G2084), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n969), .A2(new_n970), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(G168), .A2(new_n967), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT120), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(new_n975), .A3(G8), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT121), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n974), .A2(KEYINPUT121), .A3(G8), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G8), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(new_n967), .B2(new_n973), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(G286), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n976), .A2(new_n977), .A3(KEYINPUT51), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n981), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT62), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n988));
  OR3_X1    g563(.A1(new_n966), .A2(new_n988), .A3(G2078), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n961), .A2(new_n719), .A3(new_n933), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n988), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT122), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n993));
  INV_X1    g568(.A(G1961), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT122), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n990), .A2(new_n996), .A3(new_n988), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n989), .A2(new_n992), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n998), .A2(G171), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n1000));
  NAND3_X1  g575(.A1(G303), .A2(new_n1000), .A3(G8), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1000), .B1(G303), .B2(G8), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT111), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1003), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(new_n1001), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1971), .ZN(new_n1009));
  INV_X1    g584(.A(new_n961), .ZN(new_n1010));
  INV_X1    g585(.A(new_n933), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT110), .B(G2090), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n969), .A2(new_n970), .A3(new_n971), .A4(new_n1014), .ZN(new_n1015));
  AOI211_X1 g590(.A(new_n982), .B(new_n1008), .C1(new_n1012), .C2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G305), .A2(G1981), .ZN(new_n1017));
  INV_X1    g592(.A(G1981), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n570), .A2(new_n1018), .A3(new_n572), .A4(new_n573), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT49), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n965), .A2(new_n970), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1017), .A2(KEYINPUT49), .A3(new_n1019), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(G8), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(G8), .ZN(new_n1026));
  INV_X1    g601(.A(G1976), .ZN(new_n1027));
  NOR2_X1   g602(.A1(G288), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT52), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1028), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT52), .B1(G288), .B2(new_n1027), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1023), .A2(G8), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1025), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1016), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT126), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n963), .A2(KEYINPUT50), .A3(new_n964), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT113), .B1(new_n1036), .B2(new_n970), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n960), .A2(new_n968), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1036), .A2(KEYINPUT113), .A3(new_n970), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1012), .B1(new_n1041), .B2(new_n1013), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1042), .A2(G8), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1034), .B(new_n1035), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n1042), .B2(G8), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1047), .A2(G8), .A3(new_n1004), .A4(new_n1007), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1048), .A2(new_n1029), .A3(new_n1025), .A4(new_n1032), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT126), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT62), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n981), .A2(new_n1052), .A3(new_n984), .A4(new_n985), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n987), .A2(new_n999), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1026), .B(KEYINPUT112), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1025), .A2(new_n1027), .A3(new_n773), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1055), .B1(new_n1056), .B2(new_n1019), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT63), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1034), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n983), .A2(G168), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1044), .B1(new_n1047), .B2(G8), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1049), .A2(new_n1058), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1063), .A2(G168), .A3(new_n983), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1057), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  OR2_X1    g640(.A1(new_n1033), .A2(new_n1048), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1054), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT56), .B(G2072), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n961), .A2(new_n933), .A3(new_n1068), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1036), .A2(KEYINPUT113), .A3(new_n970), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1039), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1070), .A2(new_n1037), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1069), .B1(new_n1072), .B2(G1956), .ZN(new_n1073));
  NAND2_X1  g648(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G299), .A2(new_n1074), .ZN(new_n1075));
  OR2_X1    g650(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1073), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1077), .B(new_n1069), .C1(new_n1072), .C2(G1956), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT61), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1073), .A2(KEYINPUT118), .A3(new_n1078), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT58), .B(G1341), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1023), .A2(KEYINPUT116), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n965), .A2(new_n1088), .A3(new_n970), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1086), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1010), .A2(G1996), .A3(new_n1011), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n547), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n1093));
  XNOR2_X1  g668(.A(new_n1092), .B(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1079), .A2(KEYINPUT61), .A3(new_n1081), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT119), .B1(new_n1085), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1098), .A2(new_n1099), .A3(new_n1095), .A4(new_n1094), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1101));
  INV_X1    g676(.A(G2067), .ZN(new_n1102));
  INV_X1    g677(.A(G1348), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1101), .A2(new_n1102), .B1(new_n1103), .B2(new_n993), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(KEYINPUT60), .B2(new_n587), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n587), .A2(KEYINPUT60), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1097), .A2(new_n1100), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1081), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(new_n1104), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1110), .A2(new_n587), .B1(new_n1078), .B2(new_n1073), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n960), .A2(KEYINPUT45), .ZN(new_n1114));
  AND2_X1   g689(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1115));
  NOR2_X1   g690(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1116));
  OAI211_X1 g691(.A(KEYINPUT53), .B(G40), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1114), .A2(G160), .A3(new_n933), .A4(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1119), .B(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1121), .A2(new_n995), .A3(new_n992), .A4(new_n997), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(G171), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1113), .B1(new_n1123), .B2(KEYINPUT127), .ZN(new_n1124));
  OAI221_X1 g699(.A(new_n1124), .B1(KEYINPUT127), .B2(new_n1123), .C1(G171), .C2(new_n998), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1122), .A2(G171), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1113), .B1(new_n999), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1125), .A2(new_n1129), .A3(new_n986), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1051), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1067), .B1(new_n1112), .B2(new_n1133), .ZN(new_n1134));
  AND2_X1   g709(.A1(G290), .A2(G1986), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n937), .B1(new_n1135), .B2(new_n948), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n947), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n959), .B1(new_n1134), .B2(new_n1137), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g713(.A(G401), .B(G229), .C1(new_n851), .C2(new_n852), .ZN(new_n1140));
  NOR2_X1   g714(.A1(G227), .A2(new_n460), .ZN(new_n1141));
  AND3_X1   g715(.A1(new_n1140), .A2(new_n913), .A3(new_n1141), .ZN(G308));
  NAND3_X1  g716(.A1(new_n1140), .A2(new_n913), .A3(new_n1141), .ZN(G225));
endmodule


